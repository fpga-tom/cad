// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tBmvaAGRYkciual7RTFk3+V+/aHrll69qupsewK38z0ysPDuWWwR81S3lJmHIMvE
CScJbSnELEqN/lLjKjgrGMEaCI4hhuaxIK7ijH1SU8aZjPnKiBH/JWnsMfPRWZWx
PmjBV+YIYeQj8HkDu7t+SRtgqsmdSyyYi5A3LYOVAhg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10000)
URfXXX1p/WnVJ8Fqf1NdpPMOIzKlxzPf1tn0uRinlHf9mXAYKalMEV4or1AxLAfL
ugxXDp46dB/lViJvoc4PCjBU4vNhXLjkfYkneJ3IBheRmkdIk/zJDzQfCI+HWqn9
0maiI+/EJUaUIxxCmPyuxD7dQtSw2FIKTGYHKy9lIEhYS4rNetsOjjGxz34WbYuU
7XGBdf43FWxRuiLsqwtU1ZXth3xvS2ervBRh1hfH48aPY7nTjjCmOA4+uit/QWjo
u+bH4XdpchknXpEbBcaxgLINw2TBroD6Rx/+PoOuTgllPGDKeBtUx5mL9a+EYPuL
iiQ6p6bOT2od0N9S2XWkTYj6w0nwbTppDBrWYNZClhq0zHhbMbQRI08vRsBP3xPr
t4zixpTbj8SvRg7kBSYGcqJ/jj7xuHl4b7nK8WwOTBcgns4jyqE3WQ2rKWLASifr
GegE/+5J9iETNtrZU9rPsmg34ixcjBgsFVW6vXkoznSMASxBzIHSWPrGmm6N7ddR
ylHh6u1MNUl0AtqhxYj6Jr/wi1bCyuoCM5qUWWoBChZw3QIriH3xhx3rrGIB26hN
P6R318YPmt0TjZxZnyNR/iWba+J3CmaYVSUrC1o2im6ADQ/gNSwEtZWG0Axcr8cV
e7C4P/kkh5eAMQz6eZzexaSg6BNNeWJ4TMiwHMAJvEWf4Hbzz391X71dgzWHo7tC
7Jc39ktNi4bVAtL+GUhNgaooXoTq4U3HTi5rJ+5XmEgeyTgRNPzaqT0wlloTgWL4
+Ybv7dMV6Ke69FYEbcap1PISy8g0Wjjclsxa7cJis4jw0RIqerQjlPkkNX22YR1N
PsoBRMAEY7sU6DBujAbUQhBEjH7wZh7ex+3EjnFC38wbjU5W5qExj4yAOuUegDA2
I9UZbO6jIqaiJw0e5XnvH1vysJmeewrA7LqpM/AbRdvxEo81oqolXx3noNuixWlp
CiltTM4bIPJjemrNC3iniZXdUnD2p+5Sv3G5+THIm9axMY0f4oJ5RqYJhKHpaIIU
hXDhhyCoRaF1LB7urXPPWcnq+2Mw2jjnwHQMwf36OcEhKd+Bjm2+7Ck3gtKPTEQj
deqM4fzWKD5yJ/Snrbha3ic3G4vLqHivAh98rifrF4GXaFIaVcZiz644MQ2k4/5j
awTfajWfiANPMwZK+/YrsnDEFd6OnoNuCBJAFVtT6mACGYrDYpH8g05PhjqjhjNR
wrf7T9nLCW/4XULB/jgw9G/RZrXleT6i3WPGC2gNP9AfhLF2qjVkn73a+UFPeUz1
QFrAyHTs0CVOgTOq5Lp9FDh+EA2J0yTjsSjwLjWeFgxdr7mUxKxJzFQjyrQpPBBO
B/In57DJW0VUIiAZBahE12KzmO/kQyS8h4M56HPcjpef53BCevJ6hj/0j6nxidPw
LsYDsdjwJOHfk/5dPjyfaDyaphogyV4z0hBEdQ/BOoLHtWRww/qsFF8ICAjDm9C7
MTGpP2NgYY4YaVmlcU9GwKJPK4MGx91F8DguFH/ia8CI30yd4NJrJ11m6V0v/urN
L2H1VOOhE3r6uwweZ2DQOWc+dOuS9BgCvk8SkXCkTFxIUg0K4fydV+tReO01PS2h
EISQup/Aao0rTC+ZDXLQGtbjHMbzqLXyOVC9wU1yCElUiie8y3NErC2PD+DVs37i
jOcfgcRiln8qVXDlGiHacph5p7eNaNxNSeU7mRCFREluYP5geNejEs9YH+yBrC42
WUqra8m7EGU0Dk3A3/yjY1ExDCG46tNyLUuEE2fW2Rj6zB9e7PWlNG2VmNQj3cun
qjjBRNLqK51WA+zrieguRehnUsLLIL4eB/BgGsoiPgPSv7pvvWiE1I4GvS7n4glE
IxJ5bsMK9yCSFGlJTl2xDX1kKpTn3woxI840DBfHSW1jitH3d7l2vGM1piP+Rjnu
J8+jvIjXcHiiMl5gIed5OQD7RvsfjFT4JZFkdfI0k4t3FzjWRpE9ZLbudo+/hNqM
1x25ldRV2HHIxNvpjWphevhCuhzkX+YoEIfV0a8S6by8DA65Ke3UmcFxoVv9kP9t
KktEVf4VSzXhNmjvlGO4RlJYKQGSnQO5WcqPOAIrRcqxs2++6C36IoAOO9uft8NY
wHTTTRdYOB9htlU9iyTuLMcQQQVkVxPdweVyfFLihvaZaTuRbOXbm6ALmRDSbEHo
ta3VUwN+LCP9YNaCEUjb2WZBAkdWGcM0+C1CgkbQ2B2ctxnyA0w56yuQV/B2erxw
xNKZimWPgFaf3yceOyb+wQUo2gLgwvZJp5Rzz/96H8ER1sMUnnwocIJbSWvbbFR0
gd6/gNohVUZm/ADfL0HZp/D+N0Jx2URdWCjYYTzviJ3uMU79VosRegp7vxSpXO8p
hD4OIMytrUOebIega7/ps4B2fLz/vS1iwCB0lYfyN57hUffG/UFTVYH+NhuUfeQx
f8xbMQCFKz4Y1graQ0A7DGtcvKVQNyddFUeNCSHP5VtXCDSueNyYOjmMfIxbDzYM
jEg++FFcv634sT8jlNtz/iDNZeJhIMrV/VvcWAY/Oja1llwzR5WVb9bj91tempdE
aUUBRMSs+37PTZI3SUWbjGPtlmAGPxITvY0M0NZKHZ/8cDApY9V5LxwZDR70T7gz
vllr6okc+5797p8/gjW4O6ranZgHRmLuY+WSpvgaRPPnOA1ehjolJZybTpmh1ykH
ZVLoe8hyqE3UZC5ST7yi07nYAxBfkZ6N8izDx7WxRfM7aMIdivCQP09yK6YL/L+L
p/3EZoYDpYFavkcqTHgb4wTkJzFlAOEN2vgt+wTKprndGIVaU/3H5jiIFeOX37pk
HuuLDo7IO6GbKl8wwDKkcUVxD/2yESUaY0JAOvxY4rolJbyCYBDtjqZ/tO2vghW9
JzunYVneJgZSCE+v8Kv+lIIt5pMmvqu6jmCp3K1W7mpi045+Z6orgV7VWWTS3SWn
3psKC2W7mbdx97Cfzs6bxFEd7wPzxYf3Dfp9T6uEBa9nnWOMhOK3ETdqg1hZ63FM
iWocKTOkTmgF6Qp6tmNbdpqUZqRzVfuOD7aZzbrlue+kat2AslD4IW5PGDkbjJmY
A6uBAMeEHYpaGalFY3yH0/CjgkZWBcdxV9IJ0kRWxQe09XFDuRfPWXT8en1991U/
EMaGmibRIs8pgcJEzvOfjPrLfHGRnT0Yy3hd10qobwnvzkgx+ehqQcoI2P1ULoou
ebHtdsgBH5cVJpxat0jT3zxbCGv9gJwWiKWcbMgyzwCBhht2c8tvqoC2DFwWQZC1
ConhsYWjIljM0jRb8brVS/i1HaiqfR1BWUDk2BYmZbv8U8jbwjfNVvWMeaqS5LJR
y62U7LpffVM5SkFBeCUV5DnLImedYQIv3IX00GEk4e2V1OGbfGUJX5xhtjFbTrhK
i5eJW8HUX3a7KxCrmPLVLzjzDK1FgRNkwtCsU5ju+c73KtVNjs8Eh4I54V3CvDxH
n8gqS3Apg42haGX9yamnKhwtLFmv0ti/sU5ne17mdGQOywEmtdWNRTP31aifQPyk
Y5IdX8Zvsl4sc3is7xfQgBVh1L1q54eMrMkLFwyV4vbvw+L1HXal81o9EDuLJtlQ
mw6zbB9Kk2N2QKsFIy8Kw+hlhxaql19TvsnarCSfpc50KOMA0DHu30swbGQNxDXh
TC+/ZK4BuBsk9jKW08eh7QgMwbXNQCjbxfbMdwU1HhqILIhipkGhnfiR31fxWa0O
qrLZSyAAp6DrTJmvXle/BvwOO6QYP2tOibMoGj5myjqkYZjo3jmndZqN5Up+doYU
Cr6DLQgxJgAWE6J0CSsr1zl67hAicWevL8xREYoaSb/gTcnranRHTZJjSI6Zj0s2
6FkLjBHtoT9IxKh45uPRkMUYuypcewQfkG/rXJsrZa7mkGxU8WlhAYidO85Ub9kG
GSUSXmwyY02l4nTeGu05PtiwuL+lfwxl3z/fiegQ27OE7a6x/JfXdEVY731BSbwk
wI6q2i82k7+JHFMTiZPdV83RxOaLpDFwS+MJ/pJC/de3aCDEK78MGQFm6jcOfKH/
AVdOmgmnL2XAz/ndiklSLnB0hYwiqFjabvaz94A4T4JySODl87qvZfxPe+FhQCOC
Kmbn5F5MhCSo6qzMUb2Ey4jUPpNMHAwKSn1jWloXvrtIvK/uEZn+sCGrg8cnwrDo
ZdkKdPRKMT89qUNWKMHgajwuPVvmjfeUFdIPp3lonD7cq35ml1FD+rjT7F/826up
7b7zlFLkFJB+uQ2H9acPDuHnUtRgqbmVaXyZk79yK8ah7pt32Uz0aG9i8ZInVlLN
XOvNqE14MfTJGkW6kHoDzcotCHJuGWcVLU9Oq4pXng8a44keIK5PcjvldGMWI/tG
pcAWlWLVJ29p3EakjceddfLNc/krZZEbcR5KqMIYtdqdkyNkincFfYdOzt90yvOl
2KUOTA7UhZJnJqSiRRzLU5IWXPKWwHA/PVOi/BHtlbFM+yWh6p4vihob3TBoxnd/
EINtq91UqBzbyEz7jf4dojN4xAXHn6Ef4Vk6RzDri8KdCT3qul99y2LXi6kAFpn7
lfuIA7D4JRsLhzIOPvoM3aEy3WCx2rbIo7tYUg+GccIX5J5hg6NVSnIYP5CbRtm9
PQsWDcl67jAuhTA279gKQkVXiL3Ocpeh+A1E1bVXkdvvtNYnFJTS0/4tRiPS28Bv
oRuGkHFnK+gWRD62PE7CS7R7vzP7AoU54GGNZJyWdC23PcBkqtqv05k2JV6931R9
o4fn6qy3k/rtMgZ9ClsXA0EucQzsxWeBdxitNLYtArXdwUzCSmLg/yo1NoJCVa++
zchqegQpEsTynoVmyYI6a7SaSsqjLbRM+lV5xrotrHN9sA6L4t6NqOOoZWls5Xps
I3ICgA6wPZC205MktAu3UTowCeTFB0ck+RK67kJGkAYHnCvetmVPyVZokADKjCI5
47eDZxTlkvkRGZtU94qD7Muue7bnRMrKClOjW6MCKcX4bdXcS9Je1eIq1/mp7nHy
Tp353jjsmVII6sHALDFg0+2DhUfjXvKxojzhnSQ00nt7aGqvK9FarnYIuKVc6ucZ
Nhzasy6HZmP/pigERav4s1AQjTMkhpuOjiiMoEDPPhKOo9zhKw9x1fQ/aIYc2T8e
yf6m/v34VtMJgEWypa0IRZdlllAPzRPSPKDVg9EletYquTrjaIMSNiep79PtrP3A
+O/SS9IHJslcRTAaDw9woThlCdpBO7nS2Tjc/j9KGsj7V24yYgEumQiTBSq1BsA/
YPL/nvVoTkSau/vIKZvk7L6XhbTtPUviTDePE/2hp7tI4bjFhBF3XKvH0TfGQ44S
FLkQ7kIhDESJfMWMu2uuhyiLPuNM5hXQj9TwA3dGSN7jJkBr3Y09LQTIDkltsdr2
5qC/EJsWMppwgeQ2fqJ3uLydYBf1malOPd+oG4KkcV5W9fQ2LVODzzab5Fw4wAXX
rtHosUueqpQJ4rNjqKHbX19ZkaOdygzdrUYiCxiDxN8ipM3EHk+rsitckTZ9ZhuK
Qi9PvAzgetDuX8AHYwLrTQ+EB58GM1KD+PeqrD2XOqBV0XUk8r2F3dvm20TD38Pp
5YS7YNa/QvnyH7woRnCxZvQgW09tO3L2XO8W0JqXAW/85mCVbjZBO8Vs7kKGSrqN
bhvif6ivrFE2RDrj+TwVCQ/D2FjJLEXchMYbiDC2RSttRsyIeWjXnaCeU9InH1Th
reGPF2t8OIAh2Hukdzga81n2kS57bwx/U4jOr9uIVSbnCcvrGhDfDUKB0dcw3GjG
p3nJf2ZNvf7DkYoNtH2/4NcFs08w6VBD4jcrWAwLnIxKpq0NANHg/bvRnC0+fPcD
vGdJ/WrfRjb/Z4GW+WFAwJT2sl8lgKMctHbXx7o85mteMnJvZDWUOWnth8a4kwNQ
akOEbzkpHJatRLsBACkijoTnXKxIUsnsFDoLqCeFupWBhKsklcWm0H8xZfUOdnDR
iFY75oBuKehnJCGdP5zB/Rw1kD6dsJRFrnz3YK0DE+xyz1YHcobpjU+s5v0okyXH
HvwYB5L4cHLUK2+k/5goNnsm6Q7df/gPq0U9GOmrzV547Kb4wdiqYBHTyo2cbRzg
BMy+nTzevSWM4HBJuQmdZbsBmPE3TX2VC9pJ30MK8WCb+0GFgC5uCYiIEK9Zr7tW
aZrk508Drgbvu2ef5gdHBRO5LKqVL/Wi6w0qKz6VX582wywDtA7yoLKvAoK1wyf7
3iUq+pBGtJ+iqun5uEh4mh9HEIJT8pjRjiuoG3fBTR0U4mnHNSsNU/Ceb7eJSLTb
h17AIOIDSrcMozKtyOAqbcGGq+I28c3TR8gFxIpuKJVrm3nh0jI6ECNIK1UNjNaO
SJ4PXCajaCNCroaDjnZ/ucLeROD25Ufe+fQxR9XHhcScmbGpzKwoRAIxgff+F2+0
o2/DHnJYFqSnttLwNYI32xnwNDnnOY0gCHshdeUKW6yUAovx1BIJTeiG1kqd/0WB
uI1MTVIoop6MdTTUD3hv5PXAXyhdiSwPJOcfXstxK3vQGJ81Zev0tMVTlVncyg5+
u4u4I+ulJrdzAhzBi0hbmWs4LtyBTABQ+eCVlBvH2fd6qTGApwAiRyEffAbvXDsJ
hm4Ynn19hkWejL9KcVpONOTTUNJQD3vhQfkoy2RcL7X8w7wBoj3wzSb0VRH9+qtO
3lGFsiM0NJmzAa/snOrhEakM3Njmv0uhxM2cUC92G4Tmp1NjGZ2N6IcbC8bsUN5i
22JJKvbrAs5e1dcIjna7hxpkRCev9jEQLBuffp41t143lO0umVb0yJCpQak9rUCe
9qQn2msL4YRSM2sEhgzbvNqC3Q6y6/0CnlsSh0aeMoypX5uwG510pR+T3evIrveu
qVhf0rd2NRg2cMgCl/Ys4qrB8DJxlGdgeH4BM7I10vFT9eW96xUGNHtZFVwOQz1h
VF+7roNDgs0i4JEP8jwpHYImP7gaJrEx6sUzJ/jX9B0/W+oHVbA/mrAj6Cks9tpV
M8+8259UJKRBXzpxEDeNWoPAa0ldzyttBzvL/BI7DernJUO3RdQAg+hDkFpyzkvI
kgI66rDbUChgf4kqBbjKy+YpBy69qtzsoW1xDFhnOXimQ1UvnQdCEqPTt+R1zzyR
J8Z8mmPmR7w5m0lsHqr6LEL3dXB2IfNm40aa+pNoxCvYuOvkIl3GfxeeVF0ub/5F
ntTJWpQXy6HugFEHr1XIFPK3ZhT7I5umGE61svVAeIj/ZsRDIuZdag2BFRlmiza7
lDCDTqh/Mqx8X1h7qaB3U5ODPpqagaWnhYSzR+DaUsRaO7X/y9ocvG/h/RzKxmaL
gXzCu05kO1lADy6y3fAj2Ef1+yclFF0tuPnS6UhcBDLSBoAHRuSsfTwBKCdkmrGY
J4G5aYQCx+6/Ro8HNfa4jhZlMhY2HP0GZ0pjR88sh4LIuj0QMpVIQR26OJ4RdNTz
+/WnR/grWg3AtlsqmB3hhBDo1zIsEsb6FMbfH1+0GuOzwra7FsG/oetRuOua6hvp
sYLc4A0ONZ7bFIcZAUCzK1W8GRc/vcCzXgrsRH5YtRU5bylwkyzHTsn99GLus+Nf
78QuFK70/fYhUQkR8rmNx76XKB8+tsMr1FKbHZijFieGWCukghIkwBgv6DT4pMtb
wjdfKSGnSCRaUgz1Y7NkQfx7jol7x0t+WfBzZnubJyqSR57wSrh46sAvjtG9WDuy
k3fOHUWRbYrMw1r5YBUgh74ySt6VpzWAtHtKl+2MfkSHk5wkag8i4FvOUQm5aEEJ
o0dad3x3VEjR5wO8th9frjuzCLJwlPEXCCkqUsz/IiVNlQ1iWuhU6Rq7BfoRa+2M
d12XY6dIHuGv7izbGCJM/En/E4Tyr4R20F28wm3I5jUYH4m4BvmTroMiALFZ7nZb
PW5S5L2h98fcNbhO5/uqeQGdybdgEJ2Z5StcRFmvCTElnpetumuEhy9BAMMlIVTZ
/Aq2lWgDEx8bHDZBi3JofyX84AIMj3yk/qz52IlMJOINqknr1g2h4xKJ1Y3E/RIm
qh56rKcg2JRiY0mgSAS4ez61/SJVXpVwJEya4QKvZ+FARdCwdPbPHfMhyu9oUbca
lZE6wi7mSKwGauI4rDi6q0VpDOJthdkDDOLPI7AR9vow0uhZn6A8ofdUl1eJlZ8c
3QiUc8iaw4fM5fOj0jxRAoVxXnvJ8bXUWnwoUzWKJB1o6o99PwvSU0M6WkwmUEg0
JiwHTWE1vwfO/CFaqzAMulQBVWSYJVQ065vgiJ5juqdN5TxiLeu/P0yqzE2k3f50
UOZ6JiK2uutqyKw/qFSDjrp3jcmx/tD/fx0q/UPQ+rt9oCs8ygTalQthzLTFGE4M
v7cgQIk/3yEleQ711kjsx82+h4x/zSC0R6IgAg9YzriRWFdGOzpiJxtOUMu7NSb7
iJEYyHRg4lWOkKL37/T3YuBDOG9qUaR6ze5JVlJbM8Wcgg35PDiDSbmyrAn0eXkP
HoghgVnb+J8fznJCjN6Li+oGwAPWKPCKaNbm8G2SVA7V/fc8bgfcMJLUFU/kg4SB
rHe/s45zF2GFO+EBIiXU12R2d2qfWBs8oF1gqKf5tZcBBIi7p6dfodAK9AVi1y3F
h3lEI2Z463L3PSo3JB1PF1kiDtIyEJnKdQxV0wvO6haAR8dJcPIwyihWRhTyPqYP
wgv/hkONBWUIXprPyKgOjORlOypsbsR0mlMTLyAq9L+L3t7MJ7xXBQ2d6SkxN7an
c3cYrvTCang33xJN9mQlmkwN3xTjmPdQoAkhAqYZrELdr6ogVBiPMzlxMpLFn/aq
gjdOETQmEhRXR/t+pvBise3wQFMxnJ6N289rb/ksFJww7frfr4X/Jlt0Q4RDxrCi
MO6lOraPADx7hlgHWBAxyUuvnsVS1G2spraC8Vykk+p4y9a/gCMd7Ovdu/aFgcva
kXu54UUqq/bWryznVZ00TFib4cem503SLOSDaqt6++abozn5WTjym2Xre7pJnb23
s8iOU5+LAo3pPXXhLlB0yetkgcQIXBfjmj4J6CAGofM/9+XUioVQNJjod7UCYPnV
RsK6geFtTgP2KG+GnY4X2Z1k4wmg0DRKRk4gk0cAAex3ufTq9D54dV8tsnd5ZMgK
ftkgYdBz9R0ciQXF3cx84ODo1+IBBk6ayjXN3BsaI8310fmlp70pEUxHqEOVr2a2
HoaXxxhKcDXWCKU3XR2qAX7gjNMkNrc2fNxsaJuGLuy73Fs0zaRKdJV3b2xxRb7L
FVToKzsMe5fN1Wq3YjLJx1U3FQLfy8JB2tozQjK2UL/apusjT0UbJsmGxEJhP3HS
ZvU8z/xkkkVPpuU6HxUgct07YhP2AEPd7eu9VYse/f3PB8mGAYCAe3EAU5xxVA35
C1sNXINV8ILuqwEeExTlhC9/lfqnNM1HVdvtXIOletsJHkQQ+hfNBrwH0CcCTep3
yzcNOtjXZ9Xdzqn70SdzmdITqYOrlgyxsswFJrx7j3RhrPOEgmh0F9NrQej7/UVG
ELg9OpYtFAbzyNrgqpwuOAoZawilpaIjgaS0jZKQPI+bK+0Kr3QIH72X7sjykfts
X/ROg4Rs78rO96RRYO2bkB9+9rlFwJalUxUXfGfl/0CT1kmhAXei4HC4raxMlpe6
bb72JiLeOnnV8XUnBD0qq0XhS8iAvvdhixsmLzbwYhuwRMhBZePgh2eTkPJxPwIF
KQhgwMHx+sTW6Nhk9nmoa66Lw6cNtxWl9OtbYO25ohaOYHccTNYH8rUaR/zg2nOK
N8Qga159te1Ku3AiM+b+VNTA/iuX8zTFnFNXm8YgTDJLcPgPTD+xj1BghuuyrN+J
B/DsGLbCZUm7Sjq5vC0gdgyvvKpJLLLDCeTLRyWFp9sjKtH084kt9New/7EV9ldJ
8o6BSP8+p2RrYZXpSkMp9Fa0VLPjuS23hyhGl2e0p18aNhV/lY9c1BW8Vph3NpVy
37vbLIkNNIv10qrISH5p3A4vMuiJZBmKkiYkqLqMpKVMbTzL7gz3LohZaOmicYgB
K2ByFehNhQhYwzjcZ4cOgQy2P5yN57lUFYeHw78K4dzWWNlHLh+WIEmC7iXMFRot
mF6/rnevv+PkW8fWFsH6Ox0Bn8JssalRNFORDG3TSJmF0n1NwWpqia2Kn02govrK
vWRSLjsytZPHrAn3yvMFkHr4hbV/IL4/KIxFAiHpLMY+Nat2wqskXOIWOTYXCyKF
VM0YTN4VwvDbv6sODs/ZhMCtWPo8hA2qjUnVMC5vEtF/szKCq3DB5EIpjag/PJ/z
xEcbMgFTLSNbTstLtJb73LiZL2/M5jYnAJLiZNoA+6tmu3Fq++XArlArhbARtubb
p/Ws2r0lcB7KaTqUDRTpU0tLekaA+ttqbSetk9FTbi6W+3D1TWzSKKK+lxfGaf8s
HCUhY9qpoyVTqHBDc9To1JqGVvi0XZDbW4wfFLO57llC8X2JQc9vrm1ird6LlJA0
PnvXrg8415urN4yO5NAfbeDa11BJgqviwBfRRqQA4Yr0xRarMfnn4V2+JmPN727P
rOXexlbhnLIWYYA2CgflZf83Pqvt1PW7wvIxPt68vTQ6kaP+oRixpMEoCV61/T4J
KImm23e+DmE5h5Hscl1lSZPYuUFQzTqA3RNIoyM+ooYe6V6munpHQbdJOHH3cLCD
2ytHYzbT8nZto4ImizBONG8Fg/aPow8g4NE+pBIr09hrirrGYxB0s4lrnDuCHeO9
Tr7L290ypoN/yC8V5XVbJgj7IRbwSyesM4zSuX1wSMCP19V+sNLRXjGGHVjrEdmz
P/8KFWx8sQcVYXTqsXv8MjSXSO1kf54BWa8P0gNOptcJ4N4XMmLpi0HJGKvucHcO
KRXJLFNXgqIORQZ8NUD4Z0GOVLB/rfk4NlXTpBam2SAri5Y2n4lZTSst7D9k01S7
x0C63MmXlwkVMNXHRyCeorO8evXqCYmUCSeADso8r0nxVYFI95GodExlfwlYIbK8
OMztS9cYZ2/rgh4xJUAyUmaLrWlUuxWPgLGCqANj+GOZfdIVbA6EUqCcpZiNJBSl
/lzJ/8rMUoKMD6RqhehZam0SvJ1usRwecr96xum0DhEFZyCRuaoDhg6XpAKEoIKu
1muoCQEfLJ+C1zYK1eNMam+JPz7yBRe3TvMthQDN5Yf7Eo260yBYCgJotvSL6uzZ
GZ0ENP4UNlIpluSkv6ELo/giVrUsDN0EaNNnQPTLZwkbILdny0XBuAXbR0jv2dcV
ZclRniOBJSlWywKV0vbWsDX6fCCooV8/7Iif4ABfeYdfTHG64/nNd5gE02YDOD0U
hN5e+FLswEpskXezLrBrbqfanA2ELOVzmWIlkMYxmOmP/9P1HY73cK1vbWAW44vB
/jFyLVU+JgfZGWJzaFxBUGnEl5h2I0rsqTecBZlv+ZX80q370DdH5m0zHLzlE5jc
qO0jNRlU270nT6mSIpiScZ5truCLsqVc7Sz/qP+XYtYD3lC9aAgaJpwQPdcB4Vdj
+ty/aAY9TQHyI862hYbGOyURIYhpLIQRYykhWUzj6HrHT/Nm0jU+W/+lmgRNxUz+
ccebWtusDMnZ2G+QJHb31bIc5tcb6tzZfbDnZoBtEi4YlHjxvg8/j/kEEmkUcDSm
+d1tP/Bnv00aWjRVMOPasU45GzsaQtj0dqq73RjDJ32efTMw5NpzZL1qHOiGh3Im
F8xLyoMwYnY7/moMWF1q5M6IxeLvWua35Guw5VVMIwrnS84eSkPnmnPd93SL4agy
o3FQaGIPGzAaDT7qwTOWDhtKP4abMPDeBS1keL6whEvSW+i8hFuTsqVFMFuAGrVs
A1Mtg8UQfp0SYIStBpv8asByfekM92u3dB0JZV6CM+1WN+yrj/XZGqv7p6wWamq3
lZtMbY822dWLGnPld174VipSTdbU7RzSSLwNQhvsF4SHP/evqxVPAWi1ECfWvqjk
3febH/90PbiFlhZdJu3On+R/i5z1RYe8Ax+IL1QbNPg6l7MenSWam++qZMktoLac
YaQ8PhikaLp5zm68d5HiMNCaWjFHxGxb7aX/eJ+/nk55wy2BsgT8dmFh8VV+1AGY
mumx6ZfAzJ2a5Opa9Ed2G/o3Kp9PRlDSOaAToF6DsZrPm9AsEvD9X3lhvIkVBNoo
qyxbtGPlmBNwOzQDrxQ+zwncboYCrd2Vsc5xG8a3FwN4Mt9IMVgDxZgtCkqzSX9d
JPhnMMYd73Et5ehMsiKhW5MKae7mRx690a9SYyk00geS0W+HOM/5reOQTwJ1RTkO
ZqQJeOLCHBpCx/YpejVFkaM/N5s/aF2P7AawPGdY7jQVMa8PrhIyECWuznjXpBES
u6qMEwRVibYNX78Dg0ivTffQ1JPbhHlwScxYdAi9ZDaKzlOBbs+asqn6pHBs52OP
6MxHUS5XLxN/1ZfD9vr38EbTpvcWopTxhnY9S4QZPBZ2yCKphRejPLkrflfPRJtR
HjLKvAjdlQdDC3CRvn+sezXI5qp2G74y+TmyaLvPqmxGd56T/uigml6bCfGzGTdB
kCKx7frjNawYTBeSvnaWtP2gQXWWGAri2SdToyxH109nsbMoUsf24Nb0yjr2GKqN
u1qJwhef3U9E/4P1JknIgPwX9HqSS9GK1V5NqQhCWoGFutdwbM75vdKa/oOAcirT
TmcKITeaKU3KQoNdKnelnfXE3mZie0HIA/oQ7pGzwOkDsEHRGP0buqWqF78m9KEL
uvdncKr0VL04t3k7lqCBuf7lo63kmJIpg06HTBFujGtyYfCoS84D+E56y01u+3Ty
63YviwZlXAH+S79gtinBVzb+QIItP/vQCIgnhMlW7Mk1SB6UAK5UhZtjZR215Ywa
wgFG6EfrG8Z9ghv2LbC3RslwScUpo7+dVTaW3pu8UJIBFiatWCyEJG8nXS+nx/MN
HcoppGvLyN5M3V60Qhr7ul+b2ZNigJmr7inAmaXfcnL+L0/JabCi6YEU5Qk+py/w
N+RiTO2dbreyuQ0CB/HT3NtamTYtFCl3GFQmmfKrl3uYc+73ZuLhMNTZ65/aXW6R
RBSoPApoNKSZ8ffIP14YAUTU3e8YBsvO26z1ZK6Yklgvv9rQJPeePnWBx/fK+8YX
5oTGuqzEF2VvNMriyH6LVbz1I2IlsGZAfcKILwXQmBZEtZgXg9TKJmr2ok6rrfuW
Y3tPfX2ydelrWYNtKAe11qqP+BkJ7fV9Erpf9icgC17+PuW75D1NpJ23p2df3FmY
tYXQ1XD7O+Z9dybpEOZrzArN1iSHg3buxYGq+EF/Qz+UGJf388jdIz5kWusXWvlx
1wnvPnhf6K4BnTcT56cRNqao0FTkrQbbi6EkInrxGuVcBaE78b1QazIvc4Tyh/oq
Q7X7ia9CetXYMBLjdAANUA==
`pragma protect end_protected
