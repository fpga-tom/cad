// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:38 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Fksv5sCo+mlriCtnVKVIHiIXnue1I93X99WY4gYhMYlVUb5FJ8zQkUAZbRwZgceG
gGqOuK6kvJSfD00lFJ7I/GR/GRbOie0ckJ8Eo/7/kpDPQHPzR6QGKrloDMOtpf9s
rFRepXQsYmftsOsTh/oz9VqenwWWFYzbv3DXyIuojUU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11488)
vbJYr99HiTJjsetH4hQPe9hJdbTPQxk0x1qt2BkPeLPMitF+XB6SvY5sc0nBqjj7
llgA5nPu/GFkAXR9IFaMaBvhhF9K6+wC55pLt/YWmJduYlsDZg2KOzCWmTZdKJUQ
oZwoN8cuDRWqt6IUdxvFshY7IfsYyknw13XDO0hmAH93nzt7BJrVUwsEmCYf1ntC
2ll/bL7BSzCGIHj2KUP1zA+M3Mn7Knv/9HQFpKUbDyCgalPQ4cMplQcKkFztrkQZ
GF1/Qi1ekgKr2TqsxBJVUPTS7UqMxvQyVgEtfzTyfKMPH6Ug9jJuclhQQZg1mYJg
EQwSYNpbvy3fY6bdPVHq+OOTL9w7BVxFtIbTdhnHc78vsKdvr7PDUN4xSG3Yjpdm
mwZN+6lDUIChd2G+K39Hd5fYfa9CDTx4pmecryUYWUvqrShsA6GX9xVPOtJy01mP
EOGxl03NWVyw1GRyUXmbg0h58qibZaUxCtNgNmZ8QGj5pvmGhDqvDx0uOSUZQlFh
QUmCRKmjiuZFHVhWRUYwkRmomxvMniZiCpx9hPW2HNvonzf2hdnbn8l+FfE4KI+6
vQrZQ6abrYS8j9iZEGOYSSaB1GTo2D7+GHAXogwYWalJHyT11ggiHJzJgb9pq4Ue
vyTdw3yXIjXCYQ+H7cD78Xyz5nrbSkIaEKBw85rmR9ZhmLIX5dGdFF2a1p0nj+NP
MOW5dOU3A5lB0uqHWP1pwrG3HxE91cGIZDemQ+A30/ZKLbToTur/r3IbaGlMOFuh
pbWy8YiGcUAl+YZY99K6DBwMrA4byCXw7CW221rU0GGuw9eeX8o18ucTutbzZtdZ
THcXJTYgB4vI/osXjph7Wp8oJqvhtFJZhbgxQeaIGHXUxBTCHWeUnKTGnEPbSpVb
acBnjlxbTOAIdPW6/OrPDytsdH1QV3Lf29+gDFS78niI949xAcdcpZAwVzRxmbMg
XRKzpRY4k8CwtGxIrdfOhzRZQzjUTcw77ntHCWYjorPiLTcdv+PgTnrs6sVL5FnD
R4HknySRN1MYcDZ6bORkoHPHZ8Xy3pxF6Fyy0BnnYTI7NbnrG8O8PAfY+S2asyKS
32cvnyteDr0xB9wg6Tc74aVOY90/BJPO1hyPYL5+4ehTf1vjb9LhpEq36v9mckBm
CHaezXiI+oAF9Xg+U4xlXzNZeQWjnpVwOMUulL6EBbfTBbPJ0Hy7CjCeSvTZeG3X
Rf15Wo9a71RyNkGvplj1nMenJ9yxCIR0mvnwguS4wXE3Mz7vYA9rI+y3ZZUT3j8a
pPt/ySE81VIyrY8jFTT1JIxRgEAAYy57K1n8q2UHjdkY8u5WZtg97ICllVOWY3OL
RmQ1YajTcqwm05MjjMn56e6N7zbp8JZfq6ovB0mGlrvNbBzFb4vOl5aBGrK+deiT
DEJ4O9S3R4rRXlbAtM3EmlgH3cr12oh+G3ZbuIYiPw9Dp48Nl+qUSR8bBLo3lh7B
mHdmtANoEAewVXjEkR/d3axN9NjxaLocM/CWOW7/P6dEzlKMPs0+ICproB3K21n6
OYB4ioeqM/IT48guhyCM32YBPlrK9+zNkuVgP7D0ZEgS5oUB0bqKO5bwdvt+kE8J
dI2VHFdBhjUqHaO+szJHSPtLt0X3IXTEXReSE2QTs0AMn3blOEvKRgX4iSy+n3yc
fVuNLlMGhbAeh2n7NZBi12LcUgjYv6lqy6nU2C/dflKc07wzLcwJ4oLCW4KJG7iz
1QkiSh5FdZWZZoEzWsaNz9sQBUxCwPPovr6jjSHeCVrFIV631EKkwZ9DY+3r6tlo
GjGmEHseb1k35PwrctfKvZgESLHyJVg/uZBzKo1hR58v7KFMcCgd8MxdVWNznRUj
jHCHcDiaPubShEaW5BwOSKs4qGZbyWAf5GTr6q4C2hNZKrDcQTtVt6pc2oysrC5l
le+HXV2oZ+ZgVzX30DvYQ3+moMmO/JbvOABk+a5VtEDWg3lbH2LJNJWcUxR3zGIg
NNJxYrPT1U215i2GlKz6CD6kbuGd4OtC70owQnoMzSsXdvtTFulDgSDKYTYCzr7p
c8W0ur0suBsmr05O018mx0LbGpdzDTmndohhjCizCzSKoK4eIrGmbiv7hGTaeeZ/
ICuKy8Hcqrbbp7kvJMUR9UF6Y2aOAVf0Q2z0nKSiDZZohrBYVFA7gZImi8qDFI/F
fjl9WR39QrMVuZzwrUfsVgCZVIs81TiZbSSRuM0Vy1r2sRO4PSJ8WsA9zl57mcDT
P9STszFtq5F4vYshVHMIUde7jtkeB3EoZUXyqMXrV+/EzxLD2qBPbe5QBTzZIgAS
ehPqHnbyZDiVSMF6WjrqvVXoDxUQBgSRVbjeN2iZYS5o8z6fWKqSzHoKssMC3y/z
OEC6GKTkizKzDhEpXjft7yZgdwhoKUuFUAa3Lmd/48+dPil2HoreOsyAKhdymfts
1smQ6PI+iXZSJqULeMWx3wSchbYGu6kQVDLGEincMRri0KViS3HUgherf4QYHgvk
9jYxDYnFKHpMizY2TbezXfJsrx7Wr+rikEUkOvshL5ex9LaNfyKvp3RV1ABunnXE
md7IEmZw+ileDtiNRboCF4h6ivXbQIuyQslctP0S2GKe+ICiXZ+OeKGa9OX0thvw
m8nh4518g0TOLgEieHYZ0jZYrgzovXmvAcLLTCYkNLJduWkBMBT7G9vqoXN07cKY
x9RbtqC5GKjXXTbHae6ShIjlhnmqV8fr+y+hewtEWpCYJQRMB1mtt1MV7WKIJ2Ua
ADlLgd+g2loId85Ln2YjsJjLKVHOJeajTpvlK/tqm4tppg394imMinR6Fm5aQxMm
3CPieK10lfZ7EvlFdAgz9iJB44RqBK1vXFvOgxCDz24nYVEiUiPNcRXp8ITcHVs8
Ee38RKSR0JLvIgSU2MH2eibwxhAfd+a3OH1pLP9z3UXpipTJFqH1wMWEDh5Ik0R9
2YzbpuePwvt5APEBLAe3Pf6ExFGhqh1P4he6LPU3EF+Rf+vBt8n3yIsv3hwCy+YU
j/m6b1S/pYMkC/ynQX/Y3FeRzrePWla1SQMkfPaaiPyIsgsDutWwsq/bQg54BPUq
Mp8Dyqr2LT9OTd+knlSfx0+9lAWVF+XXF1BLgshJyK2LWCk2IH94VS9dj4hpUGto
eCNwYSxMOY6/OpMA0iXayWg2k2RIE/T9HhEt3mOG31Tsl1PWAO8UblEgmfeofNtL
u7vmNzSYAlRVKGEE6MNUTa0VfrgrCt/jwtpponkevrtvqqqY4j78wl+BipRdYBT0
YHkjEJdGr0ApxjHMcmoeJsQ7rZ4P/eTDgOfT+VugCV77KBF+JOzfVPjwexW0vT98
BJHaaAP9QXAR/Xg+OF58DbDAIMtO+nxPqHcbfFgcMsAGyBZ/A1Mhst0wPnZhu3LO
l58FUC0IR7/sJz3TZouvbqgrmg47eyw2g+clJpuUwRLGr8uJtF38sYE8RXC3+ltg
fVI2GSW7xWD8goY98wwN+2oRjNgZkAGaq2V2tQ9h0Wkqv1W6EZ/E2kGRhh7e4E6X
B8HF8vuItNCbNYJGAKyBluVNwZJAEcHbgCgKGsEQnSuWjdyfdlrFXlgkQXQrW26Y
+yLExzdM6ZDwC06eXfTZ7iGbSxxyVImafr15qLVeRybri8GRtwsHFuCT4iFStOVU
u625Ku7hgTQ7P5ZiScVF+nmebmxf8XSDfV5/GzcV/H0ZmM2gg6r5Y17tu1+Y8Voc
KTMW28lyDGxM4yU35PRBgap2/AO/U+OFCl6IdSFT8PugH0U7CgaqLixtMj+O2U3W
jpLmzuGlwAw7qSv9JDu2qrhKBRevoLvTojqsK3hdijhBVapCZUFP/2ijtu+qNB2y
0XEBfqT3nXu92NPHcvWpzx5PClofaYoEVhbcw+rZ208lbscTAfN8oJ3DguSXHVjZ
ZFGOCYEHOB9/k5yALQUcfpV4GDEBFxEu4dLireKtC6BVI06oCsraSdhJMWZoh/98
7AGATyRpOLyKmiQ6mJGsIXQYoWlQuro4n0EWAyQv6+Aa5qFTwWUYPKrfBTVvdjSk
1tltU2iSwANzxuQukdYQGzhx1w0BbsEYzMwbDB/ByHFRElrSsDlVrYXDD15MUeyp
4J23KKEtXF/9SxXpIKzHqo9dEYZ9Gzkfxtd4JxgkgijC06U3ljbM0vZ2b4Hm5g/C
3jheKm97f6F5rHM0Zrt4ACmvFVvy3mSwW/1YK0Z7nNv32eKi+fFrgXi0582CCXip
OKC9N6FRxhjArZeTI9C/ZbMLXpJRcWRgL7Pg9nLIbWR8Jp+VTQvHDgyCnTagpPIc
F4/aa8mgq8cmrxGoMV3Y906ZVlbmNxp/IO0OWrPRmVdfG5u8iL2nO1FIQ85sB1q9
MuXpijJlgumwTzb0rEXO757A85W1chUY6ro96wFtFPiIIgcuAl/W6nBqGP4OKyBU
aM1fdZ++QNnsCO2cvepniLPr5Clm0CjtwJmJe/HcYBQ0UQ1W5JkuLFQNvUTQVVNO
kpx+UkjT7XWDnDu9ajVsIGm0F9vVGRbxJEgfd6iZjegHwRfOys8csqA4djSl3A4b
K07h4LKYCdrftjVkgBxm1U3a06QRrloUIyfkLc+iuBAh7lBl7SyF8ZHfjjvgk2FA
ZluV9sRlQV3T93UZ1FfajaeYd7hCOWpukOBc0MAgtjDZfxPYUeK/CRUHD4PQCiWQ
N5LTswoDas3bXhOzXxduOCstWKqgOOwIiZCUGSxO0KoVBLpS/8GgcVIwkvVzyiiS
n5gVpPCZTPchpimonVbncUjZh1vkKJ6s0jmtwwmqJrp4EEGRxi3ebUC/EfToWSoS
Wec5UTVGWISmlNpFDmt1NATV25iJfp7UF4YI1Jvp6OAC8g5jJmEmM+Zqkv3fhkgy
/qG35VScUIuCjzmGKTj6qrsRIMv0t1an803GO60cMy3wblQGTpxW6T5WUSXQHBHL
pUsrRalS8cJHEaDb3AcIsKMrGVjXeevGe4SdGCnSWzch6kkuesg2vG0zdDIrC1gg
A4XGFUvxE/VXfG3SE24AL+pkq397ZIFajTF5MiFCw3Nua2OPtt2DI8u3Iyw6sJPn
jgdNWdmoOEmmLJRbVnQ0gCLQfDj8jQ9ZTLjYtiJueQ2Yw927k7IzLBEq8l3eK2Kz
YWJT37xyfY2x8dyz4wjYETuWeooiFZT6mQWed0W8BFwzIusEI8M5o37NbbBTpmnG
3A65OtSqVnMqgLTbCyeD/4SVLnro+oDn/F7GaEcfj0HHUih9ZxNftjkkYTwQD3UV
wk+fjBNdA3n+hXEi2s2bbtGl+jXiw80OtSr7zrr5xa0KpAPHiIQfXLRAvF+pQoZ0
asUXgnxw5PbJdfZNnczAEyYM4Uf0ZDnniN6KTVCwQb5n5UaGTcd3k3QBrW5Y5nmC
BoDq7EvnBhvVTjnhPr+igqKy72B8uqAPXTT7VuFex/BazhEB2l13UX4cKsFVShnw
NumUP5olxRPVVt/ocwC4NpPGjgZaP0GMUN/AetrS4NxZ1+vASKNe56xwYVyYsaTm
odr2hIU+lJx++Y9gP5alaZoRiaFmsYkHR7nInzttGEhQZLEJ2tdhOaip65PAX9yX
J9L/mkQ4zOmw0idyX5D4MN4sRMiAzRKpJnhS/9ucy+wMT+RGdRiMLnZ0tWp/+ASy
dfaiB2aggO6ZkTbl9GpMpyKZhbIaj6Oa2fUB/Epx9zX5q+SkK/l64Tcq3o4OPBfS
snJvI79llJzhNz7FWFAscT8zEW1D9Boh3Q49eBb2grR8eFFoR4hPZ88lVfi+NK11
ontYkG+BSQgDHRKR4eeNd96CVP2kcPPrIPVwz8XrEkWQlvJsqB9Xgno0mD4M+eQz
WC5GH115GtR1RTykMTgfhmne/vZ56+o6nOrEhG6Ujs0R0dUL0sgJbB3VPhzNaYJd
JLvyWx3L3ku43xvNTAM6oSsnMj/qoP44wvMtTYIkK5makN5eDDxx58xuug4PqFkZ
E4Vs14yO7XYkOeFLewMH2BWM6QcSU5pnow6hQ7fyofJe4ozGPoCYQtZi0MiKDX+Y
YeKZ1h59GSwKJMQ4OnztwZC08A7tZIcS7DRgRAMZ5w+Rj/JeNpLa43oxof+EXuZR
+iBD00edME4B3Dd+xfz88MWzzKhy7MX4f52W8KIguuklb/Zs9xq4UKKCV9Mj8qxn
mhFKW77gtTjKtdKcOMaWz4kZHu/wvh/iklYef/Keg5sNmBRJxmUUznoZbH4w/B72
Mpvpvp7973aC/Wqe2jj9C+pbRJMMc5G0LZi2Hdo/mJNQ+SjYH5sYMtoBaI0shq9U
3qsltg4PMfwB7QSxJZemKr0LDdVplN4YNIvmUv5T1V37mgS3a2WVOXXWC64vFyrU
K+5Z8kCNew7Cnl5VARH01P0EQJXZO5TEJ1ZJXAHL9r1dcLLpa5w7GNb1ErbhupmS
3umFr+X2p1eG9lJBaK4MyFE4a3e1GPyV6Mz4XD2K9XUsCzgYVW1kNFbRX8x0nrqk
+xph4Bg99EDYdbD292PR98LxG/50JBU8STZCWJpXOvhxlM3nbhvcXqdvkIbtY56m
Y16uIoyEzEADvwwHd8bYBHey0xqjPLO91nwaoaUu91VHGdZz9QPKr4BAuF9Bw3iz
ZVk90jizdWZEE/26xDZeDbWpF18vIuyILR3B9Qypbd7/NW4hljjR0FUcqmtwOUHM
t1nsKFXVYF5Is0ipitWEUuxestyOhVfboBg/zvTwJyRkiRCyNhKGbbNF+Yl/VqAn
oHZd5prxOrJKATmSF7edjLOYzNTSmkAlEoVse5m5crkzetVrz/OO38cDVy1s43L9
GWt6HkhZm5E41/bPbGHO/fVvpcFihDAP2GYiV2XLKBb1ZaBsoOEummAqLIA91kHQ
S9g2yxsKayaq7AvrpAa4hiVa6piIQ2cPTKWglrMOeT/lyRrmIsSYn2K9yvWLz0tw
1nMe6DlU3sXMzdz257NvQz0tIkkFPPmouGEwKDaWJtl6IDoz0yF0gd7GMWWzG4RO
1tMEdL9RZVuU8L7FFNz8dxfaGNvdHTjvqkSAo9ffh2bbjlPtKA1Pd8mgetu1O9oc
LAvO01BDQuGLzPIfbDrLFmCi4cSVvr8tJgXSDTEHlw3K4PERdvUDCbh2EvAUC3N/
StPzMfsxdYP95FB49Qg/nZSV8V7JB8KkeO0B7NML6xOjbARfzUw7DiiUuk4uY/4c
j5faVFtCKyoZVH8V8jHpTxrgKI8XqLEIu/u9yOFvjbrefszyhpd24Cycs1DrSJBM
QXhcEPLkZJuLUf2jtTOA18EhDQ0KpmzLbz+nQBbxtHmY36xcMSRi3tXTFcHnYbar
G6rgGxSjSoaHTiyHShaQ95u1PnnOwIdThNzYuxgLkAztLpQ6dOQRU1qbooXtjFzB
6oFZsXG3qqgf3OgU0bQSBBATRrOp1/k5dMkNp676qhHMpOWVH6e1PaVKpE7aV/JM
+cadPzarnliyYhzKmC+Q+XMZ5ns2L22Nv/baRTaF74xV942LPREOaC9FHmLlw9eH
+yHlKIx8M9QPpYkJsA88XTG/4CvnW7F+QL3BQpr8DBNWCqQVuKQgP+8eCJNBwXRv
VpyMyJ5+tE1tO0hdkaIYTCuuXvvy4lhdqZf/ziI8SDcEzuiZv824BPcb+J8+Mczl
SUXcmiZPkuH/qa2TxQAqOuPXFqnvXGT9wYeawUDInN6tQiSoKeZXpjwAEyiD+6c3
A8g9uVaDjhV+sHcIZOR+WTcWWjmXdDFbfKxJrkFaahqFDuslz6Rkp2m1zvSkgnaE
o+Lua86p2vMRLG9eadWdquugzM8LWgZGVkvCUuDJwAG8YpinF2TRaRBDpVtAjEc9
StHS3GABf3SXIg656pjxhhwkknoQhKqhnFRMuZJMbKIn4P4b7Ux1crttvWIqkuJG
2ANl6xQxkD+tVcOdHrqkHI3jCDOrffkTJzZjr/OfvZ2tygQ0/L6r263uRqib3Kt0
nl8hkHmeTBsYO3sLz6gaIPMjqBEJRNfnXQBc8JXNfKTMNpMiWKpF7PDznOl6ht/o
HR1CYefiKZNXh97HQH6Xkersymvoftoq4n9Kq3dWmjxkJWIJLrl/1wWlMKnq0nLH
JTPJiwRb+97JnRkTbHI89n6i8onfytSU8GIclb1j/3mXGSLFde8HcqOzDnYcfhHf
zHvGzTesZxcus3wm4quBzG582hyjaE6CgA9QaiJLVNUYF+7k8JpUMcvdg4IE9HGS
BB5tdjGsV8vrQq4xbwCgLLbKcU2N5SklhHeTUZqPBfYy6Jnffk2fkVZgAtDRNBDU
TcSoetcy/O+CJQYCdYzmzMrpuYZr4OASsKHG5v9i5nzwHtT7wPd4QmGwCcjOHiOx
GIc73wqhGXbdgToVTFZ33K14b8jwUsUWJXfTGZEtX9seJlye98xWIaStOHlCS1sM
ZO+9KTBjKRb5ThIVhc3IC3eN2MotwAAYF8xvf32offqjjLSw4ehkds1klzGr7O7Y
08tEcYXSuRv7v5QbuK2uLdwrp0zm8PCJXxPDoxLTRsdmS/Selb92AB35M5539o8o
+MBBrp8QWWsAd8l7bNwuCbjQraVvQtIIMEcs/V/EP3j0ehrYbJO1EbRUS1TAM9Z/
Brx7oWft7cwhmY03p5c2bTpD77s/xORh5YKyF5UfsvFF5ceVgyl2GL8hTQumHwyb
sqnuLBnncMKFE/FNNTwsyseh7jOOPCohPFl6e/5TLdWGeLZAiYI0jTSG/fDJjMXY
+DCZ053YFkEIItYpA8GaX2pGz91Z6w7+ju3s1p+jWiCLO72FznHMKK3uccsmNCts
xsrn9ldDugaEkXCtgmTNJxJHVURpMVmyhvyWYGKPOj1uvQNcoieuNezY8mc+tv44
t1i5hpILUYWY6pdoCk6nQMBlK80G3iZtfasl46dpY3wAs6JbVHxnb85R2iNwr/G7
PSw3Gv1P+jye5aoYF9UtqrJ87ZmdxY9L8VdErNlayzDOGmY0oF0PhL8XpF8TukYu
TJzHXc1FCwrUZr122tWWaRo9FUcZVJfjRH5OM1BjsXSGzwW1OY/2aqBtPpWfuZQC
N9XKTOxS1iTOTivAD0eClcPezurt5XqwMA5Hq4GWIrZFIDTC17hO2YCUcuQu8iyC
r6wsG9PUv//ZaJ6zQYxruAT0QGSvYX9ipMgBwnubSpzX4EcUsueVR3Nr9q/8La4B
ZvBcaFGtjf8AwKwyODFI1+yxbaKNI+qTN3l1CEfZDDAjxSCeQQUCAqIwoI+Fj62H
rP5OIxyPJlMnabW3je9+mIrIOJj/abZ4KqNkCHccD1jHrlOaVgZ9E/vymSSQRD9T
C5g5RCYaFoJ7tm2Ttnnp7BmHH8ewmHaeHpfeidZZUtehkzerUD6FlWIY1CJYdIUg
mRXhXq/a9smQOC636iA7CyS+Fr4EXwbmoqFEryZRI6r1oZ//AeiC6Xu/24GpojXq
JZFJtZHvhM3rLFMxDv5vxsDfVYd8HCIYqmXPn+c0dsamulvOpVhJy4sH17R5/+vv
TuBQU8E0NxBIjoBVJpax52WdTU6baQblrOtLgwwbIrO3LNndq6fMtHzt4gyzeDin
tgFZwQhODTQbkM5K3v7BlMqc7gc0/n0wuqQj+BZvTW6jqa6T9kweb+E4AW1GeGwL
4pPdj4B9bDnyIa1cFqyOp6A56pvMtH/LStKFS5tyL6YH+2gl2avFjC38B/KciEgm
+gUM/R1mDVtr0QZwnrORF3W/dv0E1QzDm4ptMqrlqo82fPvQYC171arnh3jm2T7B
hAozzT88sPFtoHeNv90D3GPquDLsuHMegOZDJqEDNpmkktVPMVbyrdKHExb9g5An
Totqo5cj8/hNNQsHGnqZzAyD01jiaNwXbMwyrBFLc9bE6q/s6tnWwHxCjNUiK8AV
cv80OM0gJhdlzVbSU78ZlC4CIdyrJUHWevUWt0LIJ3Kohmp28o4AfhULpWMH4UuA
DLd1OTyYJPYXeW5i9E/FnZCg0++A9bYKmO/NW2NetUk85qu5zu1MxAqDoapEM0UF
LBGi0xvRo5X39zreikrPTj9WguVsViDyOvi2FKlrk2tYb//UFNUloJ+Fchbou3tb
vtq1mwiMCnebxATXMGYvfIbAXr0ivt2fVNqybKpijyuvpLS1xFsqVUuWCpxcNns+
3YU3ICR2uYFAzM0YTRdq6/fISJXRmVSc1e+7dg/YgATZTRsBgmBgcbPp/IKtMxXA
DwiTUxD/wJ3kZkgGi5ned5bpWWyvNdHb40Yr1lpQxzLhDFhi4xM4jvQ12+TW8hhu
ffNNiiDb8Lp3Hw8xG2FVrnPr69Hy5NwP8DknCYPsbuf1nv66IJ2R1343QYbKohUi
1vuzn4EggNNY18HBUZ/6orwtbmCi1DgbomhKLJ3PdZk+Tntl/7y18lsNBdywnnI5
U6JvF7MAlzRmyXijIt/nVeO2vFYiwsoE7DXdCHqhDKudlsh8/NJvE13H7AbdyXaE
QnrP6FhAJNKXhbLBGbRLUBAg5SdHKueIJUTASdPm2fKmExTPoreOJs4WUKbk6V3B
xCnuiRtOw/GS+jg2VdsjscMW4sL4aH7X2KH7e88+hOuvdztC7EoJQzqIdRMetilY
vRQTJ8g2Rnznc8kpwajfehE7s1HpTvtxBXgv2/Ntz2MCgxIgVsTZmXZnLQ1o2a7s
qUIIw34U7CutWy7pP5zGCALeLo8SK+DLzOnUqh2qrE8wK0gdLc63/3uSTjvl9sPx
uVTOjgZX9SAS6ELmNZOjGsveOJUnHRA6hv0bkMkCljW6AUr9E53vwHjeLYRxAIeA
PahswUneCqvbtodHFgMgauz8ARhaiqryREy/SH8YNE+7uelUAByvqo/L+uaH4sYg
oiYPqeCR3MNXTfHUQ+Qu9BRjN0w+LdNUU5sjfER9Fp5Ze6cuJ+wH0OvxfYlDlq1v
Y0OXxoZtefpqqey6cCeP7ksvUt6IlrUlgPr4Npg89vm6YioePc5+k4e9jTCS0rA/
0eD5UgI2dxF4wovj4oktToC6QSxisHC1MpYgjDHII7+SlnMJnKHvN/ZbFoz9dpHR
a+DdOH48905yT1Wu2cC4RisAR2d2Ev9yFp805i3HEdy8dkDTXaY92FbQbKlitvcN
d8gxsKG24/VUZb0xSsoNiG77tXT0h/yI+44vUGW9K0taKcxnPqDW5zgI8LGarLvM
yLSzGJG/C6BTYTpLw/P7OvcGwbb+Yfn+iz1HPR/ccvss7nqCSVyV0RtjHrjnSiZU
N28q2ID9/Lvt0R5l6ZAsfy9RWoE4ShaeQ40pKcu73ys74pUNXY9BiVJKzRw/Ya5C
n8FVL7O9cI1G+bi64hduvqZLuBiUgh0LgZPIu6gEkXk727hkUGREBoeF2nzeL+ZD
4f4uLfRZIF89TsdZJAy/fzd3gx/oMowZBqZyt7W2+whkA0LM+xRDBUohVO6KFqKY
9Us2DMnVVJNMjOQ/VARAdCFEXLSSVykMI3xsCER43Q9q44Iym7f/7zAxc6djnOad
F6v8r5vs8kj6ANhY/cBYTbdOJYcOvSneunJLeMlcvLw539DUqh/FVThqNJvz0Lrt
UnmAm6lu88CE0kVfWQ4ehyft3CIaRI3QBvuit2Nq2B2U9C6ISf0M3ixsBzo2z7jc
2Y89mLF2ah3cRUfVIoDXwnphotytA+ONFN/3lZTRZvsp1HDlxEcfJwP+aNBiqVxn
bA5NnfEOBc4HWCk0JbcETR8MLdAczKJiLqhyMXCkL8j1pdbHSwNNb5ZdZZkA50w3
PTwSK6G4r8v2AXa+AjetUBlRvsKOow6BVwiyWh/NhrQuDyrOLQ6d26zOIyMhhJ+H
WA49HaJuMh1E5WYA5uYqDoMQxqqE1oaNvKnQPvlgmnZBe0XnD4ingBojS/LR4UGP
ewq5pcfC8AlJmdF9VWe1QJ+Q/o04NMrdbOQhUJT6Dgm6knPaEfUS2te3ikMjlUDR
xbdapZW3fFYitJNBcsx+LtktL/2TAkKs/2IW1B0IDi29Gj2PYtJFPyT0Ib+gTCbX
+Xu6IUKq+4J3ddk95KWIVxjp3DvsNRX4OrRyMGr3mnpfJ8DsLfIYHEIvCysfu3u1
oREIN8GRAvBWxDFMcwnqIzcsN5CJzDtz0kK5fmAXq0W85Mam1qDRJ0qICnDvbYCK
DPYNLnnRdsh1hofqSVR+o6Nj7fCcKRLPrDHM+D8Jrb8xpVZs+UKe4jgOQR3BNMH6
CScsK2kH8PC1FRNpbTiXi7FgDkul+NDEQ90iwc2MDCm1aHuYRRwL6LUFN9OOebU5
JZZDRkqgPjP2pNxLnedvRpohsm8Ws4qeSXK4uJ24W3PjMS3qK4a8JcTZ0aVnsPZC
D6qnCZiLp1CwjbcTRb5IXTUp5se4tYXeodGdXztbSS2bQJGGFL7Ly4Oqo46xDzt0
S1tGtHQbC8OKuJNE1pZ24LjKZU1wS+ZvyDCnuLwwZF7X/hkr49/jmNoZHU5PlCMs
N4E1JpBLqmLferaey2rEFMxfOoUWtUQTjDbM6tTC4YCe1CnY72HE8F1rWqdrGDy7
LHGHW2nBoL2mYWfl8qSREtbAsCIftlJhkQL/A6DlClENMl4ZR98JnLb4WYoMTtfh
ZwfkOo0Krkg4LbJw6PWDry1R9dWGBAcSpzebpudyhclWihKVvGsTEBSTXLxNLVqT
L1nTYE19ydnspqzAf7v1NRlA76BXJxnPUwV4r1P9nTxvRBaf0VC2e259vVSxMA3B
TxPPVXVcoSTXcLJHTetq/NYLeUhT0PAGuUEGYjvSxYJssvMt3+HGnx+kvx2oa/SJ
aT3uUqILTa99DCspU1MU/95+S+h0suM7E76rGvpy37jKIQF352Q5f3X7bc7HgP7N
8Z3Cd9hE6WZsdp263DDhLGFTNoHQtR5bE34saZzmSZzWBBOaeVH6FEeGkUjJyxes
IxGEO/UjIa43warY6gilsDQde0ytrzYxDfZTHI7Mc0anEVYqWFe/i7kkXjBDq0Jd
3D6jD/kD1VHrLdn+BnGYnPYkvVlZJAA4t2gbcUClDxKjWCXuGX0JIKQVAtpsYN+X
DG9Bq67jPUrhJCrGQ8jgk8ZSOaA/TuQHki5MaYeObzLhlahN5jqwvVhkjJwFcckg
h876lG1TJM5H1BQK84YwJX5iorLvMr5ze6GkAmtqiw9Ybn+4UgUogYoNLl5uLw7J
MZ4pW25AVeHC4YkaLFsm+YYF4gxU0GuLu0R0t0Rd8g8VKLMTwuZUih1FxbdSV258
/QEtZgdLoNjScYqePagGtwWZgev/82WOMCSf74Kju7XJNedV+ooYo6IBRMc5w+dd
PyycXKF+0SGcYjHWRAAgGET1JU/t3gC8uIaLEA17vKDR0zeUK1LQk/9t0/G5ASGp
CaanQVH62uLqwX+Ij2SbnwIpyFs9htpg116K5Vbw/JQcUUtrOXQqjNV5Ols8fJt2
mcwIn6885xmRwCrS7vNkEFmfJCbsgOCC8IUsNVU67B22ZGJrI4adbWc+IJ2yRmXx
3uCRKCQDtmhXDBZDyxyXuFXz8ySNoPodmLQHStShS/C7U+WzSWn1PAAAXy4ErWJe
edjk76k94ncBtCUS2N4ufK+zYxIx0f3pXlrIqlOw+jbyFCGSTnRJVrXcNDL/ptgf
4rdtIk+am2mwB5CQQ7/3i9sfzPNvCaY9W+/sz7/lvqHpMPNZb4zc8OK4fU9aVyoF
JnkffMT4r93NoBYbwbsLNr0f4OYyHjmSvOMiZVEiSok0+MC5c06Y+WyOyEvJiMHR
hZkLg3Ahs08J23QrkSXN3dLNqojLT1dmL8a48/eJpypEAx6hwZ6zgiR89O+YxcPZ
62Bpn5Ur2M2qzIW8+B99wPClHilayeETkSkxcyd+AqTEhjON6MmOAiRoMDpKICpz
l2GP3w4E+sD5LGdBUD+5lIUkdQ7sP0P1JrB4lmsQ8LmV9M+6DkxWjoc013qy596k
oT9ozmtfyKzOksyM7Tugb5ij4aEiM3yWQPdOhplzPyKMt0uzYs1Hq+GFNup25cjU
v93mAYG13KicSfJMC9NLp1vm7r+pCNvwFo16wiGpAUmE7JGBKy/V+YtNDPrDCQJ6
wB3rSn2EFt+8iwWa6n4iy0uCCMezLPn+kn03LqVDErrQvlnS4xB/cKFxY3y8o7pF
IVb3rDlnZfWLC3jGP9enSsKSB9A4n34jjQqAxs/+XviLDkmVZVI9zY0+BOtPgPnT
26gr98hSV1uxcPp/wyNvFiM7t0MtDEJuPGXeuPT2mQ9+PxaeUEDuMXf1xrukYwWy
HY921/jgXEOMPSsavyIPRCzC3i83P6exnhQctN9QjTx7vWny2B7CLQoSadmAEla7
SGJy6Zq684Lp+dEqpa3vyAhCCBNqZl8M1nGmo1t4EYpvqIHzx9GTAYFyVvuetopl
12xFTce1vPIcM9tS9TLMdIR75dpPJgGvDHHkiWk9KhTExgQlq6niAHd+mdDmWeAG
3yecOG9E7dkwOMMDIx025cdTO4gxWggZPagQlTLXGOlfEwIxNuH3WKHONpQd2nMJ
fH9bHtYfykpB/bGkewwLjyr1axOSio8UXx4X/oqneduOFyv/Z02+hQA3gq8q6wQL
MMmjQ5DrhpivLQAli7eF4vilewl7lS/5cItH32ImlPwCFoD9QF+UfHspRGKmGTr3
+uJtGBt1JvgKzrIGRvr3xF+l9L4+c4PcnBFubnbmreak5x24VcP6PZJbln75q05r
zo00jhVA6pMv/aNnOnJ8tjfEuKVL1+qMMJTYjlt88CwMUhUQKo0n2HjxWnZD17Ng
izfr2cRC8sdCa1RRVAGhMF7Ra/9RRRwKhMicm9l6/DlFGMJwdzNBdb4muEQBl4PA
rr9dT62SikYIPvQUw+Iln86aG+1UZZ1wfn2dP/sxnbCZISmWpyHymL4hLfuszgkP
1Cm58qygIF4hzHheSSsn7uhHwYw0m1c7kEZE0g9bGsPEwlD9XZ+DUBvyGO8dL1J1
xPtSE6a3SF69+DqdFVb0wR2//Xi1m7GzVp4LNvFPIfMD9frirlo1vxpgDocrVGEM
09du1GiCvpb3SI5ACgOmzN+9m5S3WI4vLWRGcvzO0kziAKHV9byzrifMg6tlem4O
ytY+AfuhwkkIpjQkQvtNUVVHdFUIhrdQHthbtBQs7dN41f8NWYX0nNfgvL99p7ev
koeMo1kljd447IDzW0CyI3M0AhexE4ouEaTktxMUpsEzW28SJHDG3rOcjpmX7aBq
HFl9Qt6jY3zNw+ZU03dw5o0DaFl8w4b09gd7Za0egeLPfIsQm9r7K7M4uU2soElx
XaVcWOTBdXuhjyFgDGy1rDGljQvUKSGFKS6jVg7+3TjPvFiEOadRG2POE/Np/HI0
rFQgrRiUBiCRkSfSAMiNag==
`pragma protect end_protected
