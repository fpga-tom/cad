// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NPBykOy0rrBexH7vTh4V6ukowMT55fc8yYU8N8bYiHsmHPV6kXYc1bR8NygZ/GU4
bpXTb3KDQkAbB941laqVseiU3QYeTDOn0y6CZam8ng3wC3wPrABFuKn+ofuFexSq
1C8cjFSO9qcQ29jVgfFutJg1zBDdtBFnVCVBts+UjjY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22000)
q9gB7W8gckiSZlAVoc/NnnUqOODSAM4nfbVx0VQResQsxhiPQHga3yOkcw6wLt+V
SjJILx5JWvDKGXoafis3DMGhiuQZet/onWG5i685pXGN8f4uQlwdqywJqb1YWA6L
HF/nEhFJBi4nKfvWzdnPws7lS4GetAZBm3oquOtUm5quWRmFTY+0WOsuJOadfHVR
PcRT13YPVHRbqDhpfO0jxeN1dzF/hvz4IufRx9UH0lcITC/6IDUJk1P8YAnlSBCz
pyG1x7h0pbOqoUne3OyP7CpShj8Ej/TlAf98Y4Iva5RzIh5Ao6BNvE7K1f2qlx2N
0+s4AjJxIiP0OgD6VbpERhex/OhFOiaheJ57oDly0T5TGB6pZSrXOUFShv0Zmx0+
I4Zj3QUcIEIdendANfrnZDgIisCW7mwedrptt2bfxoFIDq77+5KYdyod5PObV3Sw
se+/jdYlmRwbZEs27pPoHBQVafRbSpaF2GUkV+bndwQ1MZxudt5Wlw3kva//ngyg
mc5fh2wi6K/d1P0Y4YU0dZjCxH/c4P/UPHrJsMzwO6yOSsnHyj5cQPAvPQZnF+ak
k17ZExIEOULkSnmGUIjFm9B9my1DYPC9dtdS+WCEsKUWR/eEtGVZjL98Tl3afRme
eVyl+OrutVaXDagMeY9KcUcAzgquyTYRqS0toWqhmWDPIIjgYDiWmwaru0mC7D5H
Gb0nJvhmewgDnsndoR8dSi64xKoL1YdNy7pm5YHEFDgaSs4InBJ7T5OspoEiU/mZ
gPOq7kWs1Zd02L49cao1Qwyn/Dxh39DqgyUuhig91M1t0Jo+bAs2hqDwnvoXXCTt
MbiwcnZjcKmljQWHowTXGWRq15Yb91DBfbLnICiYziwES3MIIbTMITOS6J4roiL3
2wiBFmMFsp1vSWORtemrG+d2wFIC9ReNzs+8TuOin4H3TLovsHcBskjJjr4zA+9l
bJ8RZNaJuUZW0t0un6MR6ReRDqHaPyaD6iOQl5PqQ0B6oXv/MWdVV7w/8OUPi499
zRSZqXGlsoO/Q+cWHZQ2Fsia6UiLvcCU5oSc5wLfCFsrjficQ0cCc4+QzATlJDQL
ZbuMCu9x3x6S2jlGVxeygUyJDNYlGqRGdS539uMyBoSGZs/RKeEPBfFhHP2I8D1T
GHjsmxoUxlXvjgBD5F0SMFcMq5iEtBI1LOuWJ9Q9KlcfjtPtFULuN4fiTyp4Jqi7
nsFJTeafm6d4eEvOAPfDexFYKYbZypQcV3CkXNWGoYafCByLYwhxCTT1upyZj6uM
fO88sbUIHgk0rGexiaJ1cBSFJg9xO+jwH1wBxLC9Jew8IzRwsKRn5wZSMGnhGnXQ
/OkQi9nQlID1o1PVJ29UzFbx1XkaYHDib2HAF036IBZcChig1DpuOpXII3o0c3Sa
jNsfI1NlfQjD5gBON1eL7P7jfVkUpbe8O8m6SefZuTtlRXzzgaweAkANnVtCEsDR
Wep32TMp2szMjrqcmyjpjUaFnbwKtge87Dq51nZwQAhH6HDMCBLoRMmto0UmLNYZ
RVuaB80oFL/BEby2tR+4wfiARBA5LRE/YK4DTc4pey02e4dkNzOINyQA7ThjfiKU
gtT8QxY0pbhN+kesZdG7Skr7MxaYlxNwX3e0tGpxOZabAJmkMUhWksnAhYmoy1JC
Lb+9jCJTWQyxaX4IUkDaDfRE03wmsjxOo+WuRz6tvu8U0i3bnMfYuunFmcYr8Rb6
m3HcW4Le2sq2FXAIKvlAv9cNriWaG304T4k47ni89iD+PI76ehtSAIk1xJbcIdtq
KkFOazAtopQbxUv+OL8j5uBJ4nebuo62JyqqfiiqvEPMDK5tA444h2PWZ1bq1K+T
aNPQoQ25gIJaIscxXZ9kiYl4zkfRVp0a2QQC6L+Ur0IkAsQclsZ2q4HPkZwyn+SV
KMTLv8zMkI59ELeFBWTwRrsRW9Mj0VtUeOLahqmAIhCiyd0RAbiyObccEYfkWqo0
IB4aqo1GhNHh2vLpr34MmnXUjJ24Lvx9RB7aYn9sH8NEmD8lTNLLFZKtL7CCGfza
QyPdXw0PUTxECEGR8+Chjl7Dbd+Kx3S38ULxKs8zkXTG/92G+IpNlOPopLMPqvKF
2PzvGEKtxBpYSs6V8X43P8ax6IVGwxRMBErw+eDI56PdPwrnz6Rdx1SUTe38ih9O
9vPH1uput/acfeBDypA+liKa/ZPB6SC6B7PHy6tCaS3XN5+pblc36MApaU2WYeHf
/6hz1miVhoN8viufKGzAUQe/7HIqSfV+9TKNOOTt1KVaaGzIOpUPYsHFCWDsU77v
hC2KoIAHkxRHrfrurDiLHXKoc/Z/ic8dYLxTIaXBdrTpfL/MpEoVwhM3uVYqumZb
w1RouDJHaHGwB+kSB8ebt3hu+muabaPfzD9saKlfSzmtFRbtvxBzgdnuwhOdh31x
8xKw3gZNwIHhvekJYqos1/mtb829AGkno5mX1uEgt8EYCkeRQGrxZUEfF2+7fA2a
3LQYH1dtn0xEmj9dgfxmw0N64EWIi/0YqZMkSf3NJe0oGPYB1PrbJEuskyVz6z4q
RVzBVO8BE6tsaXj3gzVEKYfZ3DHvTyIbXWwWfjuO/uj2GacNak2JpTgSyMhKt4Ll
F83njgnSPryBxeUqcIFdozOyXT7ad92zfIc0M6hOufVviU9+Etp8v15YHDjugd9Z
wwwHNupleFecpXu8EmGmdsOa5H6sFfTgCjghF9hqHpkZsB0LaQc0FuJOLhDB4ieM
f2kncs+DuZJ3FQWXZ/HaxjNCBW0CK2VuiWOn8SCV2E5uwVGiWd7+UT8x6Awee2Sk
LE7syS2U4Kh6V1FKuNn6FBZwIgOBiJ/e9hHvL6utxH2SWB91R6JemLqBN5d6BZG7
VcKSs0I2c5kUf1TD41QJ0FHkbo3He91+Q+ZOf8ZhZloSO8QVz4fkYsb/4qE9AlXA
38S92q7E4fVmA2ZAFPKm/zdqYE6TLqLh4fB5JUNA0Q0ldSHfb86e/UhEOkyicq2A
Wqz+AJGbdbOikkqVRnox+GyiyQnX9blMSQB/dZBu+CkKx/T60+S5lCNoW5L4ufD0
qHtN8V/qZfKAMzuPiFIdyRy6BwQFo4nipclrws+bz7YCn5Ef2Lp+4MMjtA22Itn1
jea/9iSG67H5r2G5+77/XUnIwiTFNE3qbjnMSjTA+GRUuL/BLlWaK4oi0c9HbW3d
scY3n8qmidEQCSuuKhhF7/JlHSGGJETIg+grvTa3QzcyGX7A3V4cu6M+pLO1Ve4O
BuyelorpaTB8v8xpDe/lsnMvJktMNsbUgx2ELgwfncZ5l3MPIO5Mc1g4TJKDaOvm
SFHd4F2lUxxXDhA4mQCKAYeDLV7eh1mhMVNvnTwANjzpqoyhyKuzQXqR004vIIbS
09BptrWCIKuGw908nHEdQFNPFc7J0q5gVNWlwTTWR/+5GijnJYrYZs4hNNWmL5TF
ObYyUzQ1GjTZma4KMhLwRVYmW/1XVZ6nim4axAsLK11zi2qNBxywOKpagjbV9kxE
VHKIoCqVmYVGAMSZxs8MROM5IO34Br1g6/TlUlx9CClnl1CmTi5c2pzgqpZ5MBAP
BICMVVjVtQEQPLZcBaX2WkyHsbVCrhEq+ROHVzOZlt8IhoIR9wReEFVfsYGdy1Tu
QvvXxFsOxGacVJA2mEht63WPbH/Vi7HI5x6MrsNeqh1M7oZzwwahPlr1AoIc6KI7
9bvHmLaWTW0XBXLE5BRHPIWbTEioqVN36hz5O3RcWIm/rD1t90TNjOBAVNHypAfq
Gw3w+DpiV/zwHsDusKUOBarCZ1wJjwR01VLJBPNXyuRE+MzIwTtGiNEQ2QaM6pqR
HTTKQIcnoOO5fL3IE4hBdetKRrqfoqfWVPLJ0nPs/UfJTo6XfBx/MW/CSBlCEU8n
bOAfx0RNc301NuG873BMgOd/ppOv4dx0dP+xCA8Azn6FcVNimcVcsfEs/VQKc8P8
Aa1TFcwvkf9jU+il1RlYBwX0Lxk92a86nJsM0VUT1b0E92NXBK1/f612f4MPabpq
fKTUkvwsgAXQV55CbxT7L69WyKt47cVcnxqKqsCQ4J7NJM7bn+tzZOAmtW7Iga3n
ZOX5r4lFYL+725MEXD+Vcr5YUSEBY1we69p4NM2bh0pBQYne3n4lDQ50MMpvf4Dj
Mw+fAxDuHMmx4vmeeYwUHuRz6OktU9EWke3F36gdrbXUOhtPNynVrD/pDJ/TlMfE
nA2bQE3QDOQsfCCm2kLf0p9+ABt14hyHqo0YrfMaWtSgat8/vmKhUDGmDfIOjVY/
l/kNXzHEbB88ek3DRCAYO0dhdK+maIbgo7W8jnc7CxXaE+S8Yh9BCr3U6UPN34MZ
GPr/rW8Vd0Jw8LpMJkTln5w8iUGvrvfk0Cg4HB6kL1EKZdPQoPJ63BYqVKyAmv7l
GC7ShpIH2BCDrObV01uPuU42jkrYKNyjGUlAM7AuQT46sxV0UCdLXF7aDBBqHL9T
+9g70o6TtyLtqbEe01RPzYzPFso8cAV+nVzHjdEJ4VMKnUWNmq3GGaGHRgnCm2w8
P90K2GD1fdTObK4jAP9LlxXOhSrmcnsbXDhMBlpM7fFsc/em1xlErqccozCnddHI
JUnE3Z56JY6Q9qeCNhFpDYFe8wmJmunS8nF0lhD7wnDqWxYi5Hs3Qlbm80/wEI5p
2P51VLTmAW/OIFG0/Jv3vBoUZMR2vITBQWM0Y9evWYtPdXsq7q17TATmnmfK4qEx
fg9GpzXdDGAzKT3Unqg/YbvMGEmW+5XrwHX866GMozfPFz7gUg3Yf8IhcrrycXbe
6OkrNQ4wPE62ogAQdoOI5A67mUh8qb90wD4/TYWqtKqHZYMw2WQ0VMZEviX37S6b
2S0yM6vT3GkscTmJvINEMLUuenfmjPa9bwp2r5VgZt4bPhnzjk/HWrgnRJqOzqlL
KJ35CWIyU6Me5k4ZdlhbNlmahven7UjtKFio+Jh0pa9I3SpiZxoeYnZRNTgvlNMg
Tusjn7CmGw6eTlz8P018HayYiL4Rzc4V+e4zIGMfrNDa6wzOLzJJ9Cz8Km8Q0x42
9hgJcFxBUdcE9BlXfj3O4D58vr1j2/To/4o5ghgeUgWjwZl4UyOI0+p6De0rJ6uG
/UQSSBBvO7AavV+YlNv/3PXjkNIYNqJyX4NwW8qbLAk2KvpZQ1iA2uM0GvAZqSkG
s8gumCRUdFOP0ae067YIrhkj2yQhXGAfR5MCa8H6f78HijUBesMALvcmyU68mbSe
swlY3BLY8gl5tvFIIx7BFjLKDb6v+qzGdH0kBb4HaON/4QqyIE57EH+QofrQGsQs
ktZknD8j1pjWvt4zBU25KO5lmSYrqDOANK2m21tkW0pzPHGX8VZIzJr9wMn/AViD
i/q9rLz5d7BZrzA5elN1h+A1Bqa3V5gw414/n++Kcts4lTJgA7OkSmNsZtvEfTeh
ttHFLSp/6P3NHemnK8lumpQyJWQP6fjx4afFRMp4m7pdD1SX9q/qs30ouTMuHyGf
qirqls7TPqsmaMsYFf3ju8BJtPgKQ4BFxSJQ/WnSqRT0QCtohdAWRf+PAvAK7fO8
gf2FdxtEoU4HO6e7JuBRA5ya6tmKAdp5IWgAVgtzc1A47LlQCZ/LEDqJhT5siyKk
OlxgMf+QRzdEzFCADUXc545yRU7XSM6FbmddjJBqjbGuY6kipCN1ML4rrD5aLNA5
BIiZCMqGzA26d593EAms0XE1h3xFJOWQvK7n8uH1UZpmekS2xBI09qDeQmeyqbwL
+YE16IWFO0nVzeKVDb2epqBjTLB4we8InGf/gvw6wJk/T72CIQ4KLCZl3xzOkit9
+Nd0N/jgXOHJDGou5HQOBL4RBWcXNCbyM3uZhpeQp2Vu6m0rT6hmzoGux0elaYIs
UmFjB7CUnmWw5TYGqfT0twYHIdMd5XI7EnwEVOkOJaAB6A83mfkhAW9H0A+jxCQp
prkpfXv7FV0DUGnXjJSR/FQhRDHXTx57UTwz9pJ9vhXbEatYqvoc+hG8PWyrb6ip
LU6h5oAN9Oss5FJX9mSo/uCdmlBtCB29M6MOLOPZFRMbeCN5KoncxwVgbRZ0qDF/
H87dfuZoa6J7VThXxzJW67Cax7NegqXdonnAENmVFFXmQRhNYIdm0bL41m+xiKjy
BTQBXZWCb+juGgNyYGLbVDSjcJPzFhYKWfqc9wl6Ow7NxRUNZIEdkD+PB/vLvcjL
YL7QncIfxycXEkuFQixVlsPwu6IuBhsWypSWsgnuLQgbNqu1qlG/KUR3zsdV6fkK
edBPMQ05sCeTtnru90ruTexgJnpf4eoyNotAxOJCWgtPfmgni2ATgeayt6eqc3oG
rLd1bPT2TwJehzbgoo3IfHcfzZKp8fKDa7J1m0O7C/ToD+Cexfsislbjc+ds+fJM
JnPmoD3aVFZD1rYxIhANDc74SVwbvjPfJI1v5vIDtYpalSHVYNJbKb0mp15x1xwd
IdExfXcKmM9c9PJWNU0mpJjRza0vVr8IBSavGmHWcHeVBzSBV3V+99/Sk5aErr/s
r7yj3RFVyAtYT0rFwhoqt6j19lVTbDKLzyuaJbPn7R1PhZhiRgUqFaJ3E6oQbtHW
p5x7K1L3wVtFbGSP2rtbGQoWfCJ7btJpVtvnBwFuoi91Lxp3Wf4qZhXDxRTI9ym3
jf8I+OlvAC0Xlx1/TlCxPm94VwfePf+oXn5uhaYA06KLpLrPUMvl37DUAOSb8GrI
tvm3BX4EL001+r8dat4OrIvhy39LtbFirbQij5JcaDCLYhtUoPpTyPzmfrpXnWKq
0ucP5W8ISKziVX6tO+hw4n5xDgyxugPKzH71NXJYaC6qxTZjrxdEeQKOHcJLU4wU
r8mEZYxm/ZhWUmOdttzN2pGTlAUM4FEPDtZ45FQiPAVWNG3WecezqyJHM/9lZk/h
5HiscL4ZBIwvf18PG0ZbOp4D9NhDA+BvR2+Lage2i+oPm2BHDWfotTvBhmiabJpr
v6YKXaqs0VuxzWI9K6o8sSqVHHEi+87l/lhlCOKtQJR0asDP0+LTJdoG5nslRIeX
hpmMjSIIcizM9BKvy8at2aaTLRWvY6iM28lwfBCbGkqIGTHLuL1gNi9vh/C5zW/K
NhCcXih18twuvqy4u2Lo0UW4btUU1PvaL07aG95f64Em2UkTKRJJrsBqiAJBN8eu
0YXxl34LJ3eXA4jr8kjHudH0/4j1MghWqTLQX5R7yvtsGvWG+ZF2ZGF8gkD39swj
duTEwBwm7wjDBJhtIsp0Hxwu2b6q3pA68hHImmbYrwKtROvVxQMwHwxuwbteobLx
BO3iC8T6Eh3vZMZevKPvNnh7bf5O7UzF73fhuDo+nBRNX+3LjupIhtGoGS7N07jO
cX3UKawZuSptE4PzAqKrR9xgGTVPzuWa5CCckIr3HM1vQsECTB2/q9f5o/yQWllo
N/RbgIfuBEVoRVpbgaVHVMawdTqBtqjDMtSR8MUy2oTkr/FkQEu8TiNY/rJpxCJP
I/mkUPmiB2K4iHJhuNZjFop6Qbyhdsxz92yLWhLYHLk5HSX/B7J0bEG+fhbaXIxd
ihZLP6V7cbtqiZMxWbKjfdxH5VK3kCJpvdBryFRCRWcjl3ZVH+hso5W29vMYbz6u
k2DWKGqK22ZgynxiKyziJD27le2fKqie8hqQA3HOV+L8A/sky64KrIxyXkLBi473
ZAO0tzRkj3dwslpWa82aDOi2yOXj+yqI6rZNVwQkLbw9EmVjI0nl9YdjwH3MZVRE
1UJRxDjEynC6CDisnN6PQsDKNRrvIVlCXE7FUE0xOMRuyRtSDlFFIsJId0aEv9fN
el+wBxQbeP9Fss8+cwE5c/1D44X94G0yOXFP8VQOt2KXRk4CboYLeO3c1snxRAvT
JhYba+bKF+55YfcFFke6y4EBBpOCRdyUWtUgoWOl5jO59i4vPYEVUmpTlMaPlPik
aM6bGAep/zcesxN3kCK6bE5P1kzsdswoC2+Iq96owCu3eOANPi7s1quqbRELABR/
5f4PA2sHi3UR7plVjhVWt9SiOM9XksMIiNt7tZIbFA0PLIelpBnDa4hR9ldwjplt
oLSjWCaSzm9fT2wckJ2zrMjE2WDwLWPfLxicCOSBJPIqJMlPEb6DYFGL8vqUD8UZ
7z2ACdjISkJywvrxFZGhYN6tJa6D6JE/8IHjon9K3yNkBWLZR4d+rE/Q5QgoGntJ
oMjuFufVCl/VfI184XxEo4XVJym7ogp0FtbB74NPG7Y4mjMp1Z9trIvJ9AvGvFAX
bVIpNbN98G2i3LVM6+azFR1gpQ73jwXQeGb4SOYnY6x1nlpt+2baD9LfM3O9Z5F9
LZ85Gn+6h50Wk/by6+uAp07mZZ5RZ43WMz8TCcKDRl1M4EMqvhHbP00griAvvlUL
3qSUpppMlP2MVaV87uoLDWE1toBaKstbrw4rwMauiEP+Ezc6ewX/xoPN4/7ZPBAS
zjpljYuloEzsDAJWrhY3rjtj2pfKwp6cn9uZUcqxKBEBNjQvR0879W+X/QakVobt
nJ9IjmF2H5tlkeipbzJmLFEbxlcC89xw+OpAMk00M6qlsDN8Hvs2AVmwV1I7+sNu
E8mmNiRdrDOJmj4wskHihqT1az4qu5bxkhqNwEEF8AzN5gsOMuLlFZm7fqLS4+To
4hx1jy/xnBL3pkd3YmJfbOqN1P7gzWOOleDYn+F8mN97l/Syp9fbHRHPmsYPvKsn
bA9hMsvTggmTSVIFlJZuK8GK+fKz01TQUaszjiTAoi7MabNZQ45L6fAftXRoHAg0
QSrGtXjfWMiSgsDyQG8thK8RbTGE/Hc5Nk8n94v81hTwqxpYusziDvu6uJoPCi+y
w1ydYy/1l5A1zFx9m7unNNj83O74fm63LWmDh6EJheoVea7kJarKRqjlpDwq6wxt
O9UcAVjxms9UyVRETsuz38B3iU4HAe4zbA1KQDClZNJ6t/FgrNYPiHws7lPiQZPO
YEnE6YdhXPF99I4K4bceGmGAyKsrptt1UnMApTq6cehW0ITTUr0Ov5I3pCjTKVrx
xjBkiKQO65HhDPrNykBxkuTmJvsBE70Zw7ljCjC20XPj1xJQD072/0eYajNjXIXm
VNBGiJNl2g94afkDEGRa8bdlkgoDIwmp9yXL7bZTcKtzsIcaTtj3Cxz5kLfQpG6l
WRgbsN/cjpB16pklupg63WdlzwW9Z57LYhSYWkISFn3atDiWdzvSNX9mV5ZQ/deI
nFsH0llxBR4urKQ1r1XzmRmSk8yMF8zuQBwgKeHMB9jrjcOjTNUgA8IyulsxErhD
T+MLuUq5dThupL7+z91GoKsCzSpJlPbs+pflEsjrtTE98B/9twp/pd1uUCtJhbV+
/PomCsFkk21GvJ9wdW9f07Kx5lcPxa9Jmhim4yxJSXhT1+Z0SIZ7Sibqti+Dgwhu
5fZZDV0n4mLNM1etKWrj8H/jF+JZuxv2CbFGV2KEp4KxghCB3B8HOaYjps763/9A
CLoXQGTp0fFfHI56T4bRfLWimlT3ZabXDRmavIy/lIwmxIpF4L40mbbVXprKePxh
qFydkb7B0i725BBF5yfI/qqJ/7Umd7E+v+cN/Iw8cztVrxLF0ncJFTen1uRs3SbA
AiDGojxrkm/nL5UhaiO6H61Jv+AshA4Do+HTuvD7PZmCMq/BXa2x7c9CzxayyhCr
UK3P9ZxBZFYl100IPKWMy78EQ8+R9WCdVNtgwM+Cz8+8kO1ABqahNQiiEwb5ePRf
A9vwNEwH7JIG0eUTjk2zDeQbzvXP46TcQvLcTJboUENBYuw5aRKnGjMMW1zgdjPT
pBLeWnb25kmrHZ0vKBMFhlasI1qZwGp5CCZFPgU3jfjICHTrT48/oSKJhpOzhWge
oevjWJEdUV/RfHtJ1ffCfCo0fx/DyFAOSKT3Y1KNPeW9LKh3O4WXX64QDle9etUE
B4UHRs4OB9HWsftXM08cUV6vkDKkbiZcr4y8T3PWrnY6tmWUMn5/8lO58v13o38e
POkJuK+32v9lVtXZMfBFXOJ2We5U5b6Ed7xX2DmeIcijsN9vk3HaI96jz04iaDeW
cwL/L+f4nONZKg2ddg1+zu6ePArYySlH3ajHKjciKsuW+POo//0/8UFxD7RQRJ07
msFVuM3wPBowjgTwWmAfVZhHM22XYzw6oMTGi6EJ5Ieokv3QWAaN7qSDKyTFBE1K
/JGK2odJRP7qGE88ekx+N6dMQ/ERQHPzYGklx/FxX1s6ZjDWaxQIF7N6Gd2IZBtJ
Mxs+kvW97j50c0XyaFk8TVBPHuYy3YySV+DOBi8O7EgoYABzXwoKtW/5X47NyITx
ikpWgYvpaHeNuLBloF2C9UhjFW9KrhVQkYj4frCaKRQ0U5yxgtBfCwfO2QEoVTAo
6UHh7YF85oX+Kzsjk5Wz6NiAAKNRdAxtAI2ZHR51uNzVPooUfdDy19xscoYjC0cL
e/nOzk993eWDjmO4CZ9IJ+z3kkT5t35E4sbSLzK8kwGceURlVpamRHtTvUOkH0Ay
w/RyebqGXgZiPQbFuX3Fy4Hsk3E0WeGX3y/sf/ToRbF1JAIXhxuH/zExEVeXgwL7
8gg6UyQGviGhqk0d7tItcBhjglokApFsTtAPcViz+6Jg9BeFKqAIcDOMHmZS99XX
lFmP3z5u2Sjtd2eaI8tEq+WUnDIDK/7Y2L0pd4z8Fqw5521wCoHUpYcDFqWOuliH
8XXYmKmXdajDyOXUpuRyWbzkPz21+Qvowpe6cYKcnE39Ldvvw+lz2/xOccDEgkEO
nkPvvBDOOJNi7GxtBcVlfTVcP02RkoY0x4bfP/H/3xLVuDZcGzBLKqczM7TR7QKY
zJVuapgammN54JCRqDSco7VxufTHzpEIUTMBHt9n6Iuv2LQha4RL2pLgN6mUHXfJ
sVM/Ru2RX5xEc7SjqVTHTHWPSSUgUMhU8PF43Ei2qrEP1oRCVaGKSNNy2XQggDmK
iL5c6Ehw6YW+4BW2gZmGL9aJdCO3kweQq/8CL2Ts+GjrkLruXiSk0n8KfTcLBPf3
IVrwsTP8m/QHbMq0sNE01v1kknpeIzqKUvBENDIWE+NU0OEdw2wsKwTB+shjsYWf
0bDWgGhaZP+GDHhK+ceUZbhzQrqbxJmOTHMF5zB1wXjBqDiGG0wK2pgoXxpGnSFL
q+ggPFm1MDdf561Z0qQOSYj4W6KqtSt4A8QpRrLctoXcAZhZlqPTYywBUwO2Xr7V
ungOXxaIkCnahzS6KVrT/h5zU4bIgfFxFhurO6r1QxK+t6ooNBjrqlQZ9vt9kVah
1/+zV0HImVedexZkGNsTgIixXbkfP3pE8vXBhZWWRP7ctmnh3lMzdb8icXd7jRlV
Hu3OvdIrgwL1EvmDbaIaDg0+cryZ8M76/z9HOiE634Qtz/CkF+CpcI0P9DHE4UQE
ForbfDySWBdHE6MaERaQzMiI9netQl8yRAISQGfiyK8lOiyHBZC1+KKI4nKNC+7s
4o36PuyoMfzYCIiHMrzjVHC5KVrYAbRwmocUi8LI1y1A1HpFbWc5IpWDA4kTFxGt
bKaKv0Ig7HNZ5wV3IkUdePE8oT1jLdWwq8GEi/V4SvqItTAaXjfMNdAa4832EvjZ
WDKMXYJfE1v4mqE3l6Bx16tKObxbkC7ujxz7XKB1qFKGs1UbupGdjYySmxbGIBdr
71gLJR+z2xgHIE27B5lRD+wX061knZeVDWBkTgQiAMm4xnb5bav0wAq0Km2FHdKt
iuqPkGSlx98duTi7J/l1B7XNZQICgkzdHe5cTDQb0VN92yURy88mn4g+n2VSewai
zexpqjtjQP2PwwprJn4m10n6zRQc+3CXKpWyS9J7ghZPfsL8hXlJ+AY36JmfvkYY
wVZ04U05RcoEAWuWnI39KtzwxvXSLagIEvlxpDjsbsJ7tI0C2dtdN+HXRrxcZyWu
M+Lvv6yCTv5rAK96ZPwbjMh6b8pZL5d164xd5QU67tITN6AUAHt0tgKy7+pbwOWS
TqgzsWka6eHvr9kCX8oVmyE60qpoV64639zOkmWDtgJgvbG+VY2O1BHzbwOMkbnW
FMyeVoHWk+uwkVCBHprt9hoBL89xwnTaf24BEASg7c9a5fd3uIcVQnNIEQ6O/rwX
/f2kJMw8qzwYMH3DKKYR+mQkW+mWUqbUro+S7svvUShVB8aRTQOvigTfU8pz1Exi
oDj245fGKwhjuMupDXfNxogrvrNrPTEDSILf7lnlF69Tdma0eiCUbqSwIv6efxlc
bV85kQlUvvxq3R1aWQrxkR8wE90ggem/cWMqmb9CuCy4sHgXcFfd9rEMUV0DEToo
JV53w3W3M09xVg//9RbM0Wp6qzNrWMJV6HTwcrQrzUrvCdsmfTdpgr29NeOootzx
6VquEzZSNSIQell1PaVR1i1TsJcQZs3HoDQEgT3tVuVfcKI16rsjESer6+lKLEUZ
4GKf8HrCB83dW0oRAhcT4nSI7b5JD0ZFXYSEJsEA6SNiH8934OtRLIWaXeLf0Mdl
Ua+aqoO7OX2pItVSwlzFS+Orb/iiCQQKMBqCTM3GgIL/wBWR5u28CfuFHvNclHuD
Ity3GtlEoR2n7JzS4cBb+pfSL3dtJCuJwUu48F2Znoxzw9CyuWcs7AUFT1dc5qaK
1vx7N6HIh1UBRIqB6oKKDEq4Soq7e5Fa0y5TzVbSEkUvTfiuSHGmwANAD4XuAivD
saAayZW+jcL1Xd0iww5EsOdCNy3/76XK3C3WSL7DW6RysacSTyx0u8dsawDAiH/w
cq2xfWdjixAvGusSmarF82BnK2f3PjTDWF0LoS7aoLjVUkFJE2PpZ3Zvf1UE1/U8
OZPdfewiMYbKHN8+PYgjqFuGd37ME9ibarh3hgdRtPjEVl4fTEhokfPBtQe6m/2+
kpzIhAl+LL5Drbj9dJnaR5K8WMARH4A5EYEBl4RkjjYdVPwcyBlTHlJk6N0war85
QM5u15csUeLujwPf0icbJTbGJZuE7AkAIBg29vQyM5CjnMCG0Zbp/JOHGgz6/Y1t
9xYvTVAZrZsOib462FcFG4rI2u3f/LcSCWjKtrsZ0FHf5nHqc/pTylCwNQIw/Eec
RkJ/N8/04FzuFiVOrgCSwZWnCL+U+hqeeIT8kzyDx1MyVahDqHdDXCnE+1gXY7Iz
DCCNzzeZXFUrTTV38DDw4AliXEILWvJR3cNYy1As4wgK+o+Y3tAZRpHOsONoiFkw
C2eqObwgjZn/LcqH+6JbGIltnBN3SP9KQvEvbO8GhFzFbcDY1m+BSaz6Sr8NIZbq
RCIJx3wNXAS4A0UeYz/lJ0i+Iqj8VpAYYbXuiGP0dSi8KKeaE9RgbvGTyJfwziq3
Rcw9lHxdRrHp6YAkOx9/w2X3nja/rxGm48FzjiULVWo97x8+Maflu3M//hLZJidS
dX1R/z07Wnht1WJxi/VfecQpI2upMbGbFO5AWGo74C0faqmNupL47+YNqCcFX+5z
e+Om04wq2KBLN8b7scJX/+Wuk6gLIurP+K7GYmGR7p43L9vZGS3KgpCudjsDucAo
nY2WDasYl2ZfZ8GiMzjldrOiTy7VCQNEDpdRxxBQaxzR5HH9QsEq7p3pCtdmc6wg
t9wVOdVUFVj3Alrqj/RWgzO2Aj773g6BDMGl6yv8LI6XhgcKrIYAwwUeYDrtLZcw
T+bmLWJvm0yqNkjemfPqjkjlA7t+jfpGWds03oNc2RXQq3LEzMdg96F9uwK7wKvO
7fWHjYFpKjz+svRznykPZIrPjij2mnOtgJFQqgMpbnTh/DJ0WjwpqJ+KePmnELXO
F8TVlXKsj11ButmcAI2h+iG3SueY8tiZ8zpZwEv6cHMgQ/8iUwMWdhH1PlTBAIjq
La7IVCkUhqJW3KYieMAAgXt9r0l/dDkzdYKhXGmpukUnzU+eWI0c74PqF5R7RUZ5
4me4bjYj7Ay9LOi6hnXJw9IyoFc9eR/DvCc0TAFuUdjjyjShVE9CZOTpK1rM9oLn
xWWKZ03CrKWa+4y+JA8Pz9QtAyDXZqssI58JdpX1af/ajEerlnqWDAlzJJZqt1C+
VEDl4th4cZd8BYDFcasWVbp8npAUa7Jj+P3F3+lWiqlVXHQwQUvrKVW9tOa1PLbb
3U/E20WFEBjSL70DV9qCfBS7kqEgPt812QmDPja+EHxzGYL+b49fYThny/46xJ19
zz2fd353RinisN8UVjfs3UKZdV4ZXYp7+H1aoKGTIe4FHhoEi3lbEvFxhNmsGKuJ
GhRymTxQzZP6H3GPesNJWSmZzJuy3ekrY69WlpIgzrkw4f05z6QOMGsRMQ+FF5rj
Cruu2dzQhnFriAtuUGwmVhjSbItBksdVwliha0sf/+E5hI9QKSxA0jva/QBuMbyT
qWOxycv2zam8Q+RcUtDiTsV8WYoE4qf6zZXZso511+hyeCbUfgQGks6mgzShkFZ5
WK+xTv0bz7Yd3X65tdhfRLgnswYQjK1GGClwMJpRTTga95xtQMASfWESZ9baoYHL
qQXL+W2WrGl2Nm847dqwGM7QOzkIeFAAEYlab54E3gqN61WAHNHLCb2O0Z3ez0M8
KzTIaabQa9SrBG5C+PrT2MPDdfsqRhOGwJBpl/n2ANObnGGBMBNO/NyU+RQjGhx/
TChsUZ2e/dQUB7wF/ZwJblFyMSub6ZHuv1k39pfpzc6lBloGOJ9Vvy/MnbS4xLdO
xiKJyvIrwAIvVDlfhRu9H2itd1bjI1RGB2xVVCpJC3QLy8Dnz8pb7oGVZi1y4o27
mnkGsd75vtNp2gUfNze3Bt+XoxasqAODhckyErNe9SO5J0l+uh0mBo0QqA0F0VFR
epOGXnzQ8gZPP3VZ9QQCBUQu+/YEaBZEK6Ie8fxLVq23yy/wvIlz+M3rXqYWc7HT
jh0PbiBB9SZyqcFCQ6QgArXeIpALoNG5lBmSnc7Ws39AM1hQB7lU1JEd73bPFqxI
HjwyOmh8jDjkP+SxXu/nfFPGtexcb1+psBeqPLf0EVaq23kc7AX0oiBgslB1p1g7
IU0RcTjtqskTiEJZImCdm6LvqnMONyAnD44BWg/Rrt2fErsOF5XySN4qpYpPxKJj
KaD/SOxi9GV9iqVLqoU9X9hQKe92AkmKpxAv+VZpYb1qZpZWCHvtVXuD3WNdYPFU
9RInJo2ash6fm8y5YftnS7GTHDrVZsu4sNTY4aa4nptzTgDX/qEEeNhv0qJ5jr3L
wTwkH1Cy7HTzi6etfbO4cv5pspFaLEo/1yy90NoH/MUYPHRipAmUq9CxLmFD0RJp
NWdPi3fdMM3KJXwFKdqpO0O58Cum16DMj/b3nCdxEA2VK21DCF0bGW2xwwWDWrR2
G8h3NlGR9lhOPCNBrvLEVu0noexpqPYZ2+SLQcGGlYjbdY5o4pllKOI23qcbg7pS
9Ig9qIcE3wG6exxp02FmL/Sk4Da/GQypfQ1n2/TwnwT5Dmqr9Q6OaGAtSnlV4BKq
BO+l8r9d2IKo+qfqqDGAGClW/bJLapRjp2r9ioCaAqf0patlBTX0bmQ8PX2FGPrv
lcaIVjylZhkDkxzGbZ5EvEPB9W2Usl10TVL6T6MgbPSxLPZ8iCw4bqgajmtp/G0E
a/WSmmpEqlGX6kxifThWh6x9PyPgI83eqNSSImUq8opte4t9cDPzg0Al41HNvi66
61VLMT9XnM89snq7rTqyO5iDoOcG4CXCW4ugyNOFesBZydXDSUyY9iM22CHFeEEU
Enx16kw/Ijj3Oit1weLRIdxIquN9vYXOsAvOlAGmRh4Gughbh4DJ98V2cpOB9Ytj
wnYREeHhaHD9K7OlwQzXq96U2FFZ185J1rHSlC/ACxMuTDQR/v8iY+ur+ydCnuW9
Hpobun6ao0zmVconIWHP+OjBSuXQ88pA2uXsMBMrQ7eBB+O0taot9/bF6HP/EsVK
rZob4fzidFiFuPoEyM/IvG2g1sL963118nTWiRdUCo0DtpKHGzQrKj3lYXIp/5Y6
4VQr5/yHNUSPGgJsc/DmEdc44QMTnLrvEtcv4dVXYh7CJtAXfQNhbTVxZRLmtdCQ
WoQcf8agnnLngU2Khxp4Lz0tu7bA7DsdTyIv04sr9npEQ3Pm3xH+Gf9gKvAZHDwQ
+nkyar32DB6BAaIZROtsZAQvWWZDdeHWOgLJlczwe7JGw6uUNHzHT2ZLLcyIggZl
WL9vhsagx/B0dWGIPr3+k7aGZtp4iR02bqReQWaGQj9EUD4sXZS3EOt+/q9PiU1e
DxRVykK7VeuHMmknDa4UqE9wSg0zdizOb6j/mAYsPlyLcESYmy7OXYtovDjl15M9
N9osODu4l1io7bFe3Kqab9KYaDRXnOcMfoLqrgku42WbX7tVEz8WGOoIumtacLdN
SYz13qX32SZ0E9fk1jHu9nYc2CchLmX6boszK9EK1dIWwEdmBtCw/EE9CzJ5eiuM
b8XlSoWFHOq5Dnc/gGnlSPvYEvRHAyvz0UQbHxg8hLeZA3rlFT6eSG2kK0f1sySy
F9iZj4zfrvKyFmgEkAQdK0V4vUZ9XYVwVGXbDcZ0Pw1W+sPwHdJRf2hhI/gfHyMi
ICm7aMhtvS81IVsUgvzj5NEhq3ZPM3xYtPoCVACINrvCbC/omswxYsevnBGkDM4c
hoLuWTyUjSPcYXckdnuYwKFFkGt2Uo3ws4fO+JoyVDCoRhkHw2Vuyo2cxWXhDp8c
UbKv9ajjFCfflP8hpnXVX1Zd2I9OJ2YkON7/9T5joJwTaxFUlxRYUMWQfcbef7jK
Az+Wkk1/q15CcoEFlYHLyT4lQbzsMkA0DwfcjdVNZyJ4Z644/Qk01pN16AsSkpZo
GRpEn595hcq8XjeeCm76EjjXQKZqC/B3a9Kv8sha03XVM5n5NvvPYhjFGwA3hjxW
T+N7b0aRta57iqN+v63hiMbn+fC0ahis0yTHWz/R1BT9MGaeF7J3dfMdb4PWotNA
lVTggFTJgga9FDum+nQZf7U6+8Ls9Py3YMknMgCiAAaEp5SlShM436VQwe71TWaI
LMB9n44jBVHZVbV4bUXxIr6BhtxGjzZAkIwIhaGf3rp9daUcMz1h4GM3YqC5Qvr+
IDkSIt9V0997lFcIFQt8SwYsztlnzFO+hvPry1XJdiwGtLmkqg+YgsUuZQWB3+0y
xKBJ/zT4OUCWi4g0htldzxFuwgha21WRXYcgDMnUZlvDlQ5HyK2EmMuFeX8HUwX7
x7BoxHLuQYA/LNRms/c7+WdZvOOZRXdfgujv1FDjp26WcXdsvyzGc7ueeWdOKG9e
53zc+BswAs3ner1MjciXM/nj6DM3vleKE/qsUXL3Rv9X5VHANM+vJUjDLOpec0Cw
IEOgpyiuWrOM0ZEjFJ+zg5La4hAVy1NpuwxU1udXpcEErqVZcxWQd04aOMPlksdR
Cm/WNNzqmcCcEHT4GuzygbEZcwspLHqh+9Li79JmrzG18sW7MWoeSXlVaLxh2JHY
wABcaNHDpGHD2Tb+E5dDmOMBGQkujiBwOxS/NtejY/qySrCRi2tmvIOhF+2cwTJ7
ni9t/HUZUN3ZliP7j/ZyFHxfeq37VBYVRxvktYJUdI9QlkwtssNqCYxfWUBVU/Jd
/8Mk8dni+F/oBMBDJkqaip2grH0CTmuM5sOtHFBTYWTXuDaIxd3kzts4LoO7HysH
uN+nAzqsv2uuSjRbOBOj9TA+CVLt5Z+jfRb9rcXTlb3cDGssND4YKSqOG6xuKrry
O/cPli6bvbtUNQU1b/8opWGFjR1P47cT61j5Mx6WAyZcjTGj1fZpsaIBwjPZzHUZ
0m6Kmu9WtVdp95bByx02CDE1UwlLNT83FQYoCDOJGriOWVq+hxL8pRBztHzQqvoG
Ighfxv5Azv9PgyEusgB5BRztgWt+fdlZADuG/7uX+/Uih0StuveJvF6TA/MhsoYg
MpetrpOW98LkNwv7BCFK75e4+FPUSn9zU0s4p8RA9SImVsPUYuVgK8acb1P5AZtv
uQQlDQvHLo5VwqPRJyTyojNjIu1nJBm8/x1+h3xd7zXeOf//BQZTOCfoYAmtxumg
Sx3C/ZNX8DL8VBbuz63qY5Vjpk+p61YX+N+G/3fWcibK1ADAGEnL1Xqb3BeOp+hO
go7zLVZYsgqX2MO7ZutNN+UE3I7MocC0K12aqat8ebZvlH2D3f1Iz3wAZrZn1RH2
r3PwtpJxLcfPJd607xNDEvqNzyI2LTaa8Yotmr+FyUSv+WHv7XXxpO4nj7xRLFJS
ifY1x89O9MVMefmKPst2O3Sm3JRprP+NjSew0udkNHuq61T6OsguSQTBldTZP7aM
5KWdm9kLdh1+2Ju3S+/tDmzYZ4BRCw6pB6tE3x8Ng1iFpv5FVfaM0fryFQd5rLVL
klXoYTIPPiwC15jh0/uxBJ7VDEDNY5jYq3+Dl2QWo4X2nJV5JnJX4fZhAumaCckD
uAF5qVA2Ech28uPd9cCgGdnMZpeqF2OqiAiYquu+1AqLzogr+X/Xaz/SlI5gPDiD
hZmcOMLDF+pAdCDcBaSF2diMkyEz0NGPQ3naoUgu6nqKXqw8J7TdLqhhrQWbJLDD
zDaLKYIG+T1+79kGkTH1YO8S8I3SzQHYM4fZmA9e9OoaUK2Le+TSnyuliWLOMm2j
O1+VRtyIm9YXkGY87I8cvDL4uYP/ZeSqDBJnWtBIMQ6gcl+SEHzObrJXUzMgcJ71
/VA/WuMm1EdeKOQ551JhHd29t/oet4WqgMvQdDCQdekoVmhgF2V8bAMkWzXJJjgi
AUDK+Cvk/uw0HB3DXwHlNSFSo165ass0w6ebuUXS8WPrbIcaG6/v2jTwV+/iRAVF
XOA1n0Jfj69hdvZFvvVidoTo0ete2Use9AP+YCrYL6jWbndhSc91tSX9e1/gsNa3
ZJH5cFd8oqTFOOT+484gysI04hWTSV+Fnlts1gJcj1gpsY5CKN39cHqfZqt2LKRX
NvzV+f3QHII86IaTyYjq7/Mlpn1B2h3fCgz71LWvVCGjQ6ePK5sVtZOvN58R525K
6XSzMb82rTaDgi5/KoPKNNJpIgdACPfFP14Ci1bSSCXXMyE9uXnUBhgyxnyt/88C
vYyzzY89dsaSKP1/6KpNvcXQ1kE5ekK0hhKegZ4cEeeZL+MWKVQgSAIOFRB9kBhy
2zSwTeyRzdv3wONdFKFANEZUUUS1/WCoMSqYYsLvggoCnj2tuYVfgKqEV8uARZoD
gptmcNyhreqROkkJGAa+6y8whEwrkd71pQ3l9g6HLv4U+CCnJ66ZJJ0rAIYhZEk8
bmFtQ99I9wefi0+WcDN/USS+fjQ/gq0EtOGOP9OovaYkkEkYcGibqWCcIPUsSrTD
yic5zAp2fBOk6E3deOA/YSilAKJsskgxTt1TtFh9bq8chI9EkBIdN+UUe4crIl7L
xNFM3/OE8zA0bwbjNLa9tCGQXPi02jROxG+vtLJUSblXR4XnCwv56KCm5uDfHSMp
HFajk2yz8IL2FWWYdCCKQMXBhUtqXWqPBnXDVqBBgXyCRvkknQQf8GSueEksdKNX
AZlRD8hJrggVVmRD2cMIa46Nbiy77dy0YpgA+CDxCEXL3Uph/2Tc1tB2BBrZNZFa
FL0seS5/04R3J2MgqG2zk3xRc740TWiX2+/TDV/5Cz2Ik+narHamsGrRocvrnoBE
ThkoCthB91AfpKkQTcPLJcelRhJVuZ4zaVhZVYfYaUlkjLy47ZqS9qu/ZPgIzgsB
8mDV80R9kgp4HVgwwLyy2l49jiIBwur1DbU5ZY/ymfjdiZIkXlWEvU/plJaIhUZi
1N8/coQExPTbNDrX1M5Ztc2SYp1WnDXsSyOa1B3DlRfJ+l6AjUwD518fPFrYdHlv
1apAW/QXvJndKD6UjyxL0LJTU5laCTNaTy5XVgGdRTE1yjOJmun76IzB2vIgN9kc
0Cl+/Vdg1Dc4g+RfL7WQTdfvTkBqFSS/1GSzhuZJFqgjNmSPVI6NvP0DCGU/uxut
rNAYA2aA+QVA9O7KDT7RMhiFHk86ZHU6p0xxsqmkmzsbyyQGygRw1zMf2geqcFkM
w8v1GbCNx5AtE7zAzliMbcqk9m84RfqihGQeMPtUSW89UnZqQ+qabZvaNKNJrvl0
+lzsOlQ2LOzBYYMDfZHfm2QkYV3kVwfuPZmSlipJ0+mY86yiz06gIzSsLj/Z72dM
hFcyDLADNaCGnvQ5bynBlYt3euzf7ndmDRMm/I5rcWCkIChYt1AaxwzhiDhm2USa
hRVuaR+1MRIPS3jmHloKd68iK1j7fH62ViyeTjVt48WsSy/lAKecgg5WF/sqa0Ju
ZVNE2g/Pa9ANXDrJlutG7Dx+4iGZ+1b2oePoWEgXwj/JIaMz5d2mmIb/xsBbtlvg
Na/djNLKgteCLafeAIdgJJBZRv9+/EUjNGBDvALFxakPM4ElLe7UJpyTjNkq1RBb
sF4BmmQpkrh/vTuioqbUt35UcqAu6u6R2TEs2aMLsgZajccEDAx48tI3gjW8nn8z
/q9SfshrroRBSsnggRDJw4qOOPbovKp3DJrQ7wK+dxniJy8CPVXpJv+DWJ8Utqwz
sB2btiXF88WjhHyDH8tM9HVS0DwjvHksy+hvQ4NxHQsvcbVmaOsjUPXwlM9nJZRa
wotJgbh3MQE+vNDrCWnbxixY4D/Ko9plqVpoq9rUhLkP6f0ZZpm2YMg31DKK/9rt
KTn2J/LIHBXfNZtZtyLkMwWMKQPGH90WCbakshUPlF9GykVko7X8M6YY7kNNFspw
uWGWLcUEtR0GAOUhOAbI1aZQiee39lM8pCz81GxUeBLBCYNqN0Rwfr4YQ17dVjir
TbvLCTRVtr0eMD3H+PdpMsRJy9rL3G+CBh4ge3JkHl4G4H+y5y8CWmLUd/n1+fV0
tlU0T3cfbtgzhd6Mmum7cz3W8IX6xt7G56NAniPDHE1RJgXJHkjrYbgrixBvcguS
wrC0kmk/nZI8p4AE9f79g9e5994rlTJ/OSGhGpRx2hXER3AlTPzGreeUy8O28RB/
wg/7ZA+7MQd2OmpMtsNCK7N1D2PRxTFYu2GgHOiZSbNjh5KVF8MBKnVS2Enmo/TE
q9zqKwLhPKFH/5ZrvYRsYxVsgl7iIUA1gFc56qrU02t4+8x0JN9ouk7WH1HTBwcL
SbXwibTlyjT4cq9Sd7OgyMlxKEZBMmjmzwRhy3EKtI+O5TeSqGbo6MRDwx/fNjDf
RAFuKss+bYB8ybcUeYfrTfxYViNmA2xy9na5KotPgSzS/6m2pDLxPTKYK8S27BPi
K6rLvovfmuXhUj9KVxX4uGdM6gziAHtGm5cX7m6lth/rp37vnAyMrWAaUnNpXAJU
h8NlNBrtO/t8E9AfCo75LKg1TlkjmWv0nVQ8mCJgbxTeXe3ut+Xv4HXXldjVfB3L
NzGv1Ac32Oymr2b8t9M5P5e+MZv1l+VhVOwj15nSVqeYKZhlJXB12HKcChSUh2ox
XtwnFInS2vGF+MOZJkECX9MbM/S9CyfDkbO0rKOO3jGPKMpcL8jMUz8k1MOGgR9E
yzmk9KfNlmc3Sc4shLQ7+qs+odMYwt0f6iRenAKNCZ8JvERf1D5b9VeWuLb816Aq
vQKITgazNTQArJtJ+vk3aCDZqlynqbQT7hZiHyycw2mxqS6tlq5ZNGCk4Lp7ct4z
F0BcoHMuPvKBlEdZmgG4RkopXajUyXV40m/mYGeUYuV8p6o7gqAcLKICYC/rywfc
Ov8/jeo+4XonzW4GIdTID4RBgQ0zMWcXaH3/vJbAtqRCmLovPQQTC137RBkaS5tA
GdMnkJBG2ZLYZtJ/ROHSmDYozSaW+Ed9ow+Oxu9spgz+I3DUXSfpSD3LXlMh7hdr
yPPScT/uXjl5eBgUzugxxUGHyJX9DO60bTQyRaylJl/eTq6V+unV/Dfo12x1ghf1
ip5/d9LLuijxqFWSFf8aZVhRZGgDvQXF2DGtVCQvUXNtK2nh9p1IlOhzaEwFxgyG
X+rfA2CKX7xI+lOsjW3Rveq4h2fG2qHGGEf50NDWmatoXbaPGLnVW36vMSkZuI8v
HF8BTt5dagQkN5VD8kQx3eBJlVqD4QZFi0ErhXn/H5jfu9jZV6xPINN3shQY+Gdg
3EMOQFCatQ/HBIC34+/THAXSgF2P0iVUiZ3cALvzyWBnetDVs0MvuKpK8CwYtomH
r7+r0Y/dO3ljuHupgSmys38xpuyEGeMAdKWaWHLEi+L97r8g47B1D9Cn8VZtkAAd
WeFTdGkSnJ4atp1UcMATwqC2Zpe+HQPY6xHk7zN3PWCK6ZlkCjBi1nBiLjecXvAv
cV1Rf+hq2TmjgQWSuZ7yxpZwxQ7bfvHvCo1ZTmHW9u/PxxTIn6CqqkFJADFOWCin
8OfUIJ/+qDNF3Hija8T2mfj1iFffcCU4ib2ck6FKowR0KGnXhOVpfV+RpvVKzw/G
iL6KD7GCLDPHwYWEYPJXZTHyNyjYeOHDkw868R1NTiEh7KxKtm684IRoD5sYFGQz
7oqGDJz4j3o/2IhW48sYfmOmZjBj2Pu8e78odHKi8GFhGIQmmnTmk7zUEsJ6m3pv
P4Nvrv1F7la+EQidox67FgHwHuOGJe7llokzzPrrKiglwVhVvNfpi72wSJWzsKWb
8c02mTvOwQkhEAl6MsaCeOF+QPUp50Am9SPdKzxMBm+7Z52F4nGKJSgnoabT3LLl
wZQnX1P2G3T6QwREd/IikFgQhYgerY7cmSoQTilsioeSJ2tXYFq60gAM87dbVCSI
obWw12KjLivsMjRUAkcSkqCPcW46B2jRy+6LrZSvQ/LOVaHUXbaJxb/C4ZaLI2R4
q75xP4f/Mm2hWZMceotFwmtSjqs9fOS+tfx0PsXWD8IDemMESED4VHxrw74B98m1
2nMbfIxO+guIt/nfJDqffjhmIGM8AjogF+4PMR4oX/RUEkVmJ1WCdlH5dmtDdwZF
cPHmktAvonv/k7VM86ZmVu4kmJnb1WwDTPKCbyOJHaieyr41aO3mRtcPyjCGUYtr
IAptBw+SozIrpPwKXamq3qcVrZH9ZTzihOhksc81BZrfDRNz8n2M4HIqoDkZ0HC7
B+ZiBdDYzJ+ITWzQboGBXAmiHdm1zsGYFxLoHP9bU1TjFANdIMVdc0KbozR/69ib
dNuiyqXIyMvIKailNIU1pkeKzvDr+v6hayErLG/3BacrZUlAannwUpuQ1sr4cfZ3
CJmLmVjPkbBt2lJfRFM65u+psoccEugDRe2NEytHrlrBQgKsZc43SulOCDe47C+x
GISo8Gkadd1CWH9u3Pfz77v//R/JPlMbTC+juztq4QbeWGXSHbzlQWtFIzP8xm6j
pk87lq4kTAimjV0qUnRntLnjYCunnH/EUi2gNqPil30PKhgalSPfWnkBXTP609X+
8+eVN9op0HT77TeJlL8PhpJ+LLO5T86W3kHELEPwGMqjfZXI7ubHYhdb69uB3gCv
TX7pXuhdbymuZBOteazOXFdHAL+WzPMnMQC5kqlvoAQmrkxNCRS6RZI/87jh8TYr
uEKzC5QWdafV6t2rBBIo+d6f5s6xVQak+X1W3vGldLI7uKWAqY/C47jT19FVuuDb
EU/vJOvoeqrKINTYLAqW98ObqbO8GotPQYKlVNPgmGc+ZM6zO1z1j2O8OsUN+6tv
j0ZH3OpFXKZ8O14hwcqvX4u4vWKWd5Li9V8iFUUiSveWFTAf+IA3yUOtmvxxdB1y
iF2ZZYSyjSsaulPVs0sRw9NqOV1jvWKBBGMIQLu/mE8dEtYqL/GzPr9DKBeot+JK
PRDedzQuEuJbV8Si921bbFvSfoA4ztt747wJLFchUvmfgoz1BGM+c7/dO+MxJsD7
YsAWx9wXGKY5J3WG0+m2Lnx/qGz/yiCHr6po7ZDmvZundSGakKdsW6/BHea3wI3t
9DFOs3Y57m84tovsn5vPekfhNNh0mtMI9DEiFp4JNmnHPDo3rf+GDI9cmVxV/AB5
snEO/xAm+TK7Bt38j/Us8pF4GRNCK6DUuOzlA0LtmaK0toQI9sbjExWODYhAggcs
dnfjJRPcEtOW/cg2wgA7xq5AytdGZ5AKOYkkyUf+fA2zd8CnfmQYtY/tfQW9+CzP
+TuRSXEhVDz9TsWyGIm4oUvw7lqaLSnRh+ZYKhiQVkJwaZSBClGIVX5Mzh8tc6FA
qD+LjPoMwvPBGbZccpkRuwczfE3GiFqyC3BHZpfwv+f84icxiyxfs/oi+cobwy2J
hOVJrLur4NKudi82LBI8wT/E/pfrnCoCsrSUptyMiY/iGUD8qvuBEyDHDLUBLPbb
UY+tA/v1iFVpZhMIxW9hR4hUTJ414wQx/oMZTwh1CZe+gfuD+nGdc5KBaTyWZDpL
z3dD2Oo/PMM89ItlH42oRNwUji1ojTL3kDlFA5ThyiXefdyBYlcBh8VyldbUSI8r
6KiMzQSH9sBLcfVvs6StUgixfFFC9tH6MMHRKZQYAnCGyp/venZIK6pxF8T2njm2
oK0D4mq8j1MgFY835nt2SnRvNXbP5LohjYi8okjmEMtlogH68INNDUlut95Dx/4r
yIOwgDIUkpm/gbDf3oBIKsvYXFYlZ5hQeBI/2buxxR53PWsFNx+wHlwJR1PMcWcp
IJ210LUMUNqVRTvYwpw/2RKDcNHkmXJ7TkC40ya8ev5v2cAPheR9N1GW714fRXtT
0x5D+l/QgbuY1gVthLalFjsk8poeAuiNm2tKGQxx0Myp4LCrbgv7vYKu86LhG/da
kcC4N/T3CupnGskSLDs6nDI5o54nz5/d9TK3tpFVFb5U8WDrzWJygDiOGn/tQEFV
ghAkEGAtFgsgnBbZEPk8U2+3BVMxYHnaesd87yjEp8/4jp5+5MNaCCXHYxLUtJz2
u98F7FHmSy+rtz9fnPNOQh7wbET/pvPFWxHwRvHmbel3CEp4PKBZs/m1ibT97ulh
0IvWabR5tyb2IxF4Ow2wK6q2PbfrFAMFQkDv197iYzxKRUU12MID127s/BqQPVyK
yVh0ZY8RTKHf34acF3nUcMvkIFpxEEancPUL+C4BN5UF1JGMM5lsbh1Qp3Yp3MpR
Qn2Yxm1X0HknqxB+Y4Br8wpboSTjiWbJWZ3qVHDtPXuTpmwr9gJpadyWQ1kMzQ0+
TNQ4Rl/SzMJmCbfkfAHdjZiyR/TzQoJBfbg7U3aTGk/yKLCRzGM2hgDG0suDznF6
ZNnMpQ4Gsjap3lSyu5VCSAzGli/WHv9eT1CmC1b6l3za+TnCN2tS/hxE3mHkB6+O
KNRiKH2/ZWUYk7Kb+WybtWDZzcowDP3u0LZXQennrYWZiqpEMfa6oQf2n9w/7930
J6lAhFMZwx6QEjtC88RbZXWXqdEy/tBKa7kaIyWIk7/X5pppwaCl+mUw3xupyNc6
2FXnHDp8a3k7IwhExXCLIJ4PjLz9a1lPCzrHeP0FVMr2UXVZVt5D9SR9Xzw7HXte
8SN7c/pO6ehCbGdUCG+wLIx8K3A7ZXHP3v8v2ANf8lFYzgDCmYuFTk/+GdrzqhbK
tWyHNiWzE5quV6yQvnoiz3KvosrbSg2OYo9cI4yaLtIj7pwAYqWK0CNYksR9xYCF
dCfEJUSowngaPxy6pw9Ru1lckBDbhmGNnlM0P3+01XHue6srGsIeb5datfN8pSQi
dT4zJVQQu1Jt6vd3/VwzUZXfL4LaK6EM9tNE0z0OtfWnenCeKdESCmtXLS8wmbDl
uoUsacTwv1Y1bFuSJE+iP2UDwjgzPBzzfOH9vsv4ZWmlo3VFr/nXZ9LXeqEmq1up
XU44POFjk+oJBfzUhBkgzTl4O0LTEpyeEDvXTifNZD6+uw/uW0Y14zPbnFM1XPdb
X0V86+eP/uostvSWTqCiDYilv6kWp9BxmC+PzbAosVfZMUcNxN7fEadBVcqFfYiV
SSgdEQpVJ291xVNo7BlcYhDZKIZvzd8gErzs1z3RWPrvjWR4K9JBYdXdkMk+CI4U
rDCqy3WliOD/iYbYCfh8uQ+g4n9YVs4yhnhtQx9mq898oh+euLiBvL08l4cT6NXJ
NaktoXycIV7dDRUP9FJulGMPOtbUGsuFPbPA4W60zLW/IMuceCpnMvzbqh24oqcB
j9arLz/jhYeSsqxWGKXgMmnxqCk6XNCzs/+8JFq1CGbXSS3R+5muw8XQgKu5l9wZ
fv8mh2njABmFQ4juRzBKW1o4bQ6D7cVVBfjA3ZCLTbcXfkFXrwcr4b77Edl9YTsT
V1DO/FsCY3kM7Qac0gI5SNlBxn5husMd0RmNnCWdGjht/no0veGx3otPdCHB7wwe
q2SqZ89DCstPmDtUSRz9iK24UAEx1+9rxp/rAXIrxLH24BGs2fsEdz1Opdfxpge0
Xk0VfD1TLr7mmh4+r3iOhSE6bM953R8WvZx0Zcx6pBRLRDY0qBjcDPMhZqZSTU+x
zK+43qS76FMx94RRp1qzZDfZs2HLVpqvwh2eVTTEXFFOwbOomvK4lbyp86Y4kkMq
g5gMFbL95ODr04hmrXrjk4BhNStj2xKS9ztvwTHZ16N5nuYF/uFnGcOuLoOClzc0
dqWsWu44ZIXU4aBB2wfxJu0PcK8k2D7jm9NmUQxB0vWFkhpTeH1KHq9puQ0Nrm9Q
zFWEiW7bcSteqvIqXYmzbRcoxf2daj6h/8ZhNtkMGW4vTvcns0m2QdYI0z7wGOwg
DUBSqvYwZsu9JL2JhZnOg6fRrTO79PB1rhecgk2ZtR2OcS6tQDbx8CDrvFdtOXgg
zzw7WHsR5Pb/9oNIUhJhjfnEyBOVPA9urdGwRhQlWiYGOms19WMG1IXwiAPhtlXi
44HlDknvtCf9F0uhQ4rIu5jouztMaWKLjrOQFn+oMb2NRewOy4GTHSWuZzDaYjor
NKfI2OZS85ZUt1RjYArVHxFQhnF6SelslM3bdRN4PXjImKEcBTVCcdAgZUxfvy5F
KNsHCxfw9vq9FFbeSk/rFkvfr4ECbGLi8CN3YnNlwB0iLPJ3EGC3Ms/05xNMnatx
qSK9geu0aRsOkHXDVlOhAt8g0qb4jSfF3HaVovAlUU1PNmq3/RNH5q3s2bmX/5rD
dljT/tuOmbK/EHsNv8Hy2WOZ2s8WPkMT5vFsw3lCeUukBxWxyjKr8E+U1sUcYnRV
1b9wRK7lt1Gz8EKlBc/RABhCx6QH8XiKv2lz3soBQKE6hpfYWnXUbTFOHUNrZczE
+vURSEw5AIAr2tZ7jKf9BKrMWqHZ+Z5fqUgYbtfHZFyKujHVracZxosc7YERBC6u
EzUGIYcr29mGX6x1EMG8VxsqzivK1TN8niwZcJNd+G02jnjbbC8wBU44k/XGdQ23
5P++XKK2PGJQW8mXdPIwf559mnL51bLfrLIydtXPFsaCS5RIK5aPYxQZAsEkiiEC
dfxJA+72pFVWyMoVZIClkL6hegTSBAWnS4oIQBNV1eo6Od67eMvNOzMp9rAvOzAk
vtCzxgulCDdBNJ8txypT+VI+Z4XlN/Ll4SY/8qScnfGBNK1ttFBLlb0k/+efNy2W
OPhOeZtYO5rIXMWdxmHYOA3fFTsAuTxwJuxA9xYdOtYd5OX4GTiQf3wONbQz9YSO
95dtI4233gV3EU7tY7LOsbaimz8q2M3dWvsrAF0EZA7IebXhapmyD7WhTvJlOD78
w1MCVUmCEmULl12DEU3A3rV9ISR3gQvM4NRhdiGloZkKJlRF6nIBBumXEu3rxoEG
rngCt/Wp9k8z6AcEvIvFxqnF0uKrnYDHUnEbvnE92PbIGSnvWoPd8NdRZF44XEJz
x2diPte/srew9xM03a5b79TXWlmkI0h+Wplp7kcfA5nWkfbnIZYLCC+/Qp3J29xh
AM5SUvYNS9wTyiYIbirtKequtCylPP6HA6ytVPkRunoHJSRsK5Zk45SRDreft1lX
TD3dFPpbKaIEaRoLFVoWFV+aMn+ioYKRycoh7zMsbX/rEsb2DneqS8bSspOfnsOC
PiAKowJhgE8RuG9bFfcygC5RqlEGZRqtpUiVupMd8Vnq0Dbf6863ax82HERxh2mp
sdej+z7zV/XzZxklgU7cXg32giWin1oVBR/N2K5JIsMbrb5eOPKkEjDk4qX9gCKW
2o2DoOA7VztvWGpjosWp4uD8xBgjmMQzl7Q3zNoWmF/fx2baJLFMmfriksCQ2wHG
wGDMnXljCC8F+0fRs8R05Wv2Vs2U7XSEtD20cwp+loJBdlV+4scvRbeXs3/vHaqz
NVpeazGPnsHORSfGNTzheUQHTNUYZaUOWbjsEoXSQS/pD2KZRmPMS6E3Cbq39Ldf
+cUOQtsJNuCohqJDVOa8kyXLzCcfaQRoNknN8u41kZYESYcJYKWjHAjXEMCEQfEz
Fi14VBWEZRJa2t+B9su+I8K/hxD0WyyfrGHqI3X2SQIum++VXr6vQtPcG4T2Ju+S
DkLcDbFath83xB9UZ+B/FYFQlTiYFWGRLnh8k12AhnrFHr9Hr9HyPEfzpRwWD+CE
uBWTN6HVXbBTBqvsL4o6X7DdiRhDV50uojrArrihQ+9XBPA+ZWWnHnsEJ5kwa3Y9
YlLBAJLOWMYClCh6vl2p4hecUuDUt1L8ckD8VqFtJ1mZJJ1iHSqwHxA/UNDlwn/v
Nazrqnq0WTGnuUt1NRWjO0MWG7KB3UnkwdiLvzbsd/4XSbV2NF/Zz3mcx5tC7XCd
YAbAaPvhAE3QZz9ID2p2CaOIAIWnXKBEM9+1TIBl5cTajt7bJqsYPDAhOIG7C1tb
d45hJYs1Uaki8+TuRrFF5B1p7vi3p7E5bugKqjNEerzOsOWfp/blHdnV7O+AslQk
8Q1/RDSJKcaYWhM12hSqO5b5i4/wXK5DgGDKMKG86bqcEBAkW7+VxKkLQIOOZp+n
iBwLDZwNq8CSYZXtqYJYvfXHHOT/jJqpllUu4o8DSdXJ2CvsZPKS7Uct6cFfbcJ+
plQJJuj9j6b4w60nO5pmgUWE11ZpQ3Lpg6JatTgJtyyGTDZzkh6uLl5CZc1tGBKR
nIC1KXZxatRyozpG7e4xVCSGbxbqkeFatwg8+6Ee7+oSJFXwmalCUzSaCYxEa84i
bnWHHO/XapdeH9XY4NHkifOuuauwVmMJP2vZNZ7lIh1l3SVhJnHHcDQypNafH/ot
ecybLRlr8r5z/q8wx++UYYKzmMImk5AV7W1q8p00EVrI2LKMQgm0G/1jO3ymCTgF
vBwdbCCDUvy5zFRD37Jyh599CcSFIZin0PyyUrHhPOE40sdV1LrtT2p1c9jdLtiR
/s+6JwXvE1Q/7/N7wkuD6fye+vSQTPVoZiZmNgFANb1lrrX1kfEEP3R7cZVa19A4
H5ISqHngNIYlShdkCQ5IF86xdvPuRAr7aSghSDTlM23dwVMDSThM4WT8xZWIZ2NQ
YeaMM8EAzN5hwbfQ0GGCcWyjP3rqpkLIkopesrWcLYRLbIIGcBst2QOuof762gOc
/RuIQwS0wY9REQXr2w/6tQ==
`pragma protect end_protected
