-- megafunction wizard: %FIR II v15.1%
-- GENERATION: XML
-- ddc_fir1.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ddc_fir1 is
	port (
		clk              : in  std_logic                     := '0';             --                     clk.clk
		reset_n          : in  std_logic                     := '0';             --                     rst.reset_n
		ast_sink_data    : in  std_logic_vector(23 downto 0) := (others => '0'); --   avalon_streaming_sink.data
		ast_sink_valid   : in  std_logic                     := '0';             --                        .valid
		ast_sink_error   : in  std_logic_vector(1 downto 0)  := (others => '0'); --                        .error
		ast_source_data  : out std_logic_vector(23 downto 0);                    -- avalon_streaming_source.data
		ast_source_valid : out std_logic;                                        --                        .valid
		ast_source_error : out std_logic_vector(1 downto 0)                      --                        .error
	);
end entity ddc_fir1;

architecture rtl of ddc_fir1 is
	component ddc_fir1_0002 is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset_n          : in  std_logic                     := 'X';             -- reset_n
			ast_sink_data    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			ast_sink_valid   : in  std_logic                     := 'X';             -- valid
			ast_sink_error   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			ast_source_data  : out std_logic_vector(23 downto 0);                    -- data
			ast_source_valid : out std_logic;                                        -- valid
			ast_source_error : out std_logic_vector(1 downto 0)                      -- error
		);
	end component ddc_fir1_0002;

begin

	ddc_fir1_inst : component ddc_fir1_0002
		port map (
			clk              => clk,              --                     clk.clk
			reset_n          => reset_n,          --                     rst.reset_n
			ast_sink_data    => ast_sink_data,    --   avalon_streaming_sink.data
			ast_sink_valid   => ast_sink_valid,   --                        .valid
			ast_sink_error   => ast_sink_error,   --                        .error
			ast_source_data  => ast_source_data,  -- avalon_streaming_source.data
			ast_source_valid => ast_source_valid, --                        .valid
			ast_source_error => ast_source_error  --                        .error
		);

end architecture rtl; -- of ddc_fir1
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2016 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="15.1" >
-- Retrieval info: 	<generic name="filterType" value="decim" />
-- Retrieval info: 	<generic name="interpFactor" value="1" />
-- Retrieval info: 	<generic name="decimFactor" value="20" />
-- Retrieval info: 	<generic name="symmetryMode" value="nsym" />
-- Retrieval info: 	<generic name="L_bandsFilter" value="1" />
-- Retrieval info: 	<generic name="inputChannelNum" value="1" />
-- Retrieval info: 	<generic name="clockRate" value="125" />
-- Retrieval info: 	<generic name="clockSlack" value="0" />
-- Retrieval info: 	<generic name="inputRate" value="125" />
-- Retrieval info: 	<generic name="coeffReload" value="false" />
-- Retrieval info: 	<generic name="baseAddress" value="0" />
-- Retrieval info: 	<generic name="readWriteMode" value="read_write" />
-- Retrieval info: 	<generic name="backPressure" value="false" />
-- Retrieval info: 	<generic name="deviceFamily" value="Cyclone V" />
-- Retrieval info: 	<generic name="speedGrade" value="medium" />
-- Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
-- Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
-- Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
-- Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
-- Retrieval info: 	<generic name="reconfigurable" value="false" />
-- Retrieval info: 	<generic name="num_modes" value="2" />
-- Retrieval info: 	<generic name="reconfigurable_list" value="0" />
-- Retrieval info: 	<generic name="MODE_STRING" value="None Set" />
-- Retrieval info: 	<generic name="channelModes" value="0,1,2,3" />
-- Retrieval info: 	<generic name="inputType" value="int" />
-- Retrieval info: 	<generic name="inputBitWidth" value="24" />
-- Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
-- Retrieval info: 	<generic name="coeffSetRealValue" value="1.38247945E-5,2.58330329E-5,4.21390631E-5,6.35768949E-5,9.10562604E-5,1.25559828E-4,1.6813907E-4,2.19908739E-4,2.82039922E-4,3.55751678E-4,4.42301257E-4,5.42972963E-4,6.59065707E-4,7.91879341E-4,9.42699898E-4,0.00111278385,0.00130334157,0.00151552013,0.00175038571,0.0020089057,0.00229193091,0.00260017793,0.00293421203,0.00329443079,0.00368104869,0.00409408296,0.00453334097,0.00499840923,0.00548864438,0.00600316636,0.00654085378,0.00710034183,0.00768002278,0.00827804912,0.00889233949,0.00952058733,0.0101602723,0.0108086745,0.0114628911,0.0121198558,0.0127763603,0.0134290781,0.0140745903,0.0147094129,0.0153300256,0.0159329017,0.0165145388,0.0170714894,0.0176003927,0.018098005,0.0185612296,0.0189871467,0.0193730405,0.0197164255,0.0200150708,0.0202670214,0.0204706179,0.0206245126,0.0207276825,0.0207794402,0.0207794402,0.0207276825,0.0206245126,0.0204706179,0.0202670214,0.0200150708,0.0197164255,0.0193730405,0.0189871467,0.0185612296,0.018098005,0.0176003927,0.0170714894,0.0165145388,0.0159329017,0.0153300256,0.0147094129,0.0140745903,0.0134290781,0.0127763603,0.0121198558,0.0114628911,0.0108086745,0.0101602723,0.00952058733,0.00889233949,0.00827804912,0.00768002278,0.00710034183,0.00654085378,0.00600316636,0.00548864438,0.00499840923,0.00453334097,0.00409408296,0.00368104869,0.00329443079,0.00293421203,0.00260017793,0.00229193091,0.0020089057,0.00175038571,0.00151552013,0.00130334157,0.00111278385,9.42699898E-4,7.91879341E-4,6.59065707E-4,5.42972963E-4,4.42301257E-4,3.55751678E-4,2.82039922E-4,2.19908739E-4,1.6813907E-4,1.25559828E-4,9.10562604E-5,6.35768949E-5,4.21390631E-5,2.58330329E-5,1.38247945E-5" />
-- Retrieval info: 	<generic name="coeffScaling" value="auto" />
-- Retrieval info: 	<generic name="coeffType" value="int" />
-- Retrieval info: 	<generic name="coeffBitWidth" value="8" />
-- Retrieval info: 	<generic name="coeffFracBitWidth" value="0" />
-- Retrieval info: 	<generic name="outType" value="int" />
-- Retrieval info: 	<generic name="outMSBRound" value="sat" />
-- Retrieval info: 	<generic name="outMsbBitRem" value="5" />
-- Retrieval info: 	<generic name="outLSBRound" value="round" />
-- Retrieval info: 	<generic name="outLsbBitRem" value="10" />
-- Retrieval info: 	<generic name="bankCount" value="1" />
-- Retrieval info: 	<generic name="bankDisplay" value="0" />
-- Retrieval info: </instance>
-- IPFS_FILES : NONE
