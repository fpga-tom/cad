// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gQnbA0U5kse/sJ8j5hcEGgyrQ1lGFy+lijnn3WpJ4XBai7qa3yeWpHikeboppcyh
/d6ZtRKFDqWUR//4VvUIcQtdO1EgoT+8IwB8JM60Jgqz9tazrOnysXIAL9+FzyrH
4dOatjKsYTP5TR0Jhx/lBM8//9m4MRIWt4XRa0W/Ixs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27600)
LpEwpu9Yd01+kgJVPUxm9wS0C7b0S8FGnirmOBzh6viaGY015iP9ZkD5Vd4NbqUJ
yK2BcpT+K5Aj5fAcnqwVJKH2c6CS9u+XVajpA98dm4CNffoyCiH6MFD0QwLDQYUs
VAdF33NktmR036vEGQeXbMdaOL27Gi2y8irjNxbT5ixtnAp2dSanUdkCcM/QwSQj
bISF+R2aX09Q7PKGksV3ga1JOX9Q7Aog4H5qtdAb10YGdvFzuVOwMH5RQbekuaoE
F6OvUe8qjophWphUhn/26/jgLmHf1lSahJnwWhx1t+E/M0Oq1U2/YAPacyJ8hovh
sz8XIPUZlpsgQRebMo4ro6AlqVT4Jk1W3uGE+h5kQF/BLJGz1Ismi0ZeByzxgO2e
cQqBLD+xyCo4StBRml5s0jolIUBSS9QNz8IssyUUrrKJtBMRgrRgnjX+3aUGZ/O9
9gMv/wJ2J8eAu8hrKoI1TaeD7KP25ISWk0iSL81ZM9wajyWszT+gpip1AMkFgXwL
EeAobzJsKp63saOGWrQo82tgLzOeXcNQg26hzc1nZPXmbDrqBH0d0Nfqp9fnmwQV
xmmh6VNxTqCEz67J2L3eeL0WQXm63+vxPCCibyHhJnrZ/S8tPU+ZkeSLmLKVkEac
ueTcg4hhEHqI4lx+S6rTXxjv2YIvsQ7T5bIYc9wDRxdXFJ2W64ORw7x6A+KUds4X
o71Kpi/i1DnNMPHI6mEc2IyChdULGKgAFYySe6vhBG38YVysi/gQzyUxWq/SL5x1
JsmXMcEBJXhUngD3w8ibuPtQikKINJ8hW55MB9+cvkBQS5D+7My5XnGced7JOrtG
C5DDjnKlvw10ZspZSnBAwWHZRq6PVm3K4srsuX4QlgCrtmtl4k18yiSbRYaKog6W
yWj6U1LYZ8DYqqfxPoUeXgoy/0av+kPGnBkVTWzlHn4u/QIADg9BK1/RNE1S6RhS
3GvEiyYOK4ad3/FG587sthh/peqfLBE7yV+SlAwM/QXeN4s6RX/BOAxzZAMMrVpu
H0GE7otJh+87QQlQ22aPomu8CItxHbjRvoLgVHR/x2mxNHNTI+R1gbDLKWbmhGUB
eVkJZPGmMBJ6pGI+GhR7jm4yN0DGpRO/LD3TA5ptUFISuj1t+uaXzYMcC5IrFBk/
psu5L1cYhVai77igBm9CwDNfOlKZ3kxObf764cGvV2buaCQunCaLyoJw0Bv0UFD2
hZ189YRqDNiTPy0ikoDmch2iWZCkp7H+3+aMYIn4CT4qsgv7U5mLR7TsPJIoNcoZ
UIvus1K7+4gBmRvXI+1YOPKO4tIzTIRZasV+vbOI6tyP0xUgVqlQWkqIFHkYNazU
43CNN3ynMDvg0UcgJDHXanWDYfQuyFvsP5VmKLg8j3+veVTxfrlVKCdB3kP/+km9
LYIw+vL727KnPK/UPwEDmQIOlaEOzKIvSJ+EE3qoV1En9oPpcKEwvJSYoS8UgXrx
K6I4N6aYFQBevqmXfKymJa6sKaIRM35VdvPqOe2FHW7iUx+/kiVRwIcZJkWm9FfS
cVEtpPQDHHA10b+BH2tddiCo35bzCUlcETn8axeqyw3mJ+zBwtB7iiahrRsNGSjg
KlUjvpuU7lNtmFMMb1hS4V7Pa3h8BpYJqH49k4eumRQkjSGgyoDpMA5SWdhofhsu
L0JnJw5ZU+aRIYBSAcABt/tQWzrjiZpdawswsyQMY3Fa9gOmCCn0BTMvnTgsADPr
i9AKq7GV0oiGawp8KORjjZDjpKGUrGOhGhlLf2+2hhRnOfGYOGs2ibM2iqdjZFUg
oDeKpfaOWh/a+WECFiuF3mZ3hKqyIH3EZBya4rhFsU+zfviwjUxFNTP0n+hnPfeg
epB3gc25prWsfNqRgVP7dsPsLXnC0Nti0YVC8db+sHTLS8i1juSmMvERCfcb6t06
lvQV6m50oHWn9irzvm760T7FEa5b+9ShGQcs4uNceM9BL0OTUAwMw0JbOUrg2kbA
gyVhQEe3nZZrW5p1VgtkjFzhoomTwYu5DCWNNvV63Ex++qxG4zHa9DtpXE3QIWBZ
e09OiPfgIZObbAc8MvdLadHBKNQUuVGisuAxsG3QF/L0MAFrWaBHvT9odErnh7GJ
psuySt65WCEeibvaGuA7OkAVE4OxXu08qy8Wg4WecPWcyJePaqQiGEWA/TGxq9eY
zFdgY7WMXndiFQO8lLY+6iGSQ0TizgCiYOj37vrleJyQAXdhgdwlyQgSMGg8ioIJ
x0usiQgG8xHvbqleWDS8sKC7ZiAvnd9+wSV8W1SktS4V29+lSKMhZK8bUjoivPWo
LLxjWUEXHcOAdisTFhE75Jwoydcs4jzwfMxZ2wgcK1Xi6LsKGSI/2yNXQMr0vL4c
nc+Lm1nLD2C+54jyGVmGZ+AOBQbynWzdgQ5cuMrz2rN7K1Hf0dYOoOQJj4A9gFFg
nG6wv+NFIxPgeR0WqbUE8AgR9YQSL5toIkhhpYL9JTc6PEnmxADyaajZu6RQFnhv
Zuxg9/B+suLesWx0xfuqZ0S5l7N/OSsW7t79adyGANDaq3g3pq7X/vh8w9lf24n8
06IIbFiKgE8HB5/Uh8MrP9CX3RlLCBE+GSc+OOIXw4Eb4rF/RdNsqJKj9/SqBBEK
HnIRVzBzmGwh+KUxuPK1vZoHD9omJHcpedQT8IpeUdEJHdObmJZ1ICKygr3oWebD
c3yRNOBESd/uY7vNtcqaMnmoOHvNwoa5LBVqn1ZJg38uO6gBFfF4+DL38lkYPaF5
Pa8kn2+FUl3w1WdFHCVVR0B1G6LG7dhWC9bdaKdYWwDABmnodE8DD/NBnlRSSlMd
ip4f/IrHn/555DvvmAl3zte//CTEzf4Ecd3+QTz6d44pCWnT36mH2pAFDsbYKH3n
H07TNOXEksFhrs5B0EVFUFur6JpTgV6CdiIw51sHiyHecXBqVHg/uYB25FS672XA
bZFWYh+vgq28vsHSb30Z+3ycXPMqmIurdxzAS2C9ee+2To6G/spLm8yF1Z3cMkQV
wVJdlr8ITVfb6EdV5ms4YkypsibJs0pvzZIloi9hicKkwyoH+DaOeGxa+wrF4ZSC
NnvIyRrG17kPvrvmRWOoYRt6f/6r+VCgexFauOBKmn1bP6S5Tv1PEJWdni1XQnv0
brnhaW29+n1Xk2pqHje81zU9486Y4cRYuAFK2XsWMAzHPyuIadqz9m9AyTxYWy0h
C2IX93QeM+eHoZqGa8d3VnavebRycEOXqVMyIgxROjS0KBbwwwZfLa/BCVx2d5JX
MaPlO6BnYM5mxc9sUoFz44PIcw5ZjzWYOqTqznKtXjeoJ7Xw6kXvDMdPcdqyg9ua
aQY5vOXgr5TcfZ7f5HENLsee/Yll9ffTk3xJiQTwIMpMTqCfu1CBUYkno/1CMnlo
IEc5I3csUEo5XkGMrkONb2Fu7FpeIBWswBYYzLqHcP5EA9n70u+KNprDig/6ACF9
uapQklREJq3iKNHkUlmpyhJPTOabCZakIxpejfosnBrHr/iEcHAJEHkBr0VW258w
W8vReTG0un+Iyej01FbBs7T2ZMnb1cOjKPgWo+q/lJN8PU9NuI9f2Smy5dBXfULC
wcBfD1ycB212gW4Z/78fhOhM+ntktgB3Ep1d+T7XEDSSbdPuk/IPMamwVQ6eKLvy
uzGRwiICMQDKWiRYkEmHUqJzOFx41ygUvKBYglbZQj2NyQ51G1bt9/WsPk4unLeT
EP4Wze+4g+7ePBlpYwsktRpOMc3cpOrTfZ4SNbvmtn5EUbWFNpD7znrZrGrFlHbo
fggEbsxBlfOG5oK8iDXxOgZJ58iH/vxfBF0AEW+Lnz8JxW2w5s0dsUF8jFAuX7Fp
ajHyNvWwvuwwWeCvWgem/Le+6+m5xYkT1ton4vNZm4VDVKTtgUQ9QwOlKBhZL7Fq
nhVTiFLPwHPo6jr4IA0acWaTjg+3n66linv3xW06SD4HVLj+Appwmlya2dAdLdDI
fYGJZcUsPv1Isf2zA5JZ7kCi6Pf0DOPkcnS4mFSofGL5D5NtGQe/l3BVAXCvo88z
l3ODkd3jqN73PkPISpeKlmV8ixlPwHSukXqThiFs9speClBM5GAcMrbZ/keK6BTt
WYFEz1g/R20yYjM2Pr06TMq7Q2tfsOVzckmOxt1RWZihesF2M4GFqebZWnK16F8C
GQf20USfR5eXkuc4pqvVv5BPz3wpB+OedDXy/az+rfl7sxONNZMUQabSMyb1FbZN
JCxyujTW/ZSRT+GmsMorI6Ijv61d7T8Gqy77TnPIKDVMXQguXgDRnl33vc5svecR
IxUoAbemiUIpsra3wiEryO7Xl0tkHVfT7NWSy8W+W9ug6ySW3iBNYpYwOIkC/rWh
q0QqqOIahD2Nh7WwTVShLkLfHtM/F2hJRF3HPVeRFifWjX7MIqTzaCU2o11Rb2I/
7yl2WyY3fZAPVuJ43E6mayuSmlAhgtGVfC2xCqauSVBtHwsPuhZfmy/bhc7MsDrg
6l3dtF0y2e9/TvWDTpf3+m+YSmxprH9B3ejfvDlUunoXI0+4J6USs3TS+TN0mY7N
LCzZghQTG9jy6L0cBnFovO6ik6AsmSYXTyirK3XeV0wDOzMH6hv7y2BtuOCF4CFr
YJ8lPSBwR1qxfrFT1dlv1UQASNRFxgUi2TpSk19d+LA1Lk8M74GzzfdsGcCYkrEe
XmhG9g0zZn6KpLIXkcsEsQbZ3Nfp6XVv/4rwmuVWQ2KPRHq/U0ZVQ1AvmKlxH3bi
roCX+709UnHL7SYA0xX/fu+WNMIl9UmpIQMWZgSjoxdCssSKKRfWePIplgSLqg41
cOwjJx5Szo1TawQrOar2RBUeIE5kRhPsqI/2DkscCOt4Fhh4rsMQjsRIwXIwUlpi
C9amTSHU8El5qVyU5pbqtp8PLUyz3ptg+SfcthxS8N7Hsm1Oq3jfx1VaPh+JdMpd
lbe+LSFN6nSMmpsF0j2b4VacjF9l/4S/+jaYry9kVKwkWBKVdXzSNlXvq9Nznmfb
dYEXfBc8kg20szJL44GNHQfoafDSlZ6dgzFRfZTqo4QUM1XzEyovRBlQ99pn4ymU
R0VRstG1Xy0sVvJECRGssb4Mvzdrc/j+A53BSw0FSOhnhhSEXsMhyUPZ/5UoO605
M1Gq+qxjwMpsOF139jv0llEI5c7Pjmj3houYaiAEDCq2HDwJs4I2c1FIGWJAE3T7
5zUI1W46qfIAYKNaKW+L0cpL0TZpwPakH1v09vbQIBMww00BO7df7qalvJLYHrXf
p21TkHfjKtNq/nJu6eu6uyrBccHAzUmdhw018NFp429TAI129FQmR9zMkCqx8maF
8xbBr08l9+Pd/NhpITEbcw4xlcNOsgMylMvAQb3thqIXKBANGMQEAN8CSq7cEBsY
xE7UqDFBFITK51QB8wy8bywu6MVxn5pBEs4WqA+PNPOK2ubgTRqIACxuS52UBp8s
4UY4aXyip5M/mBjE8oGqmWt7N5l7jAfRWOc3tVFDYWNrn7Ccst9b9Oww8D4AC8Je
mzRBDvg51R/0X+CUcz5K4h3O+AAwyXq16eDmqvPGAtsJvBfYOo+q4ePNmWnEEa2W
sw1YET5jKHhRc7iMHK6dystrO1AITlNkkrWWAiwrcgonyMbaaUHwkk0L5AxaCAVj
ZImv3llqfUTu0eUOivv2Jjexi3JbZWUDRchhuV7S3I4FPL3j40VETclENnMc2LQv
2pbYj86owfPFnwGCJzT4zVtDldwkPmfhf9Uf8jPM9Tw8pDnjxz/vqVAab7BwA+34
jEinHUjoCa6I7BLVlAQOA7ApVhF6J4BdSRvqJ/lUkUKQJo7+/g3nrz7Kdy8j2IgV
YNXNpepd39zE3h/6jfAclNjYah0JPckVXQLQR51WiyzoEmU1dHzGfxf1beeiwIDv
yknFW67GI3OxvaZ/unTBvKcsaIU8T2x/UGWg6HXEetcqYsBKDBQZeY31PI/qkAmG
81cAtDYdo+VMtzXWmHjO0Y9yMiGedRy6BJzMmTQaUdc34EhskI2kbhNYOOqdxfCd
LZXVGAPD8sgc0YnuBqsKt2FVL/iv1E+50L8m26CaA5FZOwScpOGwIBSkR6eO6wUS
G0y7a0swCPgRshcwGCjjv5+LzMOgdSALnwkmr4AzRKD7hLNnyqdo0dilT4NYiWOe
MTnN4Mdr0FWq4U2026u0YO6OwhJLmDmr22W6s9bImMN0/jR44W7pm9jZJVHMGwbP
N8KWHY2XUQ2eOMZvVMGbJ+Zoog5bklDav7vrLrxAX42I8QhMy9hwVh4I1GPr4RHg
02R2nu9Rz3WBe6N+fPRGM7zkYHqJApfma0h36wLttXduqHx6qqLmOdqB3arvm/XR
AnsAs//Oh+jspHaW1Q84sGAdlKSFnyO/MeQ2N4Je3VDIBIvZcJ8LD1lHdDtboq9C
ynUPBojrcTRpNOJ4xwAPmGKJOqvbBo48hzaFxhiM6/MDjxEElb1yC5CHNFtKzISZ
WzJumLEJSGz0zHnNVbVAVCnObjOiXBcbcYe6eeZoRQHgcRU2jjFWgioi0gtnQ5Tt
69W9Tok+kucExW/0Lr7llLRyHL7e9aV2IW+QBYO5j2VrHg5hHbSliAhw3C5KjlLi
FrhOUuCAPHPhSnlzMTvTkrQlM0sSnxKtV/oW3LevKwRBK53ZOVPgQE7vaVYL4J70
2+APGKtHXZ4O7b4WNPljRZ9oaOT9s0MGUf0sijfPDRaw/1/Ic1VfbMJThsZF/5VE
TpH6o5kfXhTl8u1GC61urHV56WbK8ajoWKDRbOAfQA4jvcK2K1WFE3o60n8BxeUJ
aoKmHxbpMyoVOZemnyqIfdhv3xioun0CgavbCMeuz3f+jb8IRQmtJH2e4nhMwTg5
4JIdlFy+NKXh88FO5SAH4AJdTEsFZ5FnOSgr6vvTC0vT+ZpF+Wj8x9bc0gpsti9B
RPYxc6hq5i4I35J2nTCPqBsojG7VbB7v44JJ7pHGUbcAydf9shO0T4T55YVbjJqm
Y7Vkt1zcCU169bH+FqG6ChGAs7rL/hIyjFGC8UMRGiyfXpEznbsVzfuZFasvrkFb
qzXA5EfIBxln5y5X0qtGGq/Eee0a0Pr+dBsbJcmFuHwE14/Wh/0tMXzKfKU2CcKQ
H9DIBJrH3q2tmvqeIGXAaeRTC2J7M00a31eouYYF21RcOxm8fwYnZvjLbOwyjBgc
/mhlCE/63oph1B4nVkMMU4Cf+tmMytVtAMUFQAunpuNhEHhENImyuSsaiUj4gSpQ
Y5K8K+8HPe7EToIfdKhX3DDb7pYxV/Cy6wsEN0RRj7X4azuV0fbk/5khVbbdJBbp
gJLCVSFn1JUKRRaqDdzjglPkzq0cgHdH1xTYCLRrgD7D9eALNeHi9TOPaQfCBudj
cgBpt0qxRcSrcKtLIsGm+Odqo3NGqgscGw7wD/viTL6ThSpyXYpNL/cDj5G6Fl4T
Om2NTmL0HIZRcmQWtq2kNzzx7Dcv1A7NOTlbf5Gm2hAjmLpfzqFL61zD6CLdI1W+
7elOUoDOZVPbGYmWUI/E+bkr4OtzsG2Dq8RQoH4Ez1uj3hG42YNeVYDap5XsbhaP
I6qQd9Hg7QTUnoehdjzuODz/PdAO7+KexoyMdzfUwqsRa267k4JdgzA5FH2Ima9I
IjFQuLsrzhBt5c10KG9eobUG52VtowJaGkSEYIDJmQdf+LKYEFCMM71KECCHnnkB
zjs6a5s6s6xnBH8O8CwfefRkw7e6I3kSDJKJBRjiFwiY96PrOc+PvKaDS80/k72L
70A4JQZNWbYTAbttmFS6agPUoCFf2Ns8jGecGiZY69kwuQe9SfIh9aJOV53fBvKx
wjKj3Rt5IuzJSso/MP5mV6baqQVVUPziiyiI6l8b3k0VvLtUTAtYB1EvPM8htBvl
0CMgDWwmIcGLxq7hZZ7n3/XQuWxxaQThf8SWQhknwsncoWfhB04NxKKYVYWMDWbA
iTNszYj70GRWh6Ko3Np98YRTVPPJZkrtnpoTEG+VdAHCuoNQx+Kft3k1Y2WY1c1d
b0le+kRhqBlmIL36QsKOJTQg+HSvXzzl8TC1apF2vxCgLayHgGSwwWVgC3ePJKrE
5zL15310ITDTjhJHpSNX7nuJSV/n669Q5YFWAKZom/JiYGoo6qsjDCXrRIl6iWJb
ZlRYOoTmJARunUekaRc2zq3RNP06YJrWodSq0wjCmfxyA3gcRzI5yepVclVB6hOr
JnE+PG6jKcFEe+nSEtAaG341MJKzSX7Gbe9h+7quQj4Y3n0JOIhySkKAL1Tcozi9
UObWUmVrWIB6f9YUcTdV5BJlGcrwdSu07c/YCQzeZEALdjKvAv6XVSfGhG28iQ9P
UVS+WAwVMAhk6oeTFH3BOtBdgzg0Y3ZVb81kWel7DU2suPfKoOiruSCK6L+/KRcr
I4TcUq8aTtHJZ2XMAsBnLwuTEWZkwI40/Pjz7HfGj8TuU4Nwd7oTpC9UF+2vb/0x
oNsjrBuQYmCUmPMpisG04H63GPiMwd08C+89LykNaBoy9Z6LojOY7Wk6pmMENe1t
0fDjuFTnd8okMfjKnzX+7pPeJjeEgDzCREsWjV8T4GR1j+ZpVuZfY4Zqf5kAeXMP
xvKN+BZuO4yWt9BAt8CYFncZeeQFZzwM2IFsh3JLtsvynFH9AizxupHeJzUHVVTS
ff8hRjLZ0O816lCFktwZioljnn9IYZyWyZrYaQbuyTZw8ljBqtSpVDhHCBkjbApC
i1qAWTugovtVUtCvrP/rAqkvFsyhHCHdmtSeJzpYg2WYk7k06ShO9M9ypvlw/cYw
SbdUVAkRqgV/mDYD14S7UtXo4V4AQXBcE2/gkMl77veUQE3S55tvYqLuYeblXPmd
ke/+3cA2xF5QRb9MyQxNSHaINTm1i9QMOvFKeC17HKTCGS0TsfadLs3r72Mhurdl
rA218WRs/iJHfnOYmcb9EKe2j1zdSAkvQPVtKjtXuHNRX+shjl7bZWQ342aq0zwa
Y2U4gZ5iMAunKFBjQp0SZIJWXfzA5A7XkqSQAI3sPdyvgkruZA00p+SpjK3X5X1f
za+yC2hvQ4Xc90A/3HV7/mRKwwpSOuRmy0jPMtR9/jWxCxDJeV57uDOkKeERXkGY
I9YB2oYSE0naG3eQYSuGiJQ4+1LKkxeo8Ht1vjH3aK5Sac4VmdG4j38Qg2xsOuPn
Lw6b4nc7hpVQsCaSeDyjp0NeCfaIA05FdEQx+KUxiJB1sJvzD57bNv5JqVpgJZMB
hqWC4OZL+yw6AsnEVJEP5/lwfeKMHl2oxHiTSVhvMWsnqhmwQ1oGCgAlNwN87CSt
JWroJN5lK/GpTH4qQXSTMeTk9f6GrMJXTRlFTbDICF7Bhj81fvXjQ3zqc0NvxSxT
26SS4ca3mtsKMU1Q3Fu7Ge5l/fybFi0eXTOp1anHBUw1GhoFM+GbNWMBVpInW+Cc
W2B/GLAReHYzwD/gQ3IZvnLgZ3JK9XE6dClSsuIIU8NskBys3bDMG+9tav9C9DKS
x7V/mrt8UVa2BiDRtEQ1QHfxpywxTni46PB1ywxKCekSBdzGKvgfkqDQS/EWhy4q
T+pvJy/84uSTLnN7o9XIuAcBiGc5Y2J/ZQazbmeAFwRD4gf4k/JjyAIxYjvODON/
pH10QumTKQrZTOFakGtBQG1mmihm5fCrHF/dskYevSP6zu3JAOUtQ5QLm2wSP3zy
ANgRUJwUSIMxFS81uESrI6cDRoFs5/w2FqOck8KtCYfqQda3fn3FJD1qrr8Twt+c
ajexuFvNt1adWS7G6WTxN5c940HjP46GYZEyqd/cNH3hhfGDoieSAxJlLnVhgx0r
xzFCgOsctAHK7KLs1Op5hZZgoFBcIhcom0XdH18G06in5AAIdqLJ4HKjGnD1RySU
18it+cfsYmRZY6/wzi8FkR4dxu55TyMYWz60ZVPR/HZ6o3Qed5rKZu2AoU04g4zu
wfp2wcZPtltwIwTLu+0Hm/fNGXkf4yKwXNdG3KFog8MUnmfZlTaZHdUvcmK5Vpo9
ViiPdCUHU5M61jBq4nAShgynQOCci342B9ZQLujgtk14pwB+J1qWHZM8huGQrZqg
6h5+SKFGnO6EAlUxjObpaL0ruPKAsIGcRUebxg3qHcEJ+ystHy7G3uXqE28t6KTB
ous4sG2aKrqHYoQbaHcSfch2g4t3uR/uNs0PndxDmlr9b2Krzn2nb8YxBqciw/Uy
DzGDKnWBuaFet/TE0W6iSYHY0qQnXMInGh1rH3Y/q4CjQVWuKY91LAxWb2cAoGoo
3ByxIJSFjw0LYDf41IHSC9KFwLwFQnKmsdk2Al6tGEX1ukpzMkcyiQdCuXa5+4J9
574NBi+m+WHSqXM2Bg7CL+hUXPl5H+tPIIWyQqld7pQRsOhDtlORQuTv4azrYbyq
CKeKZSA7wVXXEojvfproTzsBFl1RQ5Ng2dQFL9s8oOXQGZbuF53cUn9fh/cUZTzD
727YOwWAGi/f/Y+hZOeQ3v04LepOoItyW/lJT5IAQFjtpcycSNeePSUz6ag19Cal
jqclzm3086V1sK4hNZJpDXhNLOgkVbdYD4f86CWa1KBexuzfp2A3Ss6FZ2F6reV1
DHtH0AculvLaxu+rXbulQ91hP4IquyFzBtPluEk9djZO2Yr1LU2yt+mdxX3LbQbf
gm9QPorGT7cQ3iiN2q74ab0f7fPT/R2F2Cyrhqhvb9zO6EVln4INX9UQmKigSsDu
LehpZavA0MUCIyiiybUYLBPRTbLt6+frPlJr7O/92yv2MXZeyP2M3RerrVcUlphP
b4SOjy88bE9AqrDR8q5dyhWQ32wr+InbXD2+tVHARre3n0VrIRVBPc7zmQQRY3QL
AxeoGhH20B1+LfCn0eCryM7IdEpN2Lw2zA0TrelmDJzj26GTol8Cc9jR/2ZukP/o
MzZsV+CjwWzAbMB+91ahzarze8ARb7MRciq3yBTniTqnQgiTVdRMQSCOPKeteqgO
S73IirGSwKeRkLEytJmDlq/K0zAGxdjsX6DhrMvBLkskiITa1eEMBl20TZvP+PCX
rExes6Lq+AX5bzFNFzYBBuhOl8gVnbK3TkuQsdXI9xLz6GJUWIW5ziBAZO00pcxh
4U59jToe18C1E0d8vPsAum+l95XFg3Fr2j2993VtLXtdgAaEZ4067ir6H0cFJo3H
JAzlP+iKYiCHBIYqLYiir2G33imlcbUcB6kY0u+f6L+jioFE6vlFlPLezj8R8Ftl
7xq61LRY1vUUA8+tchP9VsVN3B6O4Z0mk/ho46PxF0irakuxJb3fkP9Egg4ScP+Q
9fcPUms+tfgXMieJMkSLQrHSWaXseVZCckYKb0UQv5I2fZ9w8etFUftPOWQp1F0C
4ybJyNN/XwfoWwjwTYhuWeQVT5UD4L/njUKcd6TE3bYJrVo5yMksudwFWgeulhFS
2LYJ3l5s51/Uad9YOONeOvkJE/7H7G/R1KblBRTAI5cHF3dq8oJF3VX3cBwcEBzj
CESS+M6QTp+4WAUsZqhsvLwNKCYIP7qYs3XJIhBc3zdOVIi7zgzHH853QPL1ORW4
gF594XJQSanOpNI3thd7wTLdUImVoeF+atJ5CoYLVv1oVechNUI+Yc7SM/BMzSh2
lQr8iwUSpTSsQJ7N0HfiGsy37p9L+qlwVfq9EJ8ExHaZeQ3r06r04TxRUv4PZT9Q
ZYDdRyzAe9Ln573iwOgaSulY0/FGZMz1WCwQ/S6vlLYW6Y0nCVVNQB2Omo7b4kNs
qyfmuaylJc33Z+jwzUyIsGZZlIskLAgWYMqLZnuurLE/L10ln6+RzZSW3GTtyukO
687EEmaQM/0J1Olq6vHhBL71iSkHaFWqDrPD4Wjx62tIFJBVzl8qeXFgvFdHGWxI
F4/7nWo/1vyXs8WqP7vzCjqGwyjxezFCM6LxlWWuAnX0ZBjegXkQvcLl8qbygRLd
SXx4n2Z1mRZpEaJ4VMHQtxF14/11O/2I9CgetHOI41bhZmO85zGpCOoGFs8U9Yhw
Kkbh9RgJeQPAX/pxj5tj1u1vCdhKebpasPdP7khtN7FIIPC2NulWbgn3rlQLDmeO
Hz51gZW6YvyAgmkmVJq8CfHQ1wcvYLOCSykCWyGFpSGsojtK3sy1FcuZ+yatxBEY
mVwawCQqU23sTohC292LigBla/ccQkJchwpojov86tRCiN/5fK8G5M13UfIQzYkT
Byq7r0Pz8esVmmJbOcjHaZtLvYNc6hJTd5kFh0RyswUg1UgloNzZL7e+z8kIBWWs
GDOh4bcCZ9Snkthi9VBaoLnpPnrejqd1iJNeWwCZKTpPSjV4tJ4Z/kZn7t+RH/b6
L8lL9x2nR5d63vf5O5T+2JXSP2pHTWv2FaSZCeLQ9jDFW6P6C81ET4hCl6MnzP9t
awDvnPspZ67jUQ5Gp+S65C2NFSOTN5g7MnZx3wgET7EBX4ccq0R7jbd+5k9Me6pE
KyUnw7Flr1f3N1N67qhFczVaGkPABiY2t3k6lxTEbs2MMHuT82evnURZE56BT+AW
MbNpUmHIokZfNqXAtYVZPbO9zLGQVmDMQTRPDOUglla1TPWAhw4EgEQRrMN1cVom
qmZ9sx0eFuSY/+XIna/cZmwkGT3AZI2k1owod0ImgmhbNzslQfCuv8A631/OJiFu
K/lpO5IdT7c57UrqBZfTKLdcDIQkYqO8Fo/SPU2KaOh1AGbu7i9D6ktTLEkOCXNe
UqrVxkqMuU79ulMQxg7XdNd528txQOmfmDSPI3EdOY/z+acoNrcAqBgvziFzz+df
YE2ToKGzKB7Cw+1FZkSHBT9pbdH6E2/t3syKQ2CQUaoWKAv6MTBhu2CjjHHe0d27
xciEArxH49NCkqNmssAus0dY+ujkUc2UiWG4LYeZUM5uVmSjK4iWH6RNuVRAcdRY
ctqpPFazAp19wXkRdiOztJKVa6JqIXnWECBjxBRLDu8WOyyt/HAUxkXW3EGebDUu
0zWCEst7UbDXmKJsFjIC5J3RlTaRfm8DLqrBKhPSSnQUiAPnMwlrkpzsR8deNLTx
opgTYASL1n1KrKZYrVKFoZao+bDjTx26jLtKCDMEFFBZEQIiLqSlgIRIvFeBGGmI
2NdNHmNFb9SvoRgt+0sdDHCMlUrO/HpfqldW3J3kF+JVUmf42diNsj6KAej+h4/n
q0d9/DlhRKEXKr/PYMY3xlYE9eBkf9S7wFdWwzcM2cX3bh6vljeuJA03f1Vrm75q
SKPz0AKWRPenGkbZrHmXxClifPjdy0yTa9JjhnNn0RwrQp25acjL/M7zRBnIRWj+
j9aueILNncn/MNFJIhitfMo6fRi1JQuDK3M7qpeFexKSxL7cLWaxG8tqOV4zPxvA
x7A2iaHl5+P8NyOMXwJfSgzGBYGCLMtp7x9V4DC203TEidbOv61z+R4/pfSj9dul
0s8VNQZBuCaW+3mTwG33MN3DwqGFgn2phkxXqDlExN90rpiC9ansKfrPeHsZLjdi
VVsKsb+87nQU1w6N/fMVnEzhJKIUB4N084AGTcontIwM4zgEGeR9JYzlvOsFUG+h
HDKZAHO7cQz9VpGLd9+5V86uLo6tNDqNJqbjKvDDtmzT7SuUEpLtuWfUX1HQ3OJX
dWkWUUBb+rRq6lOOYmRjwwQ2vGsVfwmquVSq2jIK0K8IaIfxa8Zh9ViLRuxAhPa0
sO8hi/hrnVvjlvaw5DuJWNMyQnmn1jJnUmlnAV2XOkTjl3QYnkKWG4EMnbl+Qnml
ajtp13NWNBjLGE+ZlkPloCiYt3ceG1UZKGy7tJSopfaDSKdUB3Ub4OM7d9cjOrnu
S/0FmiqcOcpqFiLsTCcavtEcEyhUpCg4wUewpxG1PWGqwK1dT5c2vmEhgoZMwPU5
kyjPLJgMj2gE5YZpeMxghfeF/oAtdEpnBjr5WGhLy3cjClQodZYJqUtuNmdf9XcU
WCCavDbigLCpHAsGABs7K72WvtbEZNiWP5oB0WybnJ3Ome+8sukvC5hLZ/Cwgqw1
au5Dwe2aQyDHpUz9/4akYnM72vaNEfUqK6ki2P2BMSknyZV2NbZX3UFL3WnFuu5Y
G73x5iPZ+td6lSiGfpmPBOcbZtiRm1iR5l21n4rnv7Nfp9hyAsBhFtZ9CJUuZShp
FVgZhYFobdEezxgZQFjBim7C2HjUGgylFD8PeYAJNY7xoQHu5x95bMZpc7vaMOcu
W27nVEjbqvaCHuW1hhTsgDQdf8HrD2XJ4sg/UYwVfOtp4hPCh6C3g3HB19nsmp6M
iIUQRFYbMOUd8O+5+FL/ae+40lzwkE7ifAMVeN3cBlc4FT0iFGogjEchU9cDJGfR
ky05Z+zx/4DYYzJrwJTvCdn/ZDjkJVoMFICgOf42/Ppq0BBopHjVTifXMy/bCA2J
7oY9o4wwCEMhFllyhkQAqAd7oyFcFcdbPRrYWTPtYK0lghkeVxa+0eBaabLeV9PM
jDbqxfB2eZPlriTbyyRoBEW1VCsr8/ffT9QY5LyEgRfRevweWMiZONeSymJg46pz
5aSPrs/zfZTsLzf4rf5Am/LoFLtN3Ik/NLbxsGzv/ChmongKix/SnVyQfSynZ4CP
Mbe6KsKQrJTQ37KNWRMnjJC4lXdW/pPaRA4nVg7RUizSyCRFFqjxciMKsU8nVnBm
PyC60aiu1yKRmiFRCZcFpeCbjHv960fVL+Hknx54afaOhqQ/ysj7RxwPj+8ZaDlU
n6mfm01VoCki4TTTnDkDUp6MUibyTDyvx07DhJRDC5MYNr2mw8uZg1ztgVxiBmVs
Z97zOHL+n8BoFPPYvhLR37GSw9HTyUkOrIudXMbs5UNd7jhYjzTFF+RZDj3HPWyp
dIBwwPr/3+lZta+8sOONScITg5+ECP3F02pZUW2xk9q7INyB+YxmrH6dIPkcTfv9
RhE5TpWdxNxt88uo7TE/qveOIC8H5swrP4rxTof5wOOGX7DLdJmSr34aRpKr6DET
/lM39WQToX6ddxJfCqqbVARgItrrwzzQYrHYAaGfEZZ0N+9juIqnFM5XEM68+POz
kpZ8+sYnInhfwFguQE7Uuz2P7Xysgfh6mrtuRJiP1pCns+scfYx+Tq/LFngCeL++
ZvQxC9Saw3Dpsp0hT5becjey9Puv8L6W/9emBx+hevepWRbzqHJfVrnY5tbApY5w
jzqn8c0ZWEu4z1LHdOQjUU/RsLbzjVY9VULdhiTQBhPlz/lwxEsxWABQ70n2lU35
z8L2HXdZqRye0em3675T4YVA54XSfrMccEa/fTPVm3QpbiySw7yrAWVpGLjgIwjq
M4IY9UDu6Mpg3VF/of8/SAbqY6GOofqzLQuTefazcclglp1VPbIiVc+mDDapvDMb
LzNeMYaI9oU/qVuoeyDJRaEOpCoe165mJbURCaxKEv0fffvgC5RFUM6igF4K4uvl
Yt6vXtSQBbpq1ywqWZHTipi3o44N3xg+rk/C4jkklNRDul8BwUkE+FpB3Z53Q4e6
A4KWYGzED5ssq2ICpMlgRlvGJJViElZ+4eSVaxk9WiH6Xg0iwWVK6qG1gxc6hg8H
doqVYX64daWHwoOaBOllzT6q/ZiCkzOS+1XJt1u3HxxD8D8JYJSaEbNEdLFuCCcX
sSm9J9qssIr2YNcq5nnnNb+Zx6pSePnJBgrPvEYPrlritLdnsXRo4PYmaq3zp7KD
lYvsoWmd3fE+KuGXPMNH53fN49CskYZQzypejJLLRONHDDzTIhazI469A31ghnDl
hIeiH0TndmK1BkH8dK+N9E6BPRgNqbqBE8eDgkpMbujIAe59kWt5d3RxJKDQBAd+
Ag7CT9B9VpCwomI8yoIAq91ZIIfeN5vR5MZYL/oAfKtEs8316m4sjnnZYH5HtUNp
iXUevp2qZLEkgnPcczCfV8NHtIYh316qYJePwg3aUC4wStaAdnpq43cOClM6RMCP
DWaDRTzmx8Y7IejujrUtM7B0cKcDIALHy+/oZpt19XzqO0lQ/TxAy6vKF7QgQPMx
aNIHhzphX4SywqdgGq2Vr6aGxxbIL7jlGyYtbXlLZpCBM2pnln+r020NoQkXaQmZ
0dujeI/sDNeRJYU+iFrGdFCkzFoxu4tB7hqUPmVsXiuvjP6vnP3bJ2sWn91lEVW/
kU55DWeE221hO07WUPXmiSouDkQDZudFznsaWntYELkIb+ii4BlDF2UUHo662Lor
XdjXFoUlNIOi/AxfEDALCNlt2C8mub8IDd05akhllH4R3ZRxWunI7kwc7AnR0F29
wDM1nl7xe2EbqgVF5NYTOCY5xXN/LSXqY5R8hTNZx3A489fccH0dhQ5XEKpp8FA9
GyzjEjslxlKCrcciFwtopztLIhoLxuB44yCrBYoxMBDD9yVQgScT+587oRxtm53D
JhGMCC3BoWZmoAnhPqWEqnTEiokokqxNEYBlIEzwoQozb//lOGb0GgC+A2Nv4ade
k8rxDvkvwPFk8P5XRpBHgAgoK247QH6Nw2tJDkRkL6r3/c1gLgmGGxGl7tTsXn10
VOJzb8y0CZLo4/LjSMSnSe6kYVjGivLa2he92O7YMK4Gbr/7/mCpiuk85uRC6nBT
yqhY+2d6PLCBmQXjbJa2EZ8j6W3mq8yZ8g4Xey1SKCFmRb8XM8Ee4MlRl4+P8QVA
rqG49QmfNS3NLElJ1Lbht0+XlcaBrEGeXx9tR14HZPg4sUuo4/qlEjK04iFC17cN
vQbn5R6aokBcJtgRf1Lap2rw7/uL4cLWQx/LhG1a3dlCbkB8FuAlQZR9LkhLxW2/
d70em3f47wNwgX8Soj/v16/TLrEDoyJd6bDpA4AypufqTGYQ9E5lv0f1grzf/Djr
SFQO/i0Zk+APQnbaiZxFvO7qeUhuoWht7gyF9fN5A+d9ZFZ3GyN2C8YSuXbBUqak
1oseDnofm/HrpP8M/61apyUW5uIVg2WYvaBf1AcEZEWK1k1CTPvJkd6Iw0P7LnOd
HtLanKOXHCj3IOwnbaHjLgDE8/1L9rMankNZbhOdsSlXmz0V45dtxxJY3l5e5iZi
1gySWo0/lTuKqk9fZmXGlS6RSF9MvtRjVpC712FAlIA+EGFLpUEb+Xf0cV+M2DPe
h2W6HPKnQVxKvNx3ucVwfJwUugy79ftHaGBDoOZUwKC/g/RSq5GyltH8JZGsAVs4
Ka+u8R8RJII4JjMvXaM/CGUX1BwXh14p6bP75uME7/b8p5KH3z9bz1HRZcHZrQAw
Mvbp39/s6AiUNRE9E8rfcnVZQSTLFCSY+edaVBoCYrfojYHxGabG6WPa/dVgriZ/
XwxnGYIoLDAyc+RdTZFLZXqDtzZ0ZgJ2ICaEkPKGVn8bjrtvBl2WXxim4Oyhvo+Y
hFxyxdogDb2gqhJ5ienLjCylCwkA+iUoMqg9CidCxLeZVzZdqyRU9CpOytVB/zvM
kBD9NpuktDwUJTwFrSIwUiZpomlF28A5vUKPnoeVF+Bk8XpmU96l4tVMMm06yWRo
xVTceM024L60XeL7fL2eyvE1Dv8udlRDetM6LUpgX2TQg6J6syG4kM6Uwpi41+YF
qvq3MgpF9Es84RuYaK0Zf4YzC6yFXc3C81Xm37HrCr5toyEOEdUhTyphrBxEgE2u
OQ+1o67zd/H3VnPVopgygBnMShrzn3jTS9WmLQHrT1FNDHVDYFfjmzY0aIITbzbo
EkQM7EqrjQ/PFTpHngWSx26IuTTTtebtXKkqHM90N73REwHGHna7gy+bCA4oUaYT
eMwFknrXIPU1tXw5haHexP8O4qwHA2eytWkXAIm5HLdFtg0l3k5Zg7LhUYUD9s4p
40aDvIBc+Yh4porDH9E56soEL+7c2g0guJtWeCoqwJDPCrLA1S/IhrPGlU18EodO
p87w18LcckNvB0Y7+jYr2PgfNKnu4/td1KzVYstow1s74sw1rKdkgRB9QZto7j3w
7h6afkZ4jbJB38oJ4aCK0x7oUDI+vMtrISeOHpS6Ma1t9Jey39e1miuKZZAJLQLM
wy93cjSar+qWdn9qnVgMz2c1ilQ13Lr1EdjKo8PFKXZDPsfI3GoivmEinNBpacXX
TN4kJ3EIs5Z7bk1eKrWqZtG4P++K1i0eg+T0E9ustWQtdzXJrGpjVYL4Pu3GO4sM
vexaPDsxkVJECKVKh7yWSA7H5W50o7kUpjKq9en171u5XMHTY4PGYIpVlCLVKq5q
n2Y1AINkvi4XaqxRzabFonu1cdxXw8aJoOwsLZ9mkcUI/zDb0RbJvKRIqpeYXmZL
xOXPx5AxRfZZCiKtyYkhjT0n+NCOnRkfrWgEl9Egf6mZv1s9WCyIpDxx7ieit/QX
/FRDA5bFFSSX0iA46YLJ+nUYwqMvDspwfDWxLyfEIxBBERlqaOBU/ca/k30sUwhu
Dmq08xS7jTdGjtU6lXgNS/Beccafk515TYBnYMj8L3Wl4EOKNWvRKoA7pwPD6yEs
xgnn0HEMqRvrJ4xsmAtH83fCkYQiZPVksE5AqT7XRn+javb+vf/xZ3dOvmUTyk4U
QgxHjbjS4/TKhDZqzPaahZrDJB9u71zwWXAflZfhvm4bxR6ZSuE0+5HcX7tIpyo4
eiIpYcoV1VK3UP9krnWhuY/HpfGK8bZ3qRxp/VLFasV6Zf7x6tOTVyTs7O7WzBWW
yq057uBpoFEcI8/BEKyEs0E+S2k2jNfoKT/2TXrthbGuUABk0o+Dwj34EhsKnb82
TI8i7eFYEaTMWQ7LCY4Wa2omVp36YX+g3LmopyF/zPy4zGgcTarPUiC5EVy+DgrE
qqHovKtJAIxW3w27hcipmhLMbakL7emqW+UrQweoAm+SDfZUgP6en4/FzpprcLMg
Ox5dlg08BhQt4Cfl8QUjOP3wTnLl534JPzb3j9hzDxp5RZQuwmFcWIVDomWzcyBg
/r/Ko/FA7Od5r+FgwO3tXmci15qImfn+PrYiPZrADjxjpBi6EceZIbYd1Z6GQpgs
ZPriDgbj7DhGCXCfX81lIKaPleMe6drbNVbcLFXxhTyCG6N5bOcRNoDBczWhVBM4
sBtMaTlJh7neiS6DHP0TanSYvEOcZPO8U9gRs8yZQnVkhLM9/bX5QaVz7R/6yN2N
e7T6CXqGcCyjQRYRci/F+ek/pizbUqU0Xa9yhbf7GV559gYN0b3dpXYe3gU4jq48
3h5QBUH0xAUwjnFYERy/KbXAYbdNBY/xx2lw8x5fFxf6ag7WT9p1bjiWjd6g3Sfy
j81yVlGJ6j38o1uMIdPZsNGGCVL0OJOUkdt3YXfVFyu+GDpEuBewjG6yufYVa73O
AWIsqVvUrOodlEESxjVG5+JNMDufvpj+f6rV2RSS3+y7n+BFVn0bMah7WXrBDwKV
JcyA5gxeHf8NXXoN+yMHR+oJzuR5DjdRfs0WYcbjpTnGQaGXTd+qFw6NmzJ9o3oN
RsPO1vZH1bqYDLuA+M2xydN+MQI8kyLV1pTvv3HViVfPo011AsnBSTeu9tkOoZh9
LmoW8UjcK9fUteEvu4/G/2gwbHy2sHWF1gBm/GPlM5Cus55stn9zJa1UESaZNse/
WFrvTqWNCW6m6ss12vI7kF/zFj8OWHn9Wu/yeFJU3vEoyIHj7hDMguPPTTz7YyAQ
2X8XZ4d7FshG4HtFsregP6x7Mz9+EDyDya3PzMjwu9Uc3xpfQa/SNSc0wCZNmzAj
NxT0mdyVilj60WMBbif3PfIl7hMSUwzCiN6FL1PQYl11eJcQGOjeOW6Jaa6MLnqt
VaSdiB+fXwwZjYCwI7iN5tbmlL+BmX1j/ccjEdfXZeaFceOEILyqtFeXKSerAJJw
6WDu1kS7MhYy0P4L8vVt2PxGRjWWzf1booLXGjMcfBLE2tagn14kAxKLaUF0MY3E
LHiszZysRvA+4jZFTfiT0VU/DQz+KSiUMisgbNtM7cx6U7fq0LPio6RRYYM5hXRG
D4cg35J1alxwSeRNZwxYlR3PpoSI+Fyy9GHeD2Xaui6nQeSVuztOztprCf6nx6jm
md73w1RNU7955Vq09degq7D1cEU0IKALMovkU6tpSihJGaSfrqrYedqR/qLhvdOW
M5wXosrEG3DV0DHNz1DvyXfZa9YgC3ZyJzbaYdzH1lmHaL0GMi5364nXKpZTvez0
YtbUeAtWrXjHFJHCW3oaZwDUk3jZuGustvnpxJpKgYYxFBXH7FPFHXW6ziQ/oNOj
BgeqmQs/SEPMZT7T3rgGlO3KmvHTzxywTUqTgzzks/5CgXknpzdGwdJl6wMRqzZi
gPVzYtNOCPAvtA7BafJfJV3M2Xg0lqi8/FbMA+lgisn/coprDVn740QkNHUMRxJJ
6wzYniuHJIjOCpXZ4El+rcnwq8VubOp14ImScNcNWelLG41CTqXMxZ8ufr8mRnxD
ndmb8Ru7BO25Y+1ysHs+JDbZbPmFasCgkABiR5pVXsgz+6dC9kem0myGJI1tLyKc
7MV3DywrfCxHcr4zhYNE71jo5ruK+F1Yc4KXzIedEIAABiFj28rW08pgZwddJjuP
axXIq/PmOiV9fB9lXptVcK8ZGGAXyj8FAUSlYPd/dR6J1fPRjEW9iho78BRoxUKg
Kvh8gJ1r8SEgBQhaXyCYo/D3FufVJiFwcdjV2jijFIlFrcXDs2LA5dyuM9hHcC4y
5Lt+HPfCR235b1+rfxKVTpfUNQ9gphM6ZBgysjVIBLbmXYz71ZMA4otlwI9VaNY9
z1UbyL497OzMhVXfaXqwny9+VmAZCpDQPBifFJYXtB9IXelaT/zaXZhp2SQg3bju
SehzWcqdC5ykwC0Rh4v/Nj3adI+dgns2bHpAHKIapGR+CZRyLNTxiZEEJU6Cax4w
6Ph2TTajsOvhd1KiubdamQaXcLe6I8Id1hCfYDc75n2FdDRliGAGY0w7lQCK9DPs
5ZRladFf0z5ReSI97Ial2kZ/ZZEw4niP2o5nQijUuPGcbf+aaGOvIleZ9iNCe8w0
EEddbDu1JRawScM4Wfkak/O2AmYZuBkcuKvnZhA5I1UceqriajQiyVLRAC9oAiyR
dObn+XFHt0putdkdzssBXPfMSjWTobCsStojn3LM9w6rAuzs1HbQuYhMMUcGUgG8
43qo0Hb+KtWz1jFmSptMy7dFmhh9/ed3vz6O+b2oH6J4YwiKZeVbvneDwFDuRjI5
hNv37bSUnmR5+U6qzMcIIO3fxr7jS67yYnfhmz9/pCqIBf9/esiVkknaCHEcppJW
0RRZMwX0SnK6TVVKy4dyn/eSVTI+OEwznBK3w+Tovuc17TYU1/NSEajIYdQLgr4b
jgcpjD4bUUgTtPYRzAlLe+nPJ0mGK+TgmGIyT3oqBAQdnq7BbktwuH+44R3L7/vj
oxgnwVn2yPvxmpTjDHLT4hmvgd/jFaTxSaoIWmVmulhoYhGu1M5QJK/7TwcZVt2G
pTomeblGrB+I3lKWol/b92t6ZBHZBoN1SzsmtKTVb2jmXpoYunxQSP9y2IY27KW6
CHGY2vP3dRKRsbgOALEwN4c2l6IeyO3IMaJCHJu6x60nO4h4VvhkarIT71XnRyeJ
vDXTIL/7prBlvo2HD1taxm+vIMLoyKquAbQjw6rgDmTEPHgozixEkSQaGK1OK59e
Kfu+jnAT7FdaAVgMGd+ISw6hs/H31Qj1NF0tOD5UIo5IH2tTvw9YcjS5ZxNK9n6W
MgHpwrbSP74pD5fAiYAs48tJsa+fkbwYg/ijQQ6YDghNufDvRaaVwsnNfoBmBXk5
O602aah14GcbgV6rJ/O/+8mWdg3kwZb6MSmKUHpeCgAnadmj8MK2MF5GGC4n4Gt5
iU7/fujzdhe19rsFUsbMj746J18UqdPy0IVOP2Ywe7rSPBzlNamIZTlDrsbLMuv/
4yH2CH65KzwG4qC9pVR/dfzKDuUU3ihv91yB6gAvYAMq/wleKC7gvQRFib2CnxSH
hPahgtiBtN16ksDHgC9OdrnoeBKhy6F1c8PWrcQ64cMMtC/EJ0Rb9Wjm+uZkmLwJ
l6KJcnuP+AEHRf3zhsyrG3BzQiq6Y8rcGXBxgw8e6HOjR3+EhvS1AMTlefs5tcBU
3xw7NUoS7KAgYn25Fmmpa1b3zfCXtpvYExbiEZGg5/BnGTsAvZlhRCwLmczv7pEb
F4AK9a/Gf8R5WleWra1MupPxsKVuJcwXwjhwJhmzIBru1AKdBeptzSwFIfRHmOSn
i0ywm7W63qNWVuTscO3VWLSnkekn5OCPxp0mHfGMwL65sUMIZwJMSjhqqX6ZO0uR
rQVjVMmv5MokbQMVAep69wReIXm7+xzOX6ZTrLp/C+rSThwQ/wfqkLHlsWDju0Yc
bl/EsBH+zuX5cqzBuAoWOgrIdGwrrSPGT+7mSAN2ZTLUnk5GiAATR8Vhz/FFE59c
3mhbq6M7svGgUZPn4szuXz9oqGMzq0m+qZsUXWWj4XZcjnAq8113gfwo7gg1Djuc
43kWcOUWv+jbKXUWLy8x4MrDhgx5fgo4EoFRidCe9addsLYMvKJfUV7IJhUTwtAE
DqD732VfK7P7Juq7Vk0KSHIivdSGAjFGovSD0Ho7zdrklrmZWDN5UxiGRvPS8Qft
ESID1U7H/jsaIfgy0JnrwdX3NrlQjpUKOnax4tVe4pigNDF/6bq/yKgYu95+DJpC
Y43yLg2LqlXx7BIW0lUcTA5QH8cIij4OYGCU8KLHhg5GBx/EyCvUSYP6QaVMleBX
V0pK+C+KwY9yKHRkVemm2hqOS1hxUqzSKcPk1JzjWyyggPodEFWsibEUkfGUnamD
3ccf9T/QbnbUU8foV7fihOWpjEY+Od7U3He3Uja54Y24Wz6+SVjI+QjTmV8tIU21
thGJWpcT4naODvpl7xTJcbjVGnukmiXuLdWRHxZXClNlEZYng/2nGkr8urQYDH6+
Fu27dCkfNdJPX0r58GqoQ4T0H2i06YaE6SDjFqeZulWlrJE3plizOVuukwX4DpYT
xbO8J9jkKi/P6qHYnIGHMb64+W50dnvKVmv6Z/+iKWyWezVMfBnvgczft1UX/UsA
HL8mG4hRfglCRGs755WjPqKgGX1DdbaxWzQRtpKbhjCcDuPiXIYN8JxTVaeMktkP
fe+p6DHsXOoR4bGCcLnuRPYijo+qlxVQ/16yUT1RkS8c8C7RDGHmxk3+GYRYJm0g
E+f+SvMZ71R4Fi2M+ZbtMaQjI9LuRYt2ElSVXgWNOc05ayQ6jO/0d2YwPH4hwOPt
8jjh6Rdlducb+FOQngeXjVA93KVtCwD36LOsipymaMkGaCXOWlyqNb1BsLVHiMLD
gSH7oZtOhGBjAjSAHTxc9IVjO8bMB6XJYTAtDwoUT5lgXcfqqq5wIPCKx7RRkRVB
G8vvhhpBii3zMzyl2fa6P13CfQVsH9h57MEAFh5nIiP62lj3yrAVaVaNnYxXT6J/
68ggsVmDpSGa9Y9WmyRGbFOr+rX++SKY4p72kroCJOj84jYehyiVPYrxilWupL/H
k7ntde3Gc7psCa7E/htqCBwOo4I/+MXEsy4zLN4Yk/FL+AiPCzUE8QsRS76SPPkz
GKIiARSqHHvHwLxKf9PTW+XHnskYqo6Ae+3e/RjyKWatK4GJ3wM6ojoEQngtYcpt
orP389Ps2WR8cPNWiHB9x8CvuSI7XaV4EgK5en5s63vxyYJ203Z1fWj0ccYD6W1R
gMRKLx1w7QTJRYE95/cm8HH2lKhWbAsp2ara+Hun1/eaRijDj5aSyIcqh6vrvCYE
w8Gq60fWmSYqyHg3eNe98HoLmijqefUsjEILEOiFKISYWloQNiDgQMgKPAQa6aoD
Bu67dUSiw/NGN2hnH/kwf4TSkJZMJJ/bDVgkxnnyPwhJecI0vMV0Pcl+H5YIFCFR
TNl1eJHUpqfsnkTjhwqwVHUezMhVROHnQ+rhJqp9k/yeEDf+scc17ZczsjBq/d4j
j/XQwlhTX5rp4wqMrS5gUcCpuNh7xr+0x7ok9wkroFVDCQoefp4sqUUAry/WmlbB
X8iN+HOrI6GYHUAs2xDnRaKO6IZFUFEQWEt9ZTfNlPd1JIaWaaSspwJW59Qaf0Ia
nPWcYLh3MIgxrzn0qPPcXIwm12W3UeOh+co/ctZ1Zi3FK62U2rwa4mTTMDUvgu6B
R/bhevql1A1VbvRBoS3wh10Ov8iytHGV8RTnuWTN3F1WePL72Gv8qr8O2A6H+Jj+
PWlXEk54A0zeBg9+yGgElCZX0PReyT6W9NUWy8IDlXeOPKJQemGuaH+nNFXMppd2
rddD5oS/Gbb1CPlXaU7U0dzNlImIq+sxxh8V5ODtbijEGZVhaURHn4uWx1Bbhts7
AnchmNa2WkGz0eo/xyg4CRyDNMDb1yYGJiwp49cNVOqh3e4cXoo/kXnQcgdzUt2Z
jXOMvdE9967GDXUz5v2l7cdhD+54bO8P9i6Eqx/Mtkinlg/tTAr8brzhV/j8G85k
+8HXxf1vQkaQO/3082HoZS0C7pAvCZo+t0ZroIQ1z34liqvkni6VR0YoEqZ1F9Vv
4WS1pIwfMjI/7qPBXxKou4mtZgEAAT239e8br2pXgl74G6OSMtwITpCmxnpix4Qt
FlhUwZtCOUYcNm1MtIzlSas8Cw5ozxNhzUOCoao0deUzzp14iz+A9dgt5lZ/QQcr
Y4fveYFFAHknqxg1eMPheIPBb8VpTzxbEilVifYNs0ZtmVaFD9sGrOFqVegzDlP3
gbRHEVMr0Nq8Vi41/dJ4BXjBNCr2zFlNoGZAgW3/TKH18ZkDBuLWAsg0o5f8/gKn
+FyTPQqzhtMVA1WSrgkHX282aGNqLsbD2J2eThL1SKbhDd+FRg6UHX0BVjowD1Va
tI0G1rs4VWx9OimekcIfQ1c5ll23NRLR/JdTg0/xDjE71h2KVMyNMnYGAb3Ead3J
FM63wP7x+3Dqyky3nTbU/qHRT7RoTRoBfzYE9dblP4ilYCxlINW8osSNmXeN1M7Z
Qyi/u2O3hl77xD5qlUiW/GL6Tbz/nOD5y7dQMyc7prfw2mxd2CI4YoTt6cfXq8kk
uGnwFAnGno+1by96RXPfXXKuAOlXJJEhKNwgtS6AaPxMGXa/AzxVcEk4/Voa7JX4
EQ+F0/IS/xjeP0ip+NGf1pycrNn8pDofp4nhK385D4NI346m6cgCucmOg9P2jTxq
2YNVup+h162QsIPZtYaz+Lv7zcS1Ns/emMqQW2YNwsPQwxqAB/nSQAAki083+Mn7
2OhidB6WgfFI4ruBBcEhXjQ5ACFaiyzu4mcEfJPr2g13byQLORbhcAbVUIV3jymD
lYZMQRZSlqYiyVtAjSm1bFFzVBw1fedBl+G76YiaHdO88zJJSyVptd6Qy/0pL7r0
DTPsrzY42CqDOZ8jVH+N9iypY7ah+S6iNYGyBTWU109K1io3TYG6CJrk/jIGJ8wj
m8l6ZQDV9aY9d6xrSYZ6FcWRcxZRT1ghwDLKoJRyXcdnGfyobqiVMYl0ukKcu96/
R4xQOWYB4dVa/N5tSgaC1vaFLWhE66yGy8zSlAeBPMDmqGc+1UWgyHlBBS2oky35
Z9/qyHEIiGAUSAi5KlwZGrxoeAN0se6Orxb5hv1artck9lHvi0CFpocCpVBg27w2
P/d0//3yAmSKT420z2VeV43xY/S46Iw/dEC9Wd74HJLEwfkZEESWduAAe3B13W/R
cAhE92FqyxxSTqzJXDZt+Item5Qs+/x0fwVmA0s0b+8yrmpkf6U3lUys/4OdOwRD
Laqhd3XiRLLFuVEq9StYkrBqMrFxVxnq4psecodlXsvwK3k0G99VLrihQHsd7+v9
BH2ZCPRgZ1lATklssYr+hEO2F6c66rWwbBbmtWyMOhN5UIi9zAXd6qYXMTHL7DJd
rcqLd9Bg8miRcMtKART+geDLV3rKqIK8Q8HlT0HXhd/JsZSHNYLpVLtx5IaFVxpH
1H2fUvh0eMUW3uZLZZ1dtTPbLpQ5X0ZelUidPVtOkZlBGsuE9QFCG3GrXCrEJakV
mrR7CKZZvcLjubTVHARw4sY+oiBS1Vg5Oz3ocDcxUcu2p4+Tc+Y6dDVFeOtJwY0+
GxA2RXo28KAaPusv+9JUNSINzwQp+b6EpF59TUVhlM56O753hInpUB/K9jfcGv1j
hkTTdaxSSbUNhsjFt6qZNF89KVOZD4RrRQSZiHN3CwqzN65EZoLN0vYQFXub0Qot
4gVfVNEhoEnSe0EO9jMbSye6HuZinrXd4qYymCyIKIdCudC89T0KmlJvCdsNpEDH
jRCAtTOnA8epWzoo7QkgoyS1x83Kb4ycwSSoJKYB3dBx899SYJJLo5Flub0wwlwI
q8KlU1zCEle+1FvktBvpgEI4+Ao2Spp17yezpLe00bfaUmqU7etX6+Cbg1uFA0Eh
u3DIxemtcOw0CDTEVbyWoZ5JsF16qIOJVkkcFaX2HoWJ3a3dyL1zeH/ud50VISJ/
c5rOyVJyJDfNyRp+FgGr9tKiXmz29sm6fr6QHINxZJxn4kaUGz7BrknIrj2uWv1x
ENOkFNnGBdRRxbKGMXECYPjj4RgBnr0EJt6sB1tZWJERK3UySCmHztUYYJUqspDe
Qr1VHZqTOI3fQh1xhcRaV64fnbNZY7b58lT5QLYRew2J8Y0VBU+mfYsOiSd/IWZ+
4Xe2FkEtXY134mn8v1/NEbNYNKBDcVaXLtOXudC8FsQDuEFZG6fXFoHJ7eQk7cCQ
T/Wiq+Z6CrMlcVOqoWiykk57GriyfjNtbIylPt0fHbPmk/WecMGYpoM2JHEMasvy
ORuNAnfwxwjn0rBYJjpWHkKMaaOv8lBOLzg7fpk31BQ2fC7KnyYkq9v0Zfylqbb2
+YiVLeXFDEpbqzl3fktT9oXH8PwuLIcLRZhb8jrOyR3aNuRp6W2n2vNi53lbWUMO
4ijRb62iLHleL+QsoJTX01KbWmdbrNnvRXchiWCPzXmq93omfFS50jCj42xlBFpt
FH305to0TVKr38D6zDFkBO1OphDk8x1tGSGWcReyNJA63umzPICH1L1VUIh45lLV
jS4yHba3uFNaHH3wpM+REhFYC3+GU8a4rD7/wMzsTI5Lb1uLVa580i3ETTb+e6tO
/lZ/OSFS46xzk0XkkuW2LoIFq2hLAyjBgHArjZ9Spsoe9aEr4tI0mFVT3w4W4XVm
fUlfAGf1HzbXvLgldmsNU8c0uuDiBRKYt2g6MDG4GKglx/jkrm1sUsdI0UUjuVUR
DA2gl1PJtBZC+T1G9Eh+WxD3Z8gla4jC9kNZ0jjAhaZ931d/2iNe4eCwfQtzsfwx
I6gElr5ALuFAA4JlxWT5Lol3fg0aVCHSE888IXpCE/CFgyB3/DyVz6p9ycreFOzp
A/6b1OjJ95NFRUWynG4Zz6ZDDekNzpQXhqgrf9fBPVkDYrv8lVvAEB68qOaYZkav
oHQRanA+OeYJIsHMe5+C283pFGywXWLOosdTiWPWhinEiB218JWUlZaFJYpONxg+
IhG8GLC5ibwAufvm4JzvSIhVfQSN8t35erQgMmaLZdA0B4MvzhRlw9/sZTUAk8dC
UBOPqVwAaNpN0+cQUwbMe2kW8wvfSMh2K5GJt4m79TVbnOIlEnPExOdPKZ7IrPlz
R707cdECfM+fKuWjuBZ97/ri6s79hfuhXP+gn/9ci42eiuinEReu8AtSQyOkhhzF
oJNA0XIzUX3vUwE4tBtVhw/tLT6qZJYHTK9SoRBxvFK4xImpJ/I4UqLcbCz3ZB+h
10XTGYWdr8TmXPLWhU6HcKXLJjAc2ZIOxO48bqRsMx97yl1TZT49G3E9ktCQTF3q
zT1HrANW5dZ4bew2BWY/4jpC+13NxXvFbHHMCqcVmiw+Yb9reuTiYr/Rxtn0Bhsg
Y9zbQaa8fATjbK8x0CsKDRcA8heVYASfFE/guQ8zs8bw6cCZTMHpQWY1DALwqfwo
EZH0j2vUfr7zoH4reIWuwT6b1NRnMgnrXiZbHMWDAUHIBo9w5ZCa4ov8v69apC1y
5A8VJByk1z/1wg0I9SBokbC6lYA4IdmLKZa+mGlguXCPBkG7BiXr1ziYBzBJIWMz
qXjNHuLaA0nxDP2t86iW1s+DcnwWBCko48uCO12vdTlstUbYLVA4oHlcj2fnuGNE
OD6FTnzuwoA9KsUV9KhWBtsuniYzNllU7zxIt5i5i7ocxiJv7AQbDc8s979BA2vG
57ZUevGEjxoi0G+BVledAFE3vNp1ih4k+82vnSWlU3kly3QPS5CDle1fAqyLmesC
dkuTPW71X0AqlWSYlSJnhYxlewKVKeDAoN9izr46ZpnLsP9bupoTTFtnzqOlf6ze
KiymD7CrZxGlGPuKUPzwSHK77pfhFIU3N57D3c1MGHIdm1ANXZ+klC9QgsxNEsWj
XLKDZLQLRnFQ6cfcqb+bF9N+ee/iDWGc+O9cUCMVBD4mWvnYFq6bh2+PWcm2bUrY
kCxJE/foSoBKsMP+BgioxkdDCTk7OS439VKmf5+5b4vqAqBZ1mdfFZyFfz+frFjh
uaZum7wV+4mRR2xSlVWI/Splqv/YbT3Ru8bp3hbMVvZrtxHjuK9FIPwlL0QWiaiM
5nS9KF8vf46olMatdIADgM6HJV4auZFq1ahTDWepti/u1R//wS6Noa+AIDpCh7tf
yJXJ3xdm4e+d2oFVHLzJHEIObEu91NePfN6ThXMasXSqdqgZCzSXCZJVxJKR3VUA
02z3moILUE4GuB2/8STMkkCVGvApY0Eu4k4AjvURbZeGlTjDARRSqsENau53H8uT
HlTAv9h+g8XvxaGwdcVacwr8vuCume07FKAtxmvkUjKan+jE7GmUXA/Ck452YF45
TmPvmduA8vaVB/RwmHo0eOJZ+K4sXtiePoRMoBSc6w6dn4ycFArPouVhQsWA95NH
EsVGbtod4+klCIuCIcus9TklV1JZXF9pbOhp1cQSxlh3KvTSvqeoLO8CdR3/Lxuc
A2FZsX1oOGMfOIsfnHPezMwu9mSZp9sdveV7x9FpT5NzpW4AtBGyJeL5B2hFfYCV
Tl6oLcu3pJGrJaVShf7+kxJ4YPh7pVAWSUFv6Ac6j/qHPupCIiOhjhFKXk/+87+D
0fdIidVGymS1C5jfed+eBLywFTirBJtcjl1mp6Da2sk7T9UbFvBWVPP//M53IxcE
HMb2IDDgHa1bC6Heg8rcpDIv71DAk3p4z/Ngly9OQjn1LbtAqzLD/tuteSFtDMkg
j8IDD6ALnFbcLyFqZOoBJrflKP+oHxMwmVbd+x3/rJISwG0K1UKMr8BXE909nhoM
RogWFLMFB/VJTy+U2f0T1OGT0hKkaHLozRe1NyntDTkI5PzBL3vPJ88Ma9A13ejs
T4HjS25/VqY0xQvZ/9UsGgwSFyLDggtGLvJO05vC+QK/ZCpA7yzY53DQPsamMwKs
2cFOf7D051+NvZsXOTHVT1Nl6bN9cPk5D9NZp//5VJ0pkbEzl/ULScvpHcknT/te
grFZ3/iqp24uPQTGGS8Jh/ChPIVrH4tJoasL3bHAmq3i3F0NHVw757t/Rv+sDf8S
Ie6zM7E/7Am96vhbjIfLkVZxrPS9YMS3iWUSifRg4FmSlgim1/vqAH1BFLb4H3M/
HVMAa30/vA+wjgJgHvgzW9eIx8zwyXYDjzf23e+9dXISCbAmxyyqq3gp554fZ62A
WySs3NRiMWWoGU+JYXsl06zjZ7v1TQKyZklEzCFFmOh5PkJqUhG8u8HfI+Thy/f+
F2IXtA9NY8+Ac9OKfUp3KHKq85gpT/Z+15AJTT/ENQMXRXZP90aUuM9+gB8EroWb
bRL6cLsgv0Jw0+WahRC1rJq5DUAN018S7qV5f3LHQfK8gBiZdeNYV8xrTmb+D7st
nqTYW4bU+t8YgeT392ih3AZgyuSguFDFFAI4yzNXpzeDfKqZv6cXZ4nVy90M7+EF
N3Rw0RZucXiOcrSJrwfZwopd2HAJyFwx9LSs+i7dVRLfIqlyNbaADPVvZciVKxmx
cXgEgcc0GajYSNAn9Q5Wt4CAAcqeCywGJGvIqsNZ5Ff2IFj4Ak40vzbNR/6Stxlw
tc4COkQTyL+kt+fVhFIHjV4yej+HUKzsFSyzPDEisv9lJlnxwNtjru0SRUA6Pbry
rZFEmOgfhhbZqYGWJEq2TJLUOZSAsgIeNFDoVz3Sls1pJVkf+hoRYci4ZSSb7/aV
p7o4U6FXSbKXCWx06pTtA8VbXBVMpKAppgbCw6mLcIDjAoLogrKLj48K3Kt2CSIl
QQdtWvVu81slc+K6QvLRAzjmB9oGHMvoJ4Bk+kQkvFnVjUPU2HBlhKI1GTYU4pgU
EHM3D1NCYV4Q59HjYZFvoVr5yw0bIdLK0FfduthXuFJsEXCcJ9Vf2YGVcF5Y3Yo9
y3kpjagU6/N5nw6rsUy979R7Q5u61ZqHu96/VXMRKO33w3466X1QvA7lwHcLLLKF
gxCUQOnMi+MDMhigalbJ7/18pjWlw8eulVKnhab0fK+04W8AKc24Fezpf5y6ECkh
TMe9RPN6OwJKcgiDTzv09nkgX62uB4x1UGXgixa/JQjn1hbEgf8RJlr0ycHfCtnQ
S/yNh2UB8rl8vVmUVD8mUVRVgJ1RE7ZP4xRN4C3Jrufn/X2MTufoE3ppB55pCQED
jwIpCNqCe6ZZ64qjcRTfppGxiFTEc8BGju8YQxBu70/IXoEf9wJbLC9xgEVgVHBO
1HZHEHWZr1D4aJFyckdbSEQQFO4KzyB7auKO4idbcMJzsQM3kjLLoEqcEXnNQV5K
onSkmJE8y4qI/HdzayW9jFLw89cH/gP6G0IBjFDgeB8xrkBgAJb/VjZcQeLvW9ya
LZxwn6sQ+dcC7UpktnbA1vBQbHYjw0dgduARY5J+sfF6U6KSdlZy6pTsL62GOWJI
CBRtQIQ830nqzcxT3Dv5Rlb7sILiVSdbMw64XsRpZEHbNzbPXzfzeRFHfU+bpAMg
apRZD5BYuo9cXaN+r603S0YsFWNyQlzVR1FhtjLz/jgjwmyz6+MvE9LePHcnx36M
Uf1yrVDuGZO7m0W+UWKYewKo+sXDzoU4LLsUvXkdfcQ9/dfYw9sHqSIco5+Y5IoG
1VH2RdDeKppPeNxDFlIbhTCppM8K4ZQl4IXjFIk3qDuWzpSPmlepfpKhY6WUabcv
keMj/iIygnZd2F8zJbgLZkoFRZwFeWNZ5+RWJ3SsQMvc+cNxUgT+1BYBVwzHYbbm
BvBbc+Tla1kEU2AbSOxTKGoongBt0vdK07c/pBfD3ym9ySP8EKGZJZqf+0X0zOG3
DktEQ5BX5OJxgCr39+ZYIuPrB89bHKEhIYcaPvIVxzO6ytXBQNaR/QZLEJyHni+J
hIox2ZcVGyV1hhC9S9L7Nv7XQaOFV+LlHS2gcLHQH7vSS1AlM4vDbw+l+b0lTn9Q
vJhlxZlCyD5UX/5UMxL7eQuCzlR3DQd2V2ZOLTufxeOaaSX6jRIXW8d6EUKKcwm8
m0alj4WPUK/Hm7bnHMsu32/BjAt1sOS5z+yWIGcxwIadYqAO6FY2hfyhbwS9sVsL
ebZlx0oA60inqAO7Wx1tlWDr8S9cm4GjywlETCp2hhNpN7nVuCBU8J1cI695jCKT
Vhz3CI/VSjDxChTpIHxjxNvDYvObDd0+AD3ZK0sllIc6rvVnVeusMnOQgf//lNCZ
oMozz8c4o1agX3aZ3/FwVeGdebp63RhAo0ZVSqOfvRUXP3RTuwJID//4lOdz5A6R
gW1uxnxs0mr8hQ5ck7meaOHm9IH5qvYUkqILIhNYJtDSWWY+u17XEpQ1s7ltdzlo
T8tdSNNnthJNqHDkatLkZwnkH5xIOFmKyupny09hmDvSbTrFnY1d27emRf3vGC+d
vZhG6Jsyg8XmcztKls5jqA1cudqb8b+DynaqKLR+QmICPtr8r0ew9U6c4KJJddP3
OazomvLrqDTrmTyBSHnGBJEiES0kv9HtqRfYMhx2SYU8lUs+SA0VScn7PT3Slnda
OqMcsJB3B0oPJoRj1y6yrx2TW22XtKVmM6kz9TWPXbll97kjQP8DRaAOftOX/Yyz
lHmGxV5qg9Zek8FyW4QxSAWDXyYkM65m6zTg0enG2YvQl12BcZwn/C8injIO+s8N
RdZwOjCZabEjMSqb3LoilgEnLlmiseMMSGf7O+m3fYeGskrD1IVWJNlsafLB4YlS
hSxEMylZsu2347PYHLW64n+iEziP2yttR1mN7cHWAnL3gXKHHcDNsN6+YSaOXCnp
2mKLtR0gAR8jEPyQEb1gwOtoWNnT7d22HRm48oORXdHbEphhCQv5xc67uuj4k1Zk
wGIXJ4OWP+A+hHfpOFDEelgylq8gOpLFKSUnea0bIKTmlZAdd5UaIsc2QuYp9CqS
Jhj/hP682gXAf8AIOR5R7jM01kGt711AnmQQLkmsYNu1sElg7/68MhroNIcWKHzN
Xx1gpwXMkvihw2sNJcmZZbUCuPKe+Mu/ctvYBSPq5EW6be4lDV2M/pO4miAsetd1
B/iWs+RqPxaPgOjqF+hHo1nLz+O4hnB5Wx1SXqrp6oCabydZQUtYpZABs+42KTRP
xwbxSM6+AFgnKQC4tcm05XP3Wy46p+I6zK94+i+gFlKS5fWiy2UzIAOZFSf8hWaZ
eYlVfvrCMjkG3les7RPKmv/cYRT1fcVMVcBMXe9oJdfR7SJEUkd7/9AcVM2UxoXf
jXTDJxCB4wgI8J2FgwwxD7+ZCIgSXHxIYHNKNF6rauI7Y41efcTIgRu4CAjPay5P
BIqc6JBCw056WVN26EWHzVXXjgRH3gEBtp9ZcvI+CnYW/n4b2tsLF4e7eBk/f77W
mRdjaRk2oLxn29d1Ng55teuVQ6sVLDJagQG5bZjEia4j90S5rm+ufmERzOmQKR8n
kDUfW7yChAPgGbMAOUZgbGaZ9/MCLZMVZ3kA0k1r2y+wGIG2gZeKLTqAyYc+0kmi
cd41gKCJU4+aXwHlwSOhcbFSAj4Eo5Jee7Bg8gCbZ4B+3XIqnfV2M/v0UA3VfpWN
exYD2riz9+zcuK2CfBmxZf62nBZe2lhB49ENHQd5qMQDcAo+2W7OT9OtP9fhI1ME
Ct5rBlDnG1Hl3ujMQKXaU0xkpMp1cdkOV1G3miYL/TcIoVNUtpmd0cKWTINsu1/y
XBemud95nml86VnEFfb9wNwKPAOTow9/osTq11IyfOuvav6+XNedLdnRMPqF7SeB
Ljv98kygAzKbxg5EdC5YRGiMSiRtr83+2s+z0+YeGVNFiyFj72ZEu9bqdlC/SGo8
hBv8ZG27pzOh5ufYZK0ZJDkYbyVRU/9YTbPlEmJeHEBV08SBTEtQLJGKpbfuXikh
7xN5rMmUXzbUmov7CfisTmvMo+j8Q6eOFPBZH7SGvd+hSSNa5g3FGb+pB6/XUZyp
Lt0sqEd9icc6geScp4XfX7ALUVoiSy18x8AHBUgMlygvB1rE7J1I95cNR4FKE5sy
Lu02NOzaetwvstyd1xTbkAgnD8bjRIGfjEjXeEW/eXSWYnkDCidwH2RTn2sSsO9X
AXAfyI/w25xEQJ82xsHzipfHSH14/xPWR1llZMZsqufknVKYFsLdpY271N+xMW+/
yUTu1DzeT92eke1IFC4obI3RSFVInOSRN+WYzUc9EmmAlvwKi2rmZrqIMrivDk9V
6shH2RMo2hUL9+4zOXcZeTqRemAPukhop9LcE5ZIwkOS2nbHZw81DUa2POaGE6yQ
mFsbCUZEsY4eyVSDZGEZJu2FpAdasSvzB6qrqkN3KPLRmi+5MP783UmQJmlllc9b
c3bAlzxYMnlUtITM6StAp7hJnZAqAyAO3bGb8mSGTLgHDSswLb49N2/CIcZCEvvx
/GrJsREQ6aaZQZwCnrey9IC4PSHmTvPIvuv8w6ZHjegLyW+ezEdxe/FQyiifmA9s
miMj7zxsEJz29PqgWsUiJjyBEeooIVW5yAGF2UVOU8wLxTZITL+ZSBZ+2Xvv3eHU
+tyR2PttVzWITehTSNkYFjUDTAZjFTDoCXXzSVFnxHlLZG0HSJHzDfpBPmMJAJ4w
NYJXHorDq01Z5telK2u2W4V0Urz+2coVBXeGPclZjsdPbbXG09B5tkZx2Z0bGI37
bJQQxa5ghABKjXkAUZkam6a6DYEW+D5ldBzpxieka0wBNTHiME59OowJvOv0m6Ri
KrquSQZx0fnMtAckxuNijRYvZQz9AyAujEKTR/252Kk0kd3sAJKMZNI3vQfTJ6Xs
Xj0S2gDIEkL9HbMsjSrsV5e8v3F8lDuh9aHTYDdRYW8/3ltjyT+yJcFIdDwq6S/D
35QbURKf40vAvtU3ve0wYriLKn9cCW8UfyuPLdOzdiFfXROcaD++Cb5fUvu6slfD
QjUw27znRWkkETiCfCqVBbSUfFKp6LM0ONHJknj6oWo7wE7XRZHhNwTOHa5sqBYT
+ICZEQTdAt3nDJyK2x3l5Rox/j3dvOz+ppER0ldt4p88+lu1JSBGMkfN5ppBPh3d
umiXioMW4d28k40s6Rlq5umvdehqLhN0PUjboFuosPBqMaFwngypuUoBvMLWXbNY
bDAYv4ylyCQk3Bc9bNxhisZl0PsBBbxpDxirOVSoM3LsgCDqYLuHet2VTOPNLzkD
grALnxkOk0XzZjpI/QgaLDCn0YgkScDf6j/GIhs331n97D1JskdCyOlgQmP5wfqt
qEa0MzlXU605RJqvY1LmKc3QxvawMQ1vQYQJs5Ftlbwy62D4qilnhne92Ey0lrlP
UcGrIY49YFIe2jrBb1AHIL3cjCTjknuPMbfC4ELXq248LmxxwmrHUE+UDYJ+4pyY
EDRxSWSmTsy42uK4DRZJChDV2ttmdRvNhZS/0ZCRzr4D2mQavZqEm8oYVOfHg9ru
DHuPdOQmckmTUTQHPMkqemPr7m35/o0IGmA2bg1J7oY1mEJO1ok7vx9JgxKtTVMY
Eh9cMFPfzJs3SM1GDN06RCf6wU2g5xNTuUHM6CjKtd3m1jrr1o9IC4bVq+t0Dur0
uNZ5C90tv6pucN547zfSJeraTFZy6Y9DBhKdLLdWZ8CnZlWbFU+vr0erPbAE6sbX
Z2vCAApesusA2WOtWlxdrmCdQP+Pw2zvdbgKHtAmXQFiq2GNt7ucKpY+R4qNSX+/
/p/1uoAhxEWNKfj3U9Kskpalqzba6KTqVDT0lQyqFdP2jfvuA/59DL7YMYbz3icv
JcbnuNspyFDIpoJ7YYrLL0B7Uh98QN61iyZ6pwqPno+vsp9KmjI0j9//yRRHVnpK
Md9+DaUdj2QLamFOY2NnU1uUGsSu1y0GuPl8F1cDWAV6rRX8L/IXfgtuhpQ6xAjS
lfh6rFebGIDG+UeamyFJgg9JkySqoeG6ckxvCAcNng9aBsAlJi2PROI4e04SjHWu
ZSjeviiCvMm6cajVUW9fywak08gNEBh2D4iOASB2yJXo1aV/SDKk8cxlef89fQyG
WRLu0dwDk9o3qgLPlLm9ME55pBL1pCIu2ARFd4T7Jw4tOy4sPregeSS+aKIosXXZ
bOyGqsqaih+8RpHAxYSxz52dTn73uacWB2w5EIMtldhnt2QhZ0gAH04tnKQF6Hqb
4rLNYqiRfRSr53qnmIxYb1YF9C6OSUtCFQ4nZlYQ/pg1gad6Fl5Ajn1yqskr1gF+
I4BusbffkmK7OZjNs7bf93tv/aQgJpgnrE7jthEErK8u991udC5DW3pRakDgY/Jj
AXcMtMWROB+ooTNGERAJNb/cG6OFrB8S72R03UNl3Z+QpRNpRpGsGVuHDM0wzYMR
DfZKbN4+Env9YBUdeHXfrBEZYs40pnk9tftEV3gs6LaZ0imE5Bc4LEjZLFSLugfc
yAEfFzNhU3uqpDvu+9B/UOu0AODCuHFaRjv2Du39wQtUTQFNAMBK9eHdKmefAs6G
6Vwpv3YBW0C8cIbcfCYM3g9/aVcgUNq7SrlQqEbbXzCYcrR9WcRY1PT++fIEOmwo
GcbBJ2Y7MycS36MogBMgiLTMxWDWDWBUGmG6mc9SwxoQy4P1yfntIWWIWt7e4yuT
QcHtBmcMQwam/we/MhKHLEbTsKfgB1CaLN2dh4jP2ZnWDG07+iwCFoAlRLvK7ARB
ZQNSRjnYVSKMw764wABl8s16OZOFOC3Iv5Tk9Z4uQU6tfDJ9Ftu1SaHEBQLbVzUh
QMC0rLJK9OCv6gghqmBLl8p0U1zb0hPBiT54Fha7IDO7FT8Yh9LiJbWj0E/VXYY3
4SLXeljXhPeUc++ddGdNSD+Nz0yVe7GB3vbjrSgcwwVfo+G35rWe4Qf+2PUyt0Jb
Mmrr0dUf40z2lZF5pP3t0TDdGK3aA53v9Sq1jmn2FQfjLA5mEqDPkhYDt0im4mC/
ykTDfrEvtWhNV9dCbtg5uTVIj6LvjaxsN49lk49Qgl0JWV4D1fuaF+j+OoFwv6EY
2DqaMToXkOGtVWsRWeyoExlgkcs6eCIezr8GlhL5DQfW+KCCyfpNdAagoRD71d3o
bVEULq0EHycS3Y1bS/zG8TtQKM8JWakTUrL8NRPBGYvb9z5ohsc2udMJW09gpXVf
BZ8rfAsmlOXL/fZiSwZu0i3lUl6lmYaw8TdNpOAIkspXHgiUUkFWDQ45GgyP8Xk1
hTgdoroM81H4Nj2PZUJdLfBMhtiI757QukqiE0s+3yFJ4Skg7EPOu0BxbGYQIj0b
2k5jn+ElBv2oC22o46Fkz6XHnlkqkFaVHHuSdKyjAzUddjSfet7bcUusnH0MfMlH
EdMAV7JDNs2QcDAo3Scq8NG+BiqOj/9xv7EKNLxIqQKeWRGMiBRUiw8zxvSINMdc
nQ2skbi8KotBLRXhnHhpk8W7gP4AFdPpvjPRy1s0tiJ9B3l2aRFlnHLd6t8mz1gP
rU4Ntpzkqp3pP1bNvQrgajtc/iQ5usiGNvcp6Nj/5YwmOt5QrrXKBNldW77qAcmc
fg4NP8vtrFgvDHnwKEUODFBwzXacbrfl7RIhluvUgYtwJROLygP3MI3qWLWVfbPt
`pragma protect end_protected
