// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lDQQJe0G1ngw5jYF1PlXe8wrrP5lFu1yWueR2q3InP8soR6Qzo+g3P/DuiNvYDoJ
7qLVB3hdEX/SV0vqXPfl3x67gRwhaSjS4PL1SHq6+I5pc907Bje8hN2aCe9fxksA
sw732KFGWs/nBgvBT7RBzWmqz7wtWc/G+lO0ifBWOfo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5504)
73JJGrgItSYfG1Ny9GZufesBrAVm8Zw5XsT58MPCXF33i9lZenBhnWhlei669mae
s+8mo2OKXYFCjTj5Y1HN3SgA+UKuL0W8gOUbTRe4du649h6kxrwzxm32CWPt5h4u
xP/35P/fVbLQxtW9TF5BjX2hHWgM/aK+wMruFh1T8XKwVvL28x5nv3BW44fgh99o
TRXZGvjlmrWEx24K9avFiLw6HY4b/3Y6mq0zhsRLyZtwh2Tg5DFy3CWfjtUTXBQH
YVJOi8XHG5R++c8ZG+U8aZ4utYvl9zUJQBONz7E7IBluO9o4VVG2fo7XJxkujlsn
ldQd9+Q30ITArkb0mk6rnARmE35umdh/00/7qiBlYJ1JV+bSTi4GmRbcKABjHzgp
9hqtXDVXO5RNYaWGC1w5gzjAQeVgkOtaDWjvdjLmf7yO9OeDI0PCmiLgjsRGX1cN
4jP0xk71TRVBjjbKsHjjieo70P+bpcUu+FahbUH9mzjGBhKIiNdTeRzF6uyN0owB
X5lEg3epvByPnXwlA89NFYJmZaEE1BZCAzrmQG5K2ofPvEqz3ZO8W/7brtaZzEKx
Nddn1RC3tpn3Oq/b7AyiKWraBJylWWwI4C2ceU9AyIBCQ6MTvDG3L2gX7yypj4KD
Xya95iJoBJujobrl0p3mrzcXaP7rB9MBnlF3aezDuAitYulA6qDxgLUHcs37gr+b
sjEHuoFuo3T459klSiICEB0negQfqUTbCy5pNyAIteOnYancMh5fd02RcL7SlGhO
Vt3KCFz3GXzHBJebGoxlt9ZetwBdHfox1Q1nezzMXbIiajTkgUqjnvogrJSvkE0J
fdPFHi1J61oeCa8NRaJ/F8kjxiAycr5awRuGsKksSD+p4e+f7OTtNBBd0CIdKmRe
wh3yqYq69CgWZiWVcFcdF+MgJoup2GsgwH2fB3S9pqJRctuQu119zH4Y+qsE+ER/
OjIJZIULuFdCOWaBiVRICf1yx5xShmzCr/7Vehbl2DgDssb2Tau5ZAaodG8lbamD
DTIOS3vzTImUHgGO3IGZbPR/I+RYKACb/ysNBLljg7XoouX3xnVWI4348Qe566zv
+cRD9jvOaurK0ujrcwIljitKPTEFCBLwJuDCg5o5+xlt2ymWzmBKz2xoBP27VzqV
myPkiWVZYx8jKCD0u4vuDe4iCuO/4FegxK5f/UyUowm/X0OgSgztJhPmjIEatP5d
5R7EaEcsqCjgLFQ+2/tp3DCFFam7HqlBiinoUjXSyAk2cWNaxLdHX5Z2eZzDS2GZ
Pu43QvQfySikoHkDZLpTcE6m+6aii5228Oqo2aoP26ZCk7TNWdSkMHRz2RGycIac
ZDCf7NLdGgG9yu3UiTOHB98KHepaftPc2uosICULUOrzgxEYoi9Ky+wkZghxrRnO
0aktD1TV7dHO2j6xzrPsqgpwSgmdatSQ20d6CS7X41E3EXKdgh+bo4Q4fTpvkld5
sADsLgf9dlxR+O7aezu6lXFKyM8tJ3DPUHkM+3kzsE00MGK/7cZetKm6qDWdi3ma
hRt5zdZolzs7V9kD0Ii2I5C4Zc+ub3mct4qgERTyBzcUxWVa0WNPOVZHkzMG/LFA
WWwrqVsediCL8KTFc1dSAFX0n8vuj4Ldf/mlSZnvys6+4Uer4tL50WJEW+hg5vlD
Mni4RpE0cHKZqngl7kY0qHCMGqAt3i7k5h3Cf4tiyWALXK7sohxUkV95DUllDFhP
ChUpcN2c99kkbjEBRxUqsE5XsJTaEosFRcBILS9u7KUndZb4KKTr+dcz22I2gBAI
OMIRjtKLJzlJc+Ke/xVhW/uvggYMEsisivv6wRob/cUrwOkM0B8JkB7Uem5foLqR
nkJibZooMuigFa4aWQAz9oq/82ESuj5iPDcD40L2nRoGGQSzwK1iN9247LdDEp5K
AEzY1LtdgwS4dxiDFc/4D1/iUFmjiN2JlX44Hf9n/h4uLqj31pD7cFjq+NmpjM6D
AOUk9quMFRuSPZoq3LPC3N/AZSg04h+i23zeiEaIPniFHznIDe8cFro1z56EJMtT
oteEBZIUn3TYEz2jur50bH3NNLR62R0plqt8EWysmdVYygbhPcfe6/uN26KyiJUm
1+CY6y2XrJlADK7PH0DRvIt0KccqIgqBE9C0ssehkYDa3nuWAL13gkeGHLA1kvud
sLfdxdBHyCHFyY+h0cHkBF/86fe/2+fR380PHuKddpGnhdjdo/BNimfDoZMd+F7e
8JSSm/X4Ura26723AcrzpShl5mVegdB9oRK3GGNfbf6C7vQk5ruxw2QHKNJMfOfx
Y4nhD/y/Xq6Z2dn0pY0LQKl2eC5SIvBo46w9B5rDpS1ElW67xSzHFY6N2NjHSdcw
AVRuF1U9RjSmX7KPEX7ZrKzCQMuHGfKPsalRE7xvdhRmNJplsmk0uCGSukxQH2f0
VC/B5CsUhy7cRrU8G4nN+HK+4PCzXbL+VA3Ow+aEjL7mGoTtq7anLrWDfjn9REhW
dAneJHufUQ2RJqbpJspR6kWn2uZhddscJ0EV6GUvn6UYpaRFOHKp4Mt+l8WMprzK
iu2pUj7QvPTde7/lp9qAQoxM5YgIV/8eOLhKN0uyptQgtyktu25DM2FlVvw5ZJSQ
GiMnHpRTBLtvM64KiVj84OmYDhiwCzF4Nfr58C8XcrFy1UIsDY/6bpySb6+5Ky72
qOfAw5i6KnprSRWY0G4t17QhXcFO/VTQsoel1BsmMv8ilbOrvbtdPLzA3sEGvgg9
2pC3leWAix4TJ0nqWCmYTYwHNWmwwNm2bp92iw5ixXxygEZXb2/5vm010iEI27kk
7gqEDvuTeHhVOwL07T3v5weMXH/mAWRt1vY5RT+4hKVGgwz9nMDAxLq0AqZuKVUs
Eb+h/UmisqV9LCeGkAmF6sLY9qYBCQ9h14zb93cOAdwOhvpuyzZnlQPjLVAtBLsZ
IxRg0VPLYg60/yd4eZIdhURsXWlip9ZAGU51OcC/1/PjPXvN4x82ZDIkVoSYUc0g
bdxb6ZmkJIIUWLbz3cSw+s6ZKV/vVBkKSVdmoti702dOoVj6O6XsZkJrLepbjNjz
Yp/mVL3PTzeFLVMzmlOtbK4ciPgakSCePHRG5uOMcjNTeucH8yNhLC5F7Rh32bbE
kdC6Oor2f+3FCv5K0CRDa6rDZdBJicTtffUXz2BQXRDLZrDsnLsYoZLmR5w/Xe40
NgLABd8R8brQk51qYKZ5MJgr6+EQLQSS3WP43JoSY3p6UpyyYHKKmWq252ZFzePE
FgtqkRvAU71leleWSXrcbAO7sw0ls9X2YPkx96CWaZutoLq9vs1ATh7nSl3UoA+8
X1JG0z4kBIRZLm9PSjAbIvkr4/+tOSjSCEHBbT5FTk4pCSENAepQLju8z7C/wJi+
4sDLvOfrgnlK0TJuCEH6/7EpSovf9UoPEs3jHo0o4XDIUE/OvmK50BR3JYhVV0dh
pg1AUXI+z/CUyHXE6xidgzbajeM5UXz4BXQks+kgaThix3p3g2Iz/zsqRmB+rrzw
4auN4ulSxHPvNwqTHvz8sqCVLUbPKzq7/2P9mIqnfr04RZQha7SIDkMchimDQeAy
hn9159MOMXcRvzPPuAlnDo+qkJe4XCJByf62iXQXux8HX6LpZgltEdmyaZIzzzeR
fqsQnEymyWhmUPP4027bCffFC6prBMkTGUjR5spL6qOb5gKpCoZj5r3M7vM1o+2x
szKE5vHNHxYSO5RyneX7WPPkYAFinQ/6lxT18msFOH+v663GtE2AdEofWClYH2KL
L4GUmdiJjKpuvpwDtRt7NSvip+1HPty7EJM7NxJbzs61UeNp0M+brDVNFHLVtBHB
kUbO6oqdBLpF8wn+iXp6bXdNJHN1gjCkQuz/O9SFMkom17saq1UXu7vkOkwpxpXo
s1YOdm5nx7vBMZjhDJdcvybdIKvdzEOQS8UPIQMInhjUNo4ixoeYy1+TIvmW2I04
GDXV116peeO2j/rKXmIzgyQva+D22XgKM3pm656MyA5TrwEww5CAnjB8nKtsV2+p
vfEilfKtrJCt1cvToSgM6w6fKKM6SL63Jv/sy91PgOYPylJvHgdHjd8uZFss9H/c
PGJchXKOyzEBF31A2bCtaUyVFsnrFGCUJ2pxkVtFV6AVs+IeXFsmsdrAPjrAIhbA
Gh+8OPNdU8Sd2Y6VrkWofBOm3xGoscTBDhOKLAViRFhfc+eaWj5TQbNCN5lRctkK
t17xriBqvSvD4zIwm80aU+e2tumIP/w8YnJpMUjWcfPV4RuPVBsoEa25ZrJPY+kO
zKp5UlZphFEmXU0JzYtr+hfoXzq0qpgpnhbeWAxWSq/Gc/NNVzfKIhLH8jLaS5VM
0xUmRAvJYK/VZw3otTUR5JxDJG1NUeFUWntUJCPz5uOKufSkGy/JCdIHfgOyg9l5
VGm4MD40hCOZaaIgxdRy9iDlEJpl7jMy5HEakLuAmjWVCBcUKQFTAsb1CpFElVB1
7U0ikWIT2Kft5rlwdLhWsabfr2F+cyzuYumA6CA+7lUN9O++V3Jr/pOFHaftvVZK
0ArScQ6D1iS/VH9tWDJ3K/HW7eLnNqTPXlCCCK9UTSobvkF2D8QKRfo7L0qOeOOy
e9V3mVj6pMXqF9CpxiPTjTweX+9fUMZt5xLnr3jf6Gxe7J7+goJTDhgy4U8a+WNk
1A6Xd92bP+Hg4rFWEa8F98Ahoo/orhe0h5TPlVEea9j5DOb2u5ekHEayaQ1b3Tpw
ft0Mc/gjnNr5ZMrYlCtiao3ncLHDTmXA0B2UL2VOU9XyZPHM5bpJxuBtD3YHlX44
CRg2TtohV5aTaCA4fCrVFmMRqM2Tme311PTfUoV/XQp5OnbwINLUlQxCEyIUBZCw
/1V8xNbGY3GT6NtIR2OJ34R6CLbUvS3CcEfU0qFN4NLALPo6oXsRToD++c0keZsP
FD4u6FMgmMR9inusYzbR1eC/KrazKtUA6blWFbyjNi3s5UE98LrpmYLporvaOOZd
ktAeKjk4kEdINUQx8KpyJ3DYahwo8FQxlCh5Ni7rY8UR4+YoHCBsk+872JCbzy1y
azhTsikYef+hu1Tba6+M6uzEUtJSFD4iwoujmXg3ctdf9aOuOHN0ChmH46891Rb+
yqldCgnjksMkxgxWIa661IkWPEDOpVjkfVlNkD/ZugOA8qVEGpYdGOAYZQWMo0Ty
PV+bMDW2Iz/UH0PhslptLGBPVKUmAJ+n4WT6KQm1+xKruxd5E1mXe70gMQGZYUhY
tMdBA2RgalO52RWRoYJiA/NZ5xnlGFmSiPbDYtR/+QiJie36eCcmIxp03BlLBD6a
dpwWuumqxpqlAyj9Ba1KrxRa+//tBYfj9EHJWQPkKsGqn44W4uqqpa1aIfgGL4DW
0q4CZD0R8eVow74ht0GCfEp1vwg4PEzG8tSRWI3hGHm8KSc/TsaJlWOx5lWftPb/
dG7mwHo5B5faRS6WEFwDOZdEu9A8lRZzKiWE9klmnCdxexeoLT57Ab27eLPCe6Rz
JNJ596GMph+gBY1/XzlPYqVx2VCiIns9Vl1MrM8D8qERxJLwNzjPdxC/dViW6Kys
4h1VbiuCXVR2PciaOvN9fqMiH7jqJ7SawCZnN0+pbZqrAgcZQ9xKkyxYouRk/ygJ
b577vEu1nF6C3IdbfMjsnl1KskCBIJe8vtZLX6BrDUZS1pszZpQWSpjL0wFnNB3y
Or+cJuG27O4PFGPD3wthvGYVmFUh/fLjZYZ2MYJv6VVbJ3gNmzUfjMsBuXX4vK89
N5YU+qW4R68QQGHQpmF5R8chj5tp0SrfyruRWTMoIqv+EvjCv3WhsHTGq3EdFmdE
lDhD7df/6Wyeum9uqjgccTQ6XfVWmsTD5vNinyNG1d3dp1zttF2n69flrlT13X58
e8VPd0Q5Lxh5ixN1uJD1fjHTeY1e4gvrM64wZZhLYDcRtkD/nHwQXKJtg9fPTJk6
Q+gy9623wfVc1evctVCVC4q2wTXPPVedGfESxNKw8UuSMV0qxW5EmUPFZJwemKQL
bhegi8Ht9Y2R004bCot0G528d3evrCIGGn4nfHk63fjPmNzWinlJ4MHkMv2PIUnz
mxfOYGG+ITj03vr/b5ElQ7OHqjDBxOIZcRYyrIFOp9A2SGBjLDSMfZo9zsoB8YUD
U6PY2Md+YIBUsyZXpHzOPxdFDlHbT4eu4IsFTH6g7WRXwM82jk1iXC2t6vsoCfh+
JZoF1FLhmoPsWCNru3/yiX/eKv/166aMeIVxiq+S7++HA060E5sNJX0jrB9ONvwy
nQn/Mpd/qOM68v7IYXheHz+Qh9hCZlaIWO6VZkLC1EiEN4S6doJ0ngJG6QJ+gCbI
gql59NRKV+dnU/u41i9Nv2EXYR/BQeqwn0kkVsVnpMtyP2X+EuvD2fIfKmfoka0F
sbBm0mJKvEaRWx44Bs0CVBuggwfpGMBq5yyMKu4QXA2B0/faHI1O1BOhP7u+Cbb4
AYC4KZtVCO7n+F6aUf/7ynew7GBn6ambxeaCcixJFOfNHJO6XgiHnPWEhXwk2D8y
GgAzNPm4Fixy0mDjFVs5//tjfoHFZ05PQLNrVbw/TFIw4C+i/ygvoli7mylT0did
YUGBVOFuXYamjukPrdItTfnyEq3jOg50rxqBH+QLsau4UzVWS3wnFiPLMR0xBPjL
+zqKDJhDPr8xI7WWToz/yFaYnfUnijr2QSmDtQYM4eZKMFzvnGtan6/H4+qx3TC9
py8u3gvr9tYJK2DI2lG3M0j27e9qLY4sz8TlS73idAzVgPnPS2+ulzNa4eG6BYTc
JgJyH/18/ksRbXvW3YYpnThN4Q+25AHpZc5gILmx1B+U01h1UUBMiowioj/xEzQ/
Z/pT7pYQvNGd4sRobMKWIB+ptZy4AZLUskrvcb2C9OEPEFh8HLjb7ydftgP8Dksv
34F6NxOQ1xnh5dbs0M2OL02xuQ79SbuvS2Lw1CHR+Ebh+g8J/fKsh/R30K75zjQt
cpueg5YSF4J7F71USoF5DDUmZi2ynfhkS0SqJAbMCzuubFjuHmICtu2u/ypnx+4Q
WFwbvJBqIez3D4OFf8w1Kfp4AeEwnQTsbpP6VrwTK6UeDiT/y8Rf1bGDLYwvqDNl
GdeVJeJcUn2YgpIFGtjROnuJ5u7xLigpoSQ3zZCRMTMA3awQprVGTUWBpOlWl7rU
/2sa3mst6e1pLxJtx/xiaJxBZPpmvkUMDbUgRQko9VaiePguSDf0A0jeEdx0R4mQ
WfGEubqtGhjYlnSH1nP2bDdXMhpqeRP2QNr8xMmkdaX1alMfxX3th6lSX36Ej9OU
f3857CF3bOBCILQq/Lqt6MW3xPQOIm5MfXJpUlNRscw=
`pragma protect end_protected
