// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nf5s2y2wdnyVrOzL63i1EmW5sQwUBvi8upLB4S+kR3jbVQZewZsYQOSSOYqmhMHm
5L93/lDxupJFRWIdKi6nqpo5ruEwv0DxQxDSU8A8kE5zcVDyY7Vyljd3AEefP7cq
QzIWIGfg/7i2bjEOUsGQdMues3nCG4dICQHgTWRPJ24=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2176)
zNcJXoB2Ux/LkqemnUu3mH+S20sgs5J8aHMbEonse02mtO7TEFTrkF8CWZ0MSwDO
LGxelOViDlNQIkaVW2H+rY7AjcMFP0C4+O+gifbuHKSjgepIoaaaLFh5s92S2WLg
tPGxEaxKY/EDO6ll9xn6vfLVOGpyWJzMDfT9rPmzp45i3KjFf8gZPcUQXSIRHIY+
rGyIAfQaiFP4Xb7zhJs6CzWKQdVgBXTsXzSBBnOeRGUbFyAE8VMENNqnr0PSkdGa
k9PRkSQJysH33ZNo5dBFRDtlyRS8C2NHslh/HNZNMTU06wsrFzyLVXIbP+zDTSBz
ChxFFsl6barAv2nG+q3KvzfTNNnT3dwnmxJ9Xebb30j4kHlHp+E4hlxDKr4WqOo2
HK34xtj5UFMM3COTRTI7UtX4AG5Fu+7XktvGdx8iugpjQCCT2jHWt+MyRUJETU9U
HOgn0JYmBOOuWrQeZVdGaQvDIWfdzjMxWFBHIZMLI5RJaGXdXyuc5E2sUcOykwbB
k2Lx/SVgbtEZBEiBWxDURGF8FAOtRfdAfCJkXQTlKjqz9KJPvoAgACdFcYForQW2
1oUGb3MEStZ60t0W8BmSMAIoz5qZyEgx61WB3lzWIQonmDEOD4xyfaCvdg+f8Y/Z
KMTxYxBlBX9SqLvtDBsA73FaDUoNg7sF7J/gPJgNan4Lqp/uLFCo4aKK2lsZ10gw
cAihCBBVFm/fIsn2fpZsY+si1KeI6y7531o2C9ZD3vKveTSt3ZxAfp5YejulJ6tH
kvETdK0fHFav3t0n8FQ5CDp5jIkd99Ihf3c0G49t5pdvVpiSnufdWqW3xR38Jl7I
/LWrt217Za+oMr6V9FEKaG//CLbZqCn8Oe4dzsuKL/yzrpweF7+aiHfwg090n/FP
M20FiFuQFRPFb6AaYOaQ/6B+RvqY40EcFwU/dXQAI+ktrhA7BYUHo9QhJttiXXSe
cRU1RVqrf1Mr9UMmaZDa0EckR6gKiKFQZORU8VSfJudWC5WBzYVA1qK+eOMmqDw3
o2ApgeLMBbPXUMKqPUG96MU7O4ObqMmEDxI8+R8LAYG73AeYIMY28Y0kBtGyRXeV
hyeYfCt8DBUp19uRjpDsidNUFAUwuq+G8E/Bok/7RpxOS81q25zwsWnfumPNi0vF
UnYhjjtcmw51sR+RsDgWaV95jzkZBLbrr8tZR7xxcOyYg/z5OBanF2SoNObcfgsr
iUUsmxGLOyjza3ITQ/Hf3lpkxunTn/yPYH2+yln7VTbl2e3q3PZ7XXq1kyzg5zrU
gue0eienTgQzx2kA69Z7IR5n3WsRThE0Acr53cLscFCqTnWpab5LO2Wah9CwbwDF
HnedVhaT2KclL29YqRi5PtxoXntwVPiiYqANZC3SlbP+MnZzAfXBletbhmtzIJhu
uknFWjl/mzzAf0pMR0b81fJxSsYd8eI3qXF3/rtjjlZ2RM1m1cU9e7Fmd36orvU9
0rLJwYLYdr3xsJSbLb1PEcFh63W2jHYDZlZp29epNkNNPO8xq+lNsdJ77CpRHWOj
kIIISV+7Gpr8zTrHXACw8U2iL1oryk1efYl7AueRrs6RG4AMUOMEybojBbTk0TT9
Y9bX7+XO+7HQvyJht0hTGmIZdey4Av4VsqmZ01zVsI0PIbMXaHPF9uG+LZuXgYFX
3gY+U5VpyPU0+nQ8G4sIDOF9IR7OZCGgWJGlEXFhCU9ncsK/r6JhSfAd0JsdbqcI
O+FKrx+7SSlhDq8SxRFx7biFmDOIFSXrD4m9NTUHFUxflNTCOc2YpRrpuE0Zwu6S
WztxfqvvFK9jMtJ0ddCU8dhsUED/rp9rFTG8SMSb1l2vcUCioPH0xb1Kv+cHZAxY
en2Hn3Q23kCREgZofDOiIEAKIbekPnQ2r651IvLPkCybu2TnNKgtwAQ/Lmj6Q4D2
yUl23DhNDi8x+t06S7kVOL7UXDAO5MZaSSpVLVPnbfZD9HEhKI6Esj7XuMb+kLQl
/UCnV6BIuPxdE4ghR9aLtVJbkQMzPInVGH1zHPHnQHlFGeE6yCBrGQ6aPyveSHVj
mMPuuusNbZvuwy33k4H70GlUdVBMsOlUEeCcd1Gp+BaDHht6bKovDFULIW/I/Gjz
rRcCnwr8M21qJOeyT0BRTiNzvjsapv/hz+PIbfUuGIkEK4dbCr5ZtB3nUOndObrm
HPAKJJYuf2/rS07xwQgogTF7tqAL3sb3CHO5QwLxIAT9GrULWgMTPb1kWmgI3UmA
n6Q/Qt0hbzgx21vkY37nAsxMF4Ygf+5+5VCS6YRKPMvNpkFHCR8khOvFVjTNLnpy
fPbAUNcNz6Le0PGDMbLr08kboOK1MlMl1vssQw/Q1PkuIEHLNentbx4kCM83/6Ns
glfsZrK/IaPyHArDOALKxl+e1uDleu7jlkQvDAANxVChYUZ/4o8JCC2Zpli6dZlx
mInySYfpNX9yzmQsnAyY/skOe9qVb1qBATMxPvf0CJY1k5QRO3ZhEOv20fgDxnCM
mL5mfanUT1BoGRugbP47jsKo0OT+Y6uUmyEBGM+mEdkC03zHe3/4wyS+4jOqCpDK
Oehdp+IfmKO9QCDtTvNh4TQENfHHAkipi9/kLU4zZNiZHazDnJa46fSEn79PYDEw
mQ8GYeOF8FCYUUMfwxOIMhcUbN4gW9yHhsn3Z1dvkYry0hQGSS4hdi6PWIKFvavJ
7vgb0F4NmWLsTR3oaOKwTeHX8fQDo8IGKgBzzRW77Iq/wfJs6byoG68fkhcg3Qmf
zEWZGta5ZhA+cUT58C28hA2oe4r+3Wl9yjSEPmgVnQ8c1/Xq8eM0Sq/PpcYwZRg9
3E5ITFKCnfyooOEcW22/M2kHEZyr8L9sOHzlWyUMBy7+t8IFUPlaU9sXOgmQNcgG
BnnMru5oMmC/HEn5Or1cYA==
`pragma protect end_protected
