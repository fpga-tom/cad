// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mXN33SAXckA7G3ck00LiW95hZfpm7Sa5bj3ciJedrUJ6c42QOVKBoDkiN4nE4o6m
3IwmHweH2riELgl8NNSeUZQHgK5QMTA4vhWrSwM91iYUOFyARrXC6nKYBVdG5sox
Qs5oZ1kZS65gUx7N7D5/WEnnRsXKftvzLdHTeQ23U70=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9648)
DpPECOzPu80H2su5+Bwdrjqpg+kJCqAZqzFE+sPUJVfMO2tTjXJz/zRfCTPRWU5J
leKVFGjntnpSoBZLe/kxYZQgw8UEpAe105gSM2gzO32p/bV5HABdnR2S1PP1pCQ3
C0Ky02gF7IJB18XvIMGbvQOGeayraeWX3I3KCJY7JL+guiSqzDTJ+gkKznTlq8OO
EjGJG89WzFOvEpg5lw5tuL0PkGsf31w2JXEwWKfeOoxxLpaftoRGZO//0webrgyR
g4s1uJdPuNhG0vPYeaT6kDkblj3uiF7O/s0qXGBFdKvozeEsjNcVMoJLhZmtNH+5
1arjk40VgVh1CO3HTlGSk2Xf47/ahQGL6nRp9qFwY/Ez3neXJY+F6h4FApAuLKoJ
nQlJwl9Npfay4bF55l1GvL8anYrqw8NlV0TG5zSr8IN4OsTznsmAnmbF8yqWLDP0
JKbk90jXcb1LrJ+swXqaACdfSVC/KtbCK7yGpgs/pg+4cNGW94mYpEBRVhuPyZG8
j50cRssiyK6e/8sws5sNl39TKSwFugASW9L0yuFxrQUO1qnCGnlcZNLlcu0hxVfv
fIVlOXxAxomCZvJ8K3/nfpvjxDDxysgDtYK2iM4CaG1eyaDIq4rRp9xA2cEPVJ7f
QPlwNp9NuXOym+l7N3ySH8YTOBsQKOSCwn7UNNQHMjrbfele30kf+teWu4ZNHkgH
w5ZwgL8TjAXP5GaYIFGrHNHBKm7Ccyeh3bhxH9FU1Hwu662rfGoUo3EsV39monbQ
G3kk4iKsxdcosNw6wGfNvbdLFWa1YDNbeRRwMgVwmz4AeXbuYiO5IEHbMEh9ECC8
RGct/IApVcdYfG3Iv1L1sHieAh9UIqtWaAeo604tqK1KX6vQiPuC075x/G/eNOoR
1qJlhxxVEB+hMdQRtGz9p+PKpKrdkOI80AqFfmu09lMVf/7HdbkwQThNiy4rC0B0
2ozlKyTBxwj0iopuvjyUqvLracrD9W2PNgS7WOlzxeANtmfJLqpppXQ1r1Bs1l/5
sQQFMNxrV5Ovn/CqHyu7zH8RHVVk39DpG2po0mu27D9/MUl7IhSweB+kXF6yzkZO
Lx2MCMnP1ew/JNEYiyJ88OYutEjU/zOncsA7Q6MRu4MkD9k23pFv//MJTGx47j7b
J9ucL5cmiDsycmTPfe3b04o+xQOJPewZaegPpneba/3LFewAJL8V2ssssNkW36+8
JwbSD1JQETUlmafFKvuhmAXCvS7SuBWU6i27FFK+4hIEX5mMjy4I6ubRIDhAQYJC
Czy7BdQAjysVybRCXBecaKORl0CNMQZqsf7Xgvw5EIQBMssr7ZExfOq5+nB7PYfP
Q+AxbNZZraFQ9BaHGGnWxzoOEoinQhKslE6RATcGeEVK7Zju+KgqZ2OUUknYS/vG
6ApqKFhWCtmdKOEx9nUwJu2B0yRuazaNDil+y0cbYoc9p1U/6rTlQag3s4CIMUNo
BZr1+x5Ea6sB1o0vjU2h1307G0QA6XDod8aqKupacGwRPEx8iRLfLFqw6RVbjgQT
fj38eSJVxYlO29zlCp7A+OQsXqPP9JDw/94Sz0ZDvpwM/esM+xRzPybZs9dJwevM
UzxduhFMsxe7M5PvJ+ACWpVTNkp++LwkeVqld824Utv9bBpDbrk/eaqvHyXA8rej
3jxUDFfGZPVEDD0j2B+6X0qwOhv5PT/Mnu5mufyoFS1kJpwW5q0iYTkVBQNJZagj
hYK9ekx+lA6ONTMKAFhLLigPslhcCqjwggAkP2CzW+YrsBZTnJVbTCS6sQrdIzWj
zzB3aFPMnMKWl7MU4HpVMwq7WcB84bw3zf0W0wW0bvLMbhVbP0dbWzOdbWvrtO0O
kBEL6nqm8NYSHEqrYKri7CZZZOyx+1jQCs1kLO5Rgzof840nPHmGvEj0shRUKWId
Sh91bj7QSkYyz/E8LhOyIFc732RlAKEr0oa1EC7rKfJMpOhkilUEb0Uw41ihcMkI
fVaYw6CD8ugrw4S179e4M4fCQciOJ40oLNtu9lxafaWooWSOsHnEVDZb+Kt88U0O
E603PEVZvOq0fSxrGtzdDsuGdrx2nNulKELz+Emwu+vbmwcm8cID9hZ2Xzx4oH+y
Jk1kN+AmWXx/3Kr2F2pI3Q6m7lIjw67ytdBq9xdTuGAe63J63P/kGw7dTVM4Dj1f
4NZ8U/wF/rhbKBrgXRqFTcht/XlA4bZGheoxKlu7KcG2uDCSRQCyOOBaVFYYlhPb
ZfZUPCT8kS2+FJ292NhDq5q6Qgps6I3umz4zFbalRlIfieI3/S+IC3hBn/ksj4ia
reumflkmIMnmeAHCJcTJ17ogK+v+z4mlTUQ1gOm2LXciuAe7872jebK+o5Ezk59i
S3nz8EpYVsZPNSRo0Vh0enU0slBl4Bw5O13veRaCc5kdNHii2UgSyrC+LJ9HHUIf
J2QLUSt1fV5oMpXjGIU5qHKhXSdUKp/mpBfAFEukMmpxVum0HGzo8CbqIFKt1UgK
cALYUH4XarqiGVttYs0hdhdArsMa4ZYNc4/7XdiH0wNjKsp+71kcEOEM3HN/7MOr
iVLviZfSP/2C8ZX0BB2zoG8/WhEiUj1S4z5iJV9Ykj9Bwn5Gea8IC2SgcZq7hZg6
TzW1WniDxSttV4NH9XblajpkwPf2a+zqEgJOAWAG/qLCFUtNuUTqj+04blHelinU
qgaYUG4JCuMpGwWO55Brhi5iEUGP4CI4YxgdZA8LQEOMf5/btgzg1KGwWjl1Sr/q
WlXwbvpNeeHOmKJeDfSRNvHMRHh1FB7lkHJcahu22UvexVn2Fg8SaR1bUhxRPjs6
CCYo1t1risD9Xj2CQW5sFBiHbK9uCgP5DCRtBkuEL88bOVzmpCBQo5tIDxGZXN7n
ydIpQ+Mux7kIC0d2DrekVigmWDZs7QJxKukXYnjSA4eLg8cg0Z2ghPEjXNa5yqAX
FxGjnVE0fP7v3X9E5aD/MFuoMfEFNJLVIfW9J30WNorsiWgbZTq/vCoU51EkLEOU
chiM4ogcH0lm7SJyV4JDkphqfXyMMxd3jVSmuenis+0kP2PCfUc8irOy74BmeRMP
xCzVREddUywnx5i2X+X6R+5rfPem3VKtSsDhG0x+2g3WIoQwSFIV6CTcll3akjbX
LrH5l3hh/SU7pnoc98AeO3cgenuwqHMqOUUiJgFR+yAEXt7cfQMlG/TjJBrPtT2t
87O61uTJ/Bxi2rbAOLiMyO/0jdRJI9qwJ82oLe/c6qVPYWKIeCStmfVpdnfCnxFw
OFdfXEQjDgR4WxpHUWZmSnZDJPQOiw3BrANBFQLWrR5SWL2RiETquig30kCS/4wT
OfUygXqBZYQKKayk/ZdNgjH4r8Dx7xqIk8uof7/NdQzv+P2mLyoSedsWwup2YjGZ
xzskbtrVqAzy7NTdKChefiO5VRsadPJ/B1l3zmAo0vz9gI60N3W0BtGjgeywR6oO
SnV0LmljTBhrrTAqO0ftNfIkXQPT/4SFxOxWv4vFrPtSedG1IiNDRME8ggiKfgsO
U3L8XXr44sPGFwC/eNlTcG24QGqQv1p/142NSoKZ2y8pOCsZDuPkWxtRn+/N47n2
w5bLOVG/miZfZ4wmyjC4VnMuglqRmWbH3z20OR7py1dwzrIfTM84oJlet7Ggp9F5
v7E/221OxL1Z68qKS5WhZqpCEwzxrX/wL9DdNu1fvy6tnxvkVGO+dtWmCTrLHHcG
cGq1ZXEMcukAW27V6UHq9PAHr3ycElt9Lldra/tah4ghuZKRsv2o31Eou78Dmqgu
C/m1T/Hmory7TolpXJFAeYcNTd4D0z1+slcigouQ89N+43qPFDSIv44uOQg+i1iW
JUgK2cpVQfBr44qAtF//0lkmFi4FoCTYgBC4gqqXjrH3YRuaYzPoKTNIiiprTB/C
SKBTzLemh3tOmZ0EVFhev3mbbU9Yaw7wcBwcN61G647Hm2O+B6sfJQHB6JVWyX/U
037hc4FSIWAv10yQBa3ejCMlUepNV5AtItyt4NQZ0qh24E8QSWrETnBJ4Yzqe0Ym
1ti9t/ObvPd7uki8PSudbkf7PNbIZHVDAts8MYymp/0N++4SqiYRUBMfgKVDBnaO
SvtrQUbLwh0n1sUgHCHz8zx1Fq9n1ic4UjWRax6UtPCCdwaWISH0JwV73wSnlYpR
awEOy72FBrwEk8qRI9C7D/eEQ2iRneCVs3rBTspue1zObuipMI1GAQtquvgX/s4Y
haA5dzNgrtnnLP1m79x2VSWqJPLXXXTfOdWIKrSLoJBS1zIRWrFFAtmJueEP6RBm
TB4HCbUuRBQye+S6LgZ902Ni6xVUU/SjuUNjozZEU7pnY7W5ljNhvNw9o/tLJXAR
GzG3OLgN5ZNKCQu+l4Q2q6nqeiQ+lpuJJWie3ioCYfdMJeLEwfSE85+9JO89yQV4
6lNOJzw5OPP4YcTQdWEb0nvt9nVSHhnrX5vV/+gCLrVD1iwiXo40/KskHq3Eq07O
SG08xRetrTM+4EIvKqMkzUp/u9iNCEONKmLd2/4TfmZvIR3B/tPDN10xtRTywHX9
z4RDChpR13yfm3WdO/F6H006xc2tsFU+khbiKt29BZaMHIjX2qeaESrcn+oLJ31O
7fvyK6HUZUPS0iO3mkH/9D2faYMPdDBKN+HDCRFYXU7JSTkdiZn2zCTMIXJdSkPC
FpI+88ir3f8G5Wd/i3uc8MaVdgI+sFFR+ukxOA0xoHSwbx+cZiSgpLW/Mq/Dm8xe
WQa4d2nE/QTEKGmfz0gpHYfDoWUZ1nJLnguiwdiJYTvCM2ckkvd28bTlgNkno3XY
s+TXG4qE318kvc3wIONHFY7MQxMmSvsvhoiYvhyFK9tRNwxFsbS545DFFivORRgH
gzplaTTrNMUGba1hzPoNEBOMOHvS5sEOh+XaGN1Ahh7g8BZmfod9fe32nzyaYFsj
DMdExH3m8EA5B7u3XsIjD5Uob5ii+42HsYoAj4tMvxLfb/6cL1IB9OIqIFZsAqbM
U06EOF4MYwehhIrLgtSZZg7mMM4SLeM+Nywj1D2tCSro3ef/hdq0rCofFfuHoatF
x8DraM4PVUmw5BBwVLv8i0CStDntwTiLoZGv0qTZAogdO0cJ4BeomqmkG2Ry/jqn
w2Y8Kw+B37Dcqe8itzsqa/a/0DiIKQ9kdpKJmJFylFvb4fyaXwOGXbuwHEAr7jFp
OstGGYYBM6G29s+mec2WFKXBKGluovVhha6+pLzYi3pr+Kn2NzOGH/B35BWwYAt1
tyeREOXmwVsQw8a0aaBy5v1De63ne6sQ9y5rQV22sS3fhll8WkjGF5nue+7rOPXb
HtTQEnEKgN8VRnancXgUt4qYB5EtF0QhG9LUmsF2EZO0x3JCGXVQm4kt3DzLDTa6
sGjHTYnxnYjxFHE+CdCSdZh9EdD6RIuvloh2lcZ2bRHM2O48YvbFZEzBaHxMK9uH
5mMy/f2gOlDJ9Z/wif+ah3KwXdLco3wltRavQb4SZIsy8V18duI06T0b+T/JIpTi
jTOREduWl2aVlxm8vPKTt+pi5FhJkcTYJo5oQlifuu2X6K2Qva1hRnSGWZUAfD0o
+v1D8fW3J4IKn41E8MJXRDwUW3AxnCQgiEyI5ImFknKWuAKgY0CgVlkuLxUCt71/
JxMP7Iao4nEVfih/ckD4K2P8rsSWgbMEW+sjLkykm3+gZAdzMxwQX93HjWRNvhnc
98flPoxUP/ZA+rGd5pbcOwGG+Z1AcUgaYBESxNSD5YwyazdRoE+eJFCG5ZjjWshd
9aE6cc5+jXE/ffr1tpKvR/qIYR0ifw75pKNjC77mmtRP7oX6vhB6BtY0Ex8rgBA1
rjC5n01Gd6RirUN2qutkdBg17vi2KLaPKOFtJ6WsiQ6dwOmdZGbRU75TW8Ou1bbG
Ch7Ai4pti5jona5totxXcZNU2PKfc61ZVPOBu2g7WCD+OL3fwxEPuA7W2nHzaEL9
6Yi1MEPt+4+ERTdymyT8SMnsKeM4SoGHkE7RP64zVmd2CeLbptNyR8YznUKRt/vN
eFnPjX5pkV8tFMrRB0YaSiEwnI+GnqYdVStCNLIG1j4HGXT6h2U4lhH5UV4CxG70
kym6HE00wi2aBEqpxt9BHeaPP1pC3vGW+P/Q7WyJfbuHogSzFxwwz98E1Sr9zuTO
SawVUNWGMTt81DarKK/d+QrpHvoIckmSFAukm3OwF8oNN2m/KuLPzYe/kuzRjZ4h
/gIKW0UJkQFO25h24mrQQn47g61bhjOEhnYGLCzvB0VP5p9izwYfKpjbpgvBX+JG
uBFrJJpyITVuojy7RiWkuCKlQH1eevYTkSlTXemqJAUNIOprhTU8Ej62eT3m6wx8
WS8OM6/QLp3L5C7hfHNLQbAlDWoRBXbKsi63vE8CkLvBLlfmoE+Qv9tUrSMol5M6
weWceXrFE84rCMdTn9pMeO5T45FxZNF4oaeemouEqCtjLnZfmVf6J4cNIPyDffUH
hpiGFmWNvpR15abCmsyJ8h24Q8JB6k4tGEMW5tsLlSku75GnQ4/hzZwVQlC+mlSs
Rz5fPvr05eC61BZ3sVu7p44zSc1razAwZZjj+tsaEzZdIV45alKPP72M5dPABELv
KMBbaUOEBe8TdqJgJzGVBp3kp99na4dmQCuHJyNjhZf2uBdZ8XuVw5fAfVjbiLos
XREsfYukvIu1dWz/fdIJbxgK47WTqgNrf1Y4hQhYZ5aBQ2C7QBHGz8Yi8FJt76cN
to8KKtyK6wcjZuBUwq1/JqjRKlf16QxYXz2x1vVvU8AeDrWULqKTy3+lXcfOwQR/
keyplX71YqxoYWvoV4Mc7rOvnjNWjcML7Oxs8GaK0mo4ie4aqiE7TSrk+OczeiHS
RqtNdZGEP0uKp2dA0PrCH5iiFOcPVzs/usUVn2mVi15ti091fPlV3zopVR7eJ/79
eVJwRyEsdIFdLPngtmGsv/wDt3sj+U9qZHzoVNmEa6TAGg4m8aQplvLzRXDWgd+l
rHoPWSxVlldkr+yYHuv7OkQYP+DZz3JJF28IL1OwL8/b9F7GsiXqNXZdsONvYuh4
zFqUUde0lcBJWq0wrz9mtSW03FeCcY7EZGoxdfbmtS2/WGdg1la4XmNz3rCPoT0Z
h3un3eBFYFhoofZBdEeQ3ZqyucT7PAX0zhcjXVipK7aZNh/Ypk2UacFQRC006GwS
ty+3jDYb5Iewnhba1DYC39hxWoiaRrmwKU0wNnxWFFPteU4ReFok25cGbQhCWAa7
NrI7ZxsLZMkGfSDrtnKVlxI4+rlEgz3xacMlktoWlQhHObj2CLj5gazexbOo/k7k
aqMJONFXHjEDhE/Quvn1ZR8QxIB8tJMpZoWM+qF6s20Vy1OchMPdKzneTR1M6lsD
pnJtWFkZZUNB9RkEv4D0fexWVfyEyNFDETxxZtGnfXHMCC1xEmqLP9r4J0LaMawO
75fq7Fg8ThjboZuAy7S6QmvjjEPDOaJBtq5ln+wlKAxP2pOfd8D8OQTB0cK8G5Tz
8puxKmcmYvQcZpc0ZdSwZoySSlvvCSNdWB0Xd/XiRbHh4Nzn8JacF6DI0gCAqkQx
gChcHDiQx/vM//63hIAVs41VWYdI/XZ9zQTIrUpn92gggzM15G6sJt/28DIpzpiS
ocZBSrYM5QjEIThSuzm2cWFoCzQq/TcivuS4GGIWNuvJxeyZQuvcq4FxgDmCSIcZ
wSEKWlGoHI9hGxpJvNAXyhlpDr9C0XEADJuSIZm5iI9H+4AlKDmumpJVUkcQFw0h
PMmXoJQXfWiiyznnFp6xj3NH2csrBXBwaZxsjQ1EAtOr71aDiueFDe3OVTG3Fd9J
/0iwvbH5ZG3qZR8eR0vdhZzAkt9UbL3pT0AK/zLRU72PBYOZol8eXpKGrKpZTTJP
ecgv1j3YHcEa2V2DpOh/M0PZ/Ylwxnh1H3RHQzf9ALi7lxj7/2yaCZa9uF8X37ha
D1mCUGrczjJtXFLYw6q/y1a0CGz8CNQt4QbSSOUy+l26ondroC1P9L3DL+BlLVbe
JZuH6sU3cuaS+GWszRsu3UoCJRlmnOsWBhq2+GwuoCsmS1g3CtoUvnrdYNCWL5tJ
+m+qZcSdVRuA0bbDGLG/vHzYn4Hm42ccoV5pcfi26HZja4jl1OVL11nfj3CkFMwO
tIkP5i3tQfW4Vm0ePxft3NSGwJwwzaoX2l9tR8A9cBGdhlzGzq6uYLjYrP2XftfR
HJeBz2vOF0FuwTvnK0aL2RkqDcz8nJKkmjgWBx9KlVjlrKDPI4pVQMQXY5q1eZdA
QMxycv6YmJ7aOHPwHA7bNSQG9uk5k+foSVZbthBBqOnHCeDcZ5JbJZUGT9ygNL9E
ei0RFQMZlT0kTnviHHxaeJmZndXNtz3ruf44S5xq9Mzk1C36bd+Zs0sxmLejCoxD
u88HhwcRBBfsVWmb5UKGalkYdGQFgLsGLoIB+N+tqQpCPS3Wv1KI4B7FekBdRFAl
Td6uoEUflSjrwUaFAT1IZnJGS23pJn3sDkilqHDAtrrLYfDsurbIcEDs+okWH9uv
a6AQaQEfs3Q5AwgjQXSDWUqKf8MqIdputsBML/ucCXAOPf66QYHqiOYZyuagVfti
60XswDo9NCXJnv3DQ0ujxQoDwrazZvIQefDYgNOwbuAQtbmsyrkvRgKW7E+EsgBK
wnDQJEvoOwQg+7saPHVARSQp7xX5zLigl2ShYh2la2gdPxGsITD/mMmITRexxDKO
AckWqE04Jt+/p81nM59E1drTapx4cbhmYbBQxJ3Hxo3fQRdG5OxBigZic1WgkkrO
d+aNYVssAFBi9nG+hJhZvEkwYqfe+KvYW+ceAHWKiLs2+AtsTgpryp4H+4hXTkDH
UkYa4hHm2IieQzZB3VAKEiOPoXxHbQD7RSNaSN9D4h8oKNGwu2IatQv8qgsGK84W
R/Baj7mSgM5aTjyxmLT6GurGqmeVKGmNoJy1eaRaqKAVo3wuCSJ1atSjB/7rtvFj
ZG8LzwpTl59P83xm+FH9qzxS4sRtWKHkayLqMr+Ab6jlVfURLjfqsta52Y78MQP4
X7Dc2B/vVrdB/BtyI8UAJx27RpjkyiDnK9bBy6YaUYQtD5kSTg6eH8f1cSAaypPm
sVtgMkv/0D83Db4XGiWSp+2J54Y4toDuM3dHDgKLUJWY2FWd5DJIVdParrlDHl+Y
/zNCUllxMpCqWcqTIqC1CmL2mHb1a6a+ljOsyfDvZSGR1yQRkfNuGb3s0kz+GmCp
IJURcFgcxPeIOM8Dpowlot0Zbjf8Wm1SqRhyP/9aA+LQ2u9I2Er5+unC7HP21f4i
RcraRGcs7ZRPL/WhGKXEwMRtz1ApR92dbZMBNk6d4aHHMg/dcTIs7dqckwluHFXl
W9UT/GXpJyaFHOhwCeCYBHFjOQWtj8m9TWlzzpdGKtrR/bWmpq07GTcvj49LAx0W
+iycyQRTfZJRy7f8MgOC3gs8YIMKHNZucN5Dcx4ekgs7FhaZ+6frJ2pciEWqXXjQ
lXJpdJJ9bHR9tlsM6OyFPo25n7gfdG8ljXh45EjgGo/BCDQuwqx39XBYImkwfoD6
aKoxa0uF7CPCNtTqHs5QmFfWETIomE+kwriHW5oeAqg573hpENhtSe85O08UVzXI
YoiO/v8KBY67NENhLYiiB01czeaA7/R802VV8XdfcW+ooUEWFnXQM7I3+FpNllmb
FgipkVXnYXuA/DVIEN4CPZr3McKRZ5Krf1BI+j/gifeQxWY2U4ciDLWXPOUi4A7D
utSD+HWG/Famsq4NAxAmUzZFuZUihPhDo9ZTBNEQhy0gRuwkZKehpg/Vd8Lf3AQI
ykIEi6eNQ9XGsn9olS3BhTJTNeLycngM7p0uAEVEEhAMCgZWegKGRTRPPEGFg8B2
7Jppqg+eQwDK2S8AVHeJ1rSEBHpdMvHmlODQEDjHRH18vtcTdpJUP9CSDcgISD0C
K85RJsKLq/HUikHz2wJQ6M24yChWib5j3adCkEHB8JumqX9t+ABTkIxJAza3uKA2
YhRoCuWb5weqslbxEP8TO+nZdREOrueXscrC7Ckspw/vy2UouWHi4jloOnx3zuve
/a1SawUXviI16KL01IJ5SgJKOOT97d8Bgy1T4WQLrs3jDfHWYf2eXasv8I3xKykY
+SPUA9drxROeocTgNdOLKZ5w7pzpTFB6D1JKQEqh8AhPbP8Y7hOfOKvFCMM6RkR4
1LSLgpa3WUcl6dNelClprxiiUrU5gMvjopIOLOY1AT9NN4MWsoDXGE/k+I+uYEWj
Pft31vgTYUCCrqrd2x1DtCiVo8ZRKnXJcQriwQ/eE/CmfwoxmKE5ZL/n6rlNL+NW
G2+/UPyT+zHY9GGQYIEnGboLvxNxjwrU+fNA8jJzIlKj2pDZQwNatIMWwCkcA2S/
6NnQTI85m9NFAR7IzedTA/xqk9kIWkErxXwzC2EDu5UCqIXOK0io7hvotcNmEpr9
4tSgaPCU+Ib+F7xFTsSD+6bK9IgVlqxZAYfu0lJ0s+gDyM8b1dRLglAqMJ1SBjrL
uN7rnDz6HKB+QnbdkqS7M9/GyJcLbmiyqiS2uAkHW4c/hN35WX7J8GXFX/z0b0Bt
b732zslAKx5WMOu9BvfPrYtCQSFgANlKuUBLmgAP6bq8J02pkqVfY1O5CgZWo+d/
Tcw3evR5PETP5JiTDHzHaFj5ldRhoAp7IOcLwEmNggV4njm9QGN+nkiTcAEanxjU
ePCRzXatvHcNxMPQ7q3r6SspF2GNVoATRR36PHlc0Y/iXov/zpgPmN6O/Q/FR236
oGbGra8rWpfT5U6AyXYuI/9sGZaBIwH9Zvvauqu+Fh/y/Nk+5pO00A+4gxDl3yuI
RQNsjNxF95PuzvQo9Uur95LB2iAXKl1tfmH8EfsXcqbiuW/xT2CI0efJTfvjQhz6
J7o92zBvfFxJ3UTCTiBhGvSU3SlhGxC3DrntB/Q3Iuz6FV6zwad6l82QQzBaV3S4
MZJHXd2T/zUiay0DgurJVlh+kNJZ2UGltb91DK6kirRuj1sC8p3ha/CQEDuUWf5q
SLaNRIDy6Fi8P0XIb6M7xAqd0PLyPn+UX6V2KzUgIPNgnw8M+djU2bP5lH8qia/i
Uh9usVFRSFGwPqpIA2zpPZGcb9Rj0I1jxEZsX+ocy5Son25I4UcZMs8tAz4LZ4UZ
Jhkj9ft18zA98+mRqimfohD53ltLl7S74KSpgZCJnIslvYODMeOFenyQTZHTd7Sc
w9vSjRAQ/Hlpi0dasXnmcHVEji/m2QrZunC7xRtzCr01vGbVULdIxh51P9QYmYT6
1MASgp23aeeOtixFZlgD32CsY3zGq1KRT90sDdn4PAYOdkNSMdHBD7gjQ+FI8wbI
blhA+xRFb0YU1lwEfIG2iAVUIUMMzVCQvyr1I8NQwWKkfyw6kLvlSNBIQIfifJ1l
AnmWbYjVckNZ7tQow6oZVlqpUr2p1Rr/I4OpoKUBNqzNj84fG31XcpCmkcyxEx9O
Zja4VjvB5/4aYtYaWPlB4AhuwtO7QD+3no7+rEa9cF6n8VYvq1ZguKp6Mc9bW4y8
scvBU9tatMmz2igkQD8fkXGxw1TBP0wCjurIH33b3gMlN/7zc1qr5LLRmWGB5UYg
K5FJnvTNAP48EtTSm6L2S9QoGIkVwhShy79hotGoEHkEPXYdfDyyeWXhU70QWa+V
7VBCJ/o2UhFjOj4AC/gbqowCMHm3VyRdCAJR1EK4jvb0b/eoYsJBWDRPnPpLqClO
uIjRnoHsjlLVUV0aqEjsqtac5EIF668AU4kofOAPLzgM7O5pEXAY52yuRrKOHlt1
aYVKlqmIj4W9/mESIALbaiBCsk+1pIpPjPwTqlkB0X1qRcjn0esidGTsSFwrB2z5
3U5luObtB/STKxDjbzEhGC61jvJhz7POx8jMGEYD0tXPssfjq878WVG/Bq0pKLci
RWOuZ9jydSO6x+ma5/WZCAI56VrevZ0kyNHxWpikymtgpmR7kZDJjxOVlz5Ig15X
rbmjmHW2eqnbYLXuRMLbPYUcgN8etLeeJClURkdbz9xwiN1VChPd7QjmP7fEmZnY
CaQDtwat9Qwz3ry4tLSEB3E46OZoscpBXYXWLofIWCEQKsnaBH6DEhDPDEvzu87U
yKucxLCJ4GRUJbaXXdkFoi25LQ1BjsxAoP5aoiQtRhjrp8XmbHizgT+hKe8i61js
8Xw8TofTOdglGCx609jkoE3+Q/KZNsnHXx29anmBpFJk+t2wD0yBdHEp9IMDWvMY
Uuuc9LZpZXHLtmbZGfnkdZmt4xprfXVS1JztwnphrahGHyIftFbcHtOjO5iyJ9zN
8uU0sRcLyfOkWVeLJHU1jkkX3volGKB8NuB3TRi3TUyOi3h5RMLB38Bd6VkWR6k2
lftkm1yRaYIimjPkPP3kzrQwNMh0LGL0MwZobZQzokklcbh3GxaoEZqDxMVIEzkP
SVia4Mo5sXE/ROHFB8ZsuvrsRvSnJje8oOwVBPhAJ8uLvkpJcUhQ2A6HGvZ4KSif
jG/XfE9evw5sQbS9So4xzkcqhu/KTDuE5ktjFoFxSGvU4w2MpusEVUgXdSiGl/Di
5qElc878/8oi9jVkNfZT7amCo5C8qZN4tUAlixuHxeFnHjuXNNp8J789V4BOW2Rc
krQUhrksKsIKA/Erxbree/BqtZa2jRJ43DpRjUp+4ZBp3ln3UgjopcGv5vhCu9le
N8SFUybHsm+Dq2T6nMOB9HCXS72aCxc3JDx+D0XCU7QYRXA38GjLUx6XZTBZymMN
IMa8jAR0uwjODYICAiytopOnpWAQyueg/JBhdXZ2JStVjlSEv1tuDRYx7np8IBGO
7fRej7nSJbGgAiyr9m/G5JBK/mvyuDeJEXJPT/pyce4LdXLmuT3itYgyKuz7QwdY
`pragma protect end_protected
