// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
e8PrABTcnMFjGpqLsJg62XNmdRFX5z5q3AGtvIuCCtfU6ID0trZnbgQ82jJqkWj2
1mh+QbXOO8M+3YAgHP1EcYtWCAWBTKvyzvRIkiAlE/ent5HJ2dQ6uGQCYFyU32KD
AjOqJ6SGvHgtqAhGHZup16K1q/RyoDtF3tHQ4czv9h4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32064)
7chbfeiLdELEJ09F7Mc2me5FXR8jt1Whw+qjz+M4IZEErvps7v5VLKojAzkXu/OM
/lywEL+8NaYZbBoiWVqrXlJsH/mabkaMmCLfg10KyUBgL19fi2m17tadEZR9JhRb
dEtTgZm18unAxbFKKIw+fxhz7evxV7S+IrD8Rk1nPo19Bag6wgKjCkCVJzk6JLdS
U1mVroAJJjBfTwMyoMK9YMPPVkZBgKxNM2NrPLwhSy9/gxELJ8YySwYKnCe1TsBR
xhU/VqCgZmbmcL1hpAHCB0nP11llcqU6OwmYw3iRxk0FZA9rF/yLd+3FyWYZW7tF
ZgUhpp+ZgLlymqBEvKO/1Kuh8IqLSxDXOfaX5ymohl3xqRwA/yEYlSiyv+UPfoSV
56ndmK6W6OvOGahLqIgtF2BYvtmPlW8y7a3PFX2e2Oyg1U9WjO4w0bQI8VyGHFWb
lGlzVZWXGhTFiI237m/20LeZEqVmAQlN6BsU9JVBUIpI+ZXIEzSBUBAgoA4NwYL4
Cv778LaWNrL7y/Mcsju8iwhpI/Cm6whE0v6aBOCGAkVQb+ERigx9j0hZ1wRww5PR
uneOt+f9HBlJkApz31Y4VgxQkyHKAX0TFlCM+q4HU0ac3qqUdoN3P3tqkK/+tXs7
aHcC51flgaU0mRF92To1WAEvBVND6bC7K9ivKu9YhNr5XMjRlyeLGozIJWYwnUgI
Gm16QUw+wAg+Y0zUhpRnx2XejXQ5rcPSs8JwzVks6kBqtnBYrrsG99gaY8neSSUd
KCF5ZD+MAXAPuqoizYBjRq5EUSI02X8GS+LU3Jh7r8Jeqr4dGqdviLRyIkwBXsXc
r0nJGX5iNmsTpDpfq3CpnFJtUWD9OpZxGq1EkA8K2Co9hT42kVdee8UlV7f4vf25
hlolDmSPt+Kz/enHRP55sbdCD3fuqlg3SGiHUMZFmxMgnAJmJAwfcC4pB8zkuGyX
i0sv3z62xC6PLienCNbsRjeMlaPzIhY4derRz2hLJc/+WaiTaIJ/yb7uNpZpo3G/
x25lI0UT92uA519VVmvnJPkkK2gh2P3phiwmIqzeBRzx2H/9VtMBeCEhRMMmjpuJ
FyOMlvuRPv+2+VD5xyaM17e5BwuNpi8PixfuN1Kr0/g4dXRq636J3afJcPmqMPpK
fRwmY1TyX1SQmNSa/Y3vLqFm8ec00o9WboXMH3Jm8pAfQhzWm/jSV/xN88FG1MPc
NQidOzJLRWPO2SX9nLLE6h1ZYWpXzqxMrAjoNH41VE4NDldAkHHAYoUBUeTAK48c
FFaVqVVeoyUZOkeYldm04uwoa0gRnj3CAFjyfAmGNAxnCsNhzqLogAj3SbbX9Z5S
HC4HeQDw25k98No01lRv/RLIMVXYCnAFEo88RZiDOsRwkrXFI6kpfzK+033AWois
F43eKUeaJEAMtk5/CG3xtKQwL45VG3eJ66eCA+w2Ivxk+sVKLjCK4fbacealrSVe
xncUYti85LOtSDm4a70/7D2kH9lc2dGOKuQ57J4Aq9pEfBOy8EGimT34EwJAlbkT
EuyPGh23nZGn6DFGlyasq0PRRumOmMTQFFmbLKtoNdjf/NAyMH1ZfCy8o1YVyxjv
akwemDaBM1rX1YefIvZm7GDtgcIM0t5b/rj04EEmn8x7WP8zUoH6cAhks6Y7e8DT
i3eXGFUvd8D2QWfQJ2NPTmUV6yxqA+HZQZM+zx5y8xwYY/zh5gCoRisuLy9ly0DZ
WAwant2DRm8nyC3lb55c8W9uNdJBKXGRO2hacQWoOJrGEnhRpvM702yNjLW+Xo9i
qaXpJS5SdbDbsiWshS9lVLqQICqclqe0bTwpcAZYri53sPxivqVik0kuY2plHCKN
HgVC0Ds8jyjaBRcTw02kEHKF8EFNJXv3J4GgRf5onPxvmsjA2Svzax6PEONZArWT
CIkieM7xgLrBu0a6Rc9uut+kBrurTQ0Mi9nS7hYU+q5P0U8u2tuXAQV8dwVbwshy
al4hc+NPXomaS0tTPseTK9iwp7vruEF1F0TLycl1RzcliJnTFcnOAdixk1ItyXdS
0GnM4ntzoUbqtEdITOws9Cy887cJQHKKS/K0F6Mose2Xc72/hQn3DQdqlfJiZeEd
mqbLPKU4cSPiHRqoAoBMqTU+G5UyKSrV8CeIzxTI4GJS34KbQkQWrHXXn9jmDH2d
ClkZsaNtVLZvhd7iYrhEtcVR/PqheXZ64cVU29MbN/M6oM0DIDQXlk2FVpzWF2uB
ZUwobx0F/NABIZWVBP4zB143r1aRzfFAqZlVWiquLv6LYcjLYahsDG63KMr8tmIi
FAkrtPhUWZb+u3yQ85nfiO8C2nIHZMzW4oUOveqyol3z1KTvQ9hzNpD/jODXizEF
wvGgQC0o96CHr4og/3fBtD65iG/YF1AWgJuOQBCaxovNFQpZXJVe7s4l2bOwGiaX
2sVQhnvDU9p8XYVrIU7/GUOdnvooEA8YafqODG54Vyy12Hly8htlQB90ZSufjFXu
QUEHs9XUmaMKOlP76JtrJb3lBV3f9teQLYadhFrDptRwym1YIfEBJsEuB+ZuQnfv
rUjdbnIW6rX91ytbFzaeB1jep5s9l+ZpCGPJ5PyA01K97onm7pDCgLMuCUvbY7+g
kyPi9aTzYLHJXmIoXlfKlrRESbrr4Lv0jlJwx0E9U644FFfXDK9Gok7R5usFmKbb
RH28dAljPV7Yb5NtPrBr+9G3FD8f509LHoreLOlVs0F+Ydzk00j/1bbQ910WGQF5
Hc6uEgp6q59fBDrfidBlIDxGuyS62a87EsZCxTXNhf4ej5DUMdWF3COYtMvtFZaM
GG4GQ+BFUIMC0dNj8o6Wv54pYPF03DfH+2DUnUihAO7XLFYmJnjkAxSe3jTXN6L5
+HF5iVSyAdCtnPbZuyUL2VvO2GSH8Wn1KNAhrtQUu/25ATqt9rj3rjMLNpJtIBuK
YhRlcBmU59YE3Haixu2LiM6zY+fs2IbCFLfyhXNngMvOgZmJAhyTCy+nd+IzNG5i
Q96006ZRqj0nr/4yuBNROIzfpNoK8FQFbF0SL/AJx1RERfEfa+EUaQFoCUsoQX9r
eGtEkVk83VZMYSbg6lo23CKExtbv3YSfx8nVyCQ4mY0kXT/5CC/jdsVhu7VhobYi
a1QldUKlLERQVuy2nYFncFz8B6g40WTquDShksv7rCOB1orqQTy7NvmD4YkVbLtS
jgVFTBWtXTRIFr+wqLadzRJmptsVoZQxNNw9qZr8QjxGgkQrrVTuM6xJsknn2k6+
9YdVFYiXNln4O38HQKwJhVj4ig+8gh2hkvz6igtwf01HxA3ylwEZ3fIwW/NQTEbq
vPEquA01Y7ybZrHpfBwwiZm3UJFND9V6XThB7eGoWU7lBeznNRegY1ENehbWDZro
ZZCO80o0/7jh4peDks8cZES6E1NJ/Tx9sRBVUjQmuBNv9pzGn1hbXHfXK6jNVHdN
xGG7uO4czzcaHV2W9Cl9RifUVALn/yBjh6Jlusoii7e1Sd7u+ODRuHT1i/jdoQJv
fItr257IxlmtpZE2Ya480rWkerZBkS9OR4swN9eXIr2D75LXkohWFbX9+WfcHdT+
sLdiFECS7MWAGzIpx89/tQAzv1rPfU9S/Pgt+eib3r4CielveHGsrak8DFVnoM78
MQZ/uavVqhRoi41uKgcVLa+Mh+avR+9ktbB12Yo9+uVZr15LCt+/0MtQPIUCvmun
F9BlBgdGouMr6eRYLdd5JNDe0POY7OIMlotOOquoQ/TIlxagVcz5MmjBmo02ANRK
xzK+gVFLUtEOnNtconx05CvfQDIfva1qi0kVD6iDdoFAZUS510eVIK8pFjX7mEOX
RLHkIkaL1RPAEIl70Nbw50FE86ZmmmplwvzgUhaGUCpdL0PrDM+v5+1GwKgkT+15
Vuvs8EKIH9c1SDk9T1kP2lUPUG20IDTA9nHBvjNavBn+wNt+wbDovhM7nGc8Rqeu
GGd7Lo05IoN0qgWFbkZ0JmjyOv6084oZuHBw93i++D6OADz/BmVqLywnZt/cK2Z9
jocOalvlUmLVaoTyIR8HL5PLHdj1Y1goRQbIDKKsaXkKiWk70NER9Ke/+24T+Gjs
kJPQ2gffE7E0mhQ0TeVjWKB/rXjTNk2Eoe8VWBncfyMoZFe+bylHsgbspN+eEKe0
xbsx+I9hwNNErPcyfjeyYlrEwepSkD9pIiqphX41sMJJeuySjZACOlVMz2TsUxHF
IzawQ1vr8Pcvq+JCjrDxNBnmmrbM9lQVBHadjYH/s+IlsUbiaUrb3ZDKoEZnJoGb
5Q5vJRsgwhQrW9cU5bSGe9mQS8YR8Cr3vrIlPR/onV/i48KLREx34MBiAGThDfl/
ZQxKaPkO5xjeVcAKYu7ea4wXIH2OljTHDxSs4yfsX/Vsy6aidON5DcVxwRbAktDL
0c/ievnnmGQOP6ice/6UXez2a6P7ho/VJowpH5y32rThnuV/p8sqwrSLV+0yva4+
WnOm9iQ96dIzXSs82M0N43/55rOqC5aAbj+swi5f9pWf2Y5XbPr4O/nsV2MAkE9O
9UWuC4jfNqucf7ieJ6m9Sn9tzkSwyR0YIeJzeHcy7hUQSak1ExbWl7tUDQHGyS2u
SPkR78X1jgSCy+rkSfkZqQri/x0QYK7BJbSF0Jz5CsdsWaXJYnR9qvzlqfmsry/+
nvaRLnQLWXcnF5flvkQYuoWjsGSi566xTUrSxE+HIQ/fNPSQSyN+rPw33c4O/VYD
Xdn9NbMa6IQWMWnyBug9Jax39McozAwkD49Oh9G5unU41wTkRa64BrbV19jbiLkd
EleLzUHQZkWXMylmU1w5wthD9QBBBUyrZDehmgt2uIag5wNA0UGjlb3AxuGspUwI
8tOMxWE+2Dg5hKfDh/pFz7PsJnQzvXYu/FdjcI/GNCdNgnTDMyxULLwcXukshLcr
JYyGpVYE/XOEEkBB5c2Btd70h+bY3/lONBKa0Fp8IcGqGoe6E6T11QrUe4zPVOvV
qUI+WM9xjgjp6fcJG7fMCE3ahIzeFqa+PHQRAA9r+0Yhic16bodFiLRHxjCi2w7G
QBg0cnVCprNQJCI32VP3Pa6oemwzvqhE9mQH7oBUN6lS89sT7CYhz7cDjO2v/lM+
Pj1SEU5JBCUsRiS//jvQ7JPJyR6i03bZvUQ4GkmEjOTyIV/zU9WeFa9OPO5bGyOZ
FkHMbVDvUgXeEFWezgxksTGAx488mcA86yfP1ozT6t6ZumEk4QrHBmQti6MnhN0x
rhDSJldqLihcdag9oH75bDskSdlcEjngttcMvvaudQzRCSmZI68kZpWqUa89/fKr
S8UZVG3wBrqr2UeaMhAu5RV56UMoPBxzBLhKvBuYft0kfHLFb3S71OeT4w7XFhRE
mw+b1drq1vgm3m1BMXqYD6j/58//6PXujsAQnEHYKuuRre7wcM9RET2i9zBadVD0
1n1+ggbV8wism7PYhSNdbtWypEAP4Enhz0GK4/zIEAK1Ux5N9t2yfiH699Dz1mcn
QTectnYevzQUZAkRCK0SlCclPeIwUHcIBD7/VRtXLSyfJc29zC4xnPT2yH5dR4qh
3kMVBS1cGX4PyaoKlDeoLq3biIp5iCMdw8mhMJaStVGSZgmlKKgDZqwNVsnsweeX
5LEQQlJZ7Wrhp3owqku8sXMxcTCa/mfxrFmzQYrV04LmQmzNvbMqaD1cYKDX69s1
inedsyk3UbDTCfaixCmyl71WsBA/1w2RS6Y7a4ZNSqBgjJS2vcemaLahghQRrEBM
r6CXN84xxhhO4Kt4i/kyVCpDTUpDsIVRzTcg/ec8Zl9JdDRTY0tKDBhi7u+0/fLU
a7C3SApMM9+/UT17nFVLP/53/T51pKqHJtbjI7qv8AzhyTUfwRgmjofe2jDQ+xp+
G1PH3u5xHUFLwYAMwgAgUoZLxu5SFVo9AlwT7c3O2dtLqRFVdKnEAy6LQU1R+819
4Iyux6oBDUFHUUfpse37us3T9cZ4KMOmNg1aasPDApJmtQXDvOzQ1qCD30kcu3UW
IEftBzQ6Z8kcLOyUMq+E21GU9x5IHDYd1LAtHt0jNoGwxGvCdXY5EyQ5Yw48kwHY
sAG7OXlW1RMymy7sYwP1RVcY/PRuog3XYqwGieTEdHvlzRtRm7fEhSi2K6ugd0hx
QlqfpS6TN/8N4pzP4EPzrnBiD3DORVKeQWoqer7/wQid59CdUICScZpHqZzYSyKp
M8AkcOPOwvTfeXhc7OuXJByzGNkzJgvano6zpJTwIoKNwu2AKjOYsaLW4k8PN5ZB
3N9oX+JfT7e19IFgymzFwS54djvg/kz7+AwQXy65PuZ5nms1Vtw1oFkkVwSbUVug
kg7DME8FgyAFzgNHYSUAX5+lv/Fmwf35iH43ef+2QkFVjUsxPj963tfq4g+Qh4eK
H6cvEwCY0OmZlLosaaxCAato/s9etm6BDThiNq9b1z8Zkvm6FlicZlCzwm065RLw
IiRBgY8Cx7wyKc3cvIdyJGudJdPTmOxeZSV8TU0yVX8pTGijBWI1Kt90FqDllX3g
Ivjy/7Hr95ZGnJVLWWgoznWcW809nNrWXBi7WXqvSkzIE0dAlAPh3uj8Go+A+tHK
RU6nszYi2y8ohN8pBxb51deV+wXuxfOJqJvvVb8w7+2mQZRj4Q7wICRB+KAWc2lV
m4q6DCFONQ1eO9ufPcBFHPG1uvXm4mIaYTTYEnsAecCC94C4kW+dxE9vKGjWRgUo
f6vjSOsAxy81Zf7OKNRD+g5BgX1gcKd+MozOCT3o9fC7UfBpkQgsDUcdi5gaKGxM
SXLNBasVbhl/P5U8wRnsEYBd0ywTjJKVcZ8gr7GKC8UMxqjvXasl0kkP8AmoDGQV
lQqyK2zzM5CWS2RhlDpmyrC8xSOzrg1DxQUtemzrMETEtM/v6w7En7VR9ROGYQsE
wKPR+sSDXenO0r8MMqIGCnDviOU3HJVknSe9Aov2U+aNUpqAnua33IuTqk7iAO0d
xOZ95A4r56kgxxuKtLnR65RFWnc4pocFZLnJ9RK5StUN/z0/vFRQ0T57W4wr+hh9
Hoj5KZocC9RRE3utYZUw15+p3NOnnggVyHLFxWL6yOZUsYYiuTD6j42ZBowCZ+K1
V6a/Gj154/SounrcxhYJhkaY/JWN+ozShEW4KyIoeE8wltJ9jDk+sQbbZl203dqN
TdLC9DKm/TuCNOIblZTLjs6JxcRIiHUb+ue8CRgmPBQppexSyAn2TWmqr3ehD6vb
qZaXPWuvoWeXWCtsOTe3l1qk9cU62EHmuAaJGJHO1E6jmdgSUHTRVIQwC4+0Jtsp
2YzxZci5uhneXklVfWpRJXJOSm5Kh/v3dmnnVkvbkH5K6j1OW9E2M1baQkTGn+Cb
k/EIXuUzNrrCw4wIIk+wOM5jSbI5uX3dKBAqxC0skYQK0szVPEczTMekyruQkc5r
MB9fNDa2GEgCaGQMerDi8d/9DkPPd3B76nLXamV53SzqSPvBJmaq0V0uYDnyvg2W
RRaMoJOBqSLMLRvmjdR7xTEVyin0NKoftyAeDWi6oUa554eQlPAUmAwGNB6vBGhy
uEfbSO5nd8tm/7DvRdgDSWh90uGRSkajmkJD3QqI0+uxHjbwifj9GqJhDTcPCsSY
js6/4oROzCIR5lb2mMWlSvHO8l9kMZCQeNQkM8iHWYy9x1VBcN6VZcSB7zl2HeHv
xZ3h99v0/izqMopEDizWfc1OXy60B1MAx+PkDgDev+9u4pvmRIMWY5qLJzszfGY0
ImTgcEBp/B7U/JF3VoWklJb8ZyWb2gQVuiznKvFpMSEZi7tXQKVM5y0Ojw7+eE5M
m7WCo0XpcNgf1SdDTXUxXAHUK1tKqeqqmttkb/hfn0LM9tJQSTbyOQqmi5yVFkaR
qbRBJ3KLYYYVOKZMEVsiW2AT4WspWMhQNWkvBnHUzz+LKFDoqLv62zuLOgMMDUyo
63eNmurY71rXss2d6qpxRzq1332+TVnFwwJL1LakB2Lvrp6xQqfr29HfNB4zUEA0
Kh1sBkUBovCDqgsE9FwBX1mZBwOmv0L0+VVCYZsKPsI4EJ4vweq0logxN+rfP5mQ
2pQVsQnpGBcBrwy5cU0MI1rXD6UiCof91a8eg0voPFsi5UpKgiiAioXWHVyNj4gL
yIj8HixxVkaC5mV3PMIdfoNIz/tl4RRloYFA7oSQuVXUxLvI9xup2Xu+tFwuwyND
JvK6dTMG2KZUQGJsmSBBE6rcgfX4KAm3vL6dVm+3IA0LsT/2jqT4rjRGrh7adhlb
uAyxYIbO1n1rTfM6i/iejKdOj3Ra/JbKrxIdmIvS7KtV+hFyBh7sgW7h3Yk4Fuq4
VPyNbHezhZqnoIBSqp1ietmTNCYpLSIjHAvStv3tZYYq2fq2RQYphvIRQPCVJxX6
0qgCt4r6UZPItyXuzY72bP+9TfDmYMLNutYk9H6t1CuRoFwXBWI8TOEc01ssxW+4
Dw/Y1Q6heedEPmzCVoUR8ldrJHVMZSPtgUglxn/XbfCfV3hm3WW9Pl1dJeQ0RUex
QhYEORyyIUoe3wnSayzlpK5JAFeo83AJZM8ucOD/DoAhvCYxVoT0UQzeUKqBUPgO
dijHIfUoor5Kdj2IAyB2bjDcYjh/v9eC/2q786F8o5Y+lod/JXMWj253gqzYy58I
FJsHWEpjrPNBb80YiaC2I30upKhJHpX3aRETODpJ9dDP6rHCwuXBFU0K/CDMlKBF
3idGpRU6TtYpr9vPDMpcxwgt+NWVAc3LQTQYBVMYZ2K5majY2bfiqycOpwx/wRRm
890tmVtzLiuYKCL7M0W2ObW6lErv+5tNiJ0Bdrl0/f4Kn3tGEwsRY7BOgUs38CrS
XEPHxp3TfV5fRIJA8Al8U886yXhw3P9sM5J5LfubNbkT52v4GpRKUGUOc23xE2UA
Mj1/RFTi09LgzdaxCmDgJYnIfk7YUBoRX+AMhFstvT5LH9pcENpqm7AbI8txv0pN
w/aNK8uB5h97w78ov/EKS2w7hNYZqV+tG7sbBW/ESDJsph64sN41PqtLSYqtYRbe
cubE4tmexVevnnGMhaVEQs/WfK57h3tHrkBiPiV2sSAr5Q4qFUvuFnSaApKN4FHf
Mp0HQuz1NyRKTcXV1//Rsy8rE5m6o3ZV3wRyU22DWxORsLUi/sVXij0kmp8+hoty
Mxh12Qv8YHula02jF5HEoOmiEnmHRZw7XSUzYloMIp9/R1sKV3LTPZ2UjU5barjc
PRVzYTcMTKkFexl01NGOs2EXWyLpkXNPSBqfyO+9EiweK4nubqU0nhEUY+m36+dC
0Q/4sEMU4C/bWh8c9FuSOojaiJTA720IDgW1p6MimtQ6gqonz2XRiyvopwfGMP7k
FTiB+7I4kmY8RoezguKpq1Ehkjus+yNya2kvgPkuRoBm6/AgsEb/nRdXY0oDJEzO
6sCpFC+lrvHcZ44tMKJD6i1FQ/Fzgc2tggGJhCQYR3h4ojL01aoFR2OquvLKHsw/
vXGJ2R2du59eKil/rUBxjPDCQgu4AYq5IaOpca9DyGybsF4cRH6VWI7DmbyMQWdw
cWSqVI9M46IWH3kKFAN2lQPwkbmfjif2mHBifb18zbkDLIlzuhPHYMrXL8qVcxoZ
ZBxJGyitgjHQUGkNyWeXGIpvzdgqUltyI1C8lJJ2nFPhxWSlG5m7v3SaOQm8OQf6
HA1Xz6fvrW83hOptyQGmT4cqffWPcf3Y7wwM0NTSRFuhT/iw7eVUu2GueijCDZ5j
qVhcQILK9Ra2VH61809j3w3t9PGKnd+TT8oRy834K/uUZCjMJ8pFguFi8s8JDXup
qBX2gmO928wbNfVFSFS20/5l4MNpFwVKHX6nOP3bYBwi2YcaekM7pEudepI+Svn3
OdUSsCqCyFmy/PI6BUpEaFSNXejRYjhFprjnc9lTchrszSgJNlYd4tL4dUNIsxoJ
nvDpfq/jtZ90LF5Ue++km7qmv7xZglTym+1jEOFAmZkRYTEPVLHB6K7OEz99Bf+M
IS1j5LExq/RXwWxb3Q43SYwfuJig+MdGsns7z1FB2SanMBw3u26pfTsNBIfDU4/7
9t500Dr+WvN6a33kLWIbOkVauh20Pazv5bEoN03NtdRpICD643UPYrPYs/pwGTFA
osJYB5mXi9rKk2Qf48yr/m4gmzBn4N8b5SXqCE8/y0bdE1BP/361vQmh5x9ZVzTt
SIWwM1Te8cr4E4D1TXN0GBH1jxkLthmV3hhBg9dz9SoaYpCGfuN6TCpagJyVdU3Z
4gEI+9jVUEFGE3mtqgXLbgqzFrnGYDiY0mATPxEgLuti5GU/xO4sl0vKVpUofVuB
FsRremcjFqg7b0KLkMjRyyO3U4qm92kyzElOU0flJc86xqJMyndDQRrl4w5WXqiV
IIl2OCnudXJx6vFyAmIYbh6QjwJ0i64PDPZDZQDwB5ondotyixZkSHZFCOJ/PF5q
hB3+Ubu2x2FSd8N37KxiGuAdHCJtJhTZvCpeiLowV9hqP0sgTuK1K6aQnuqAhNO7
JoLckBdrV9JdxfzJ4pA6pCe0Ab6vOZimsH6KUmGEYfug54A7yulsA1lO7U2KD7on
otcGczcUh1DIiTN1Cnue+BGLhbWKF+f0+YUw+45Uyeevniw4a76c2W+WwwXTe7vx
eI8eGh24AETGOA3k4n3DGMRmw+7OX7PpqOdvDau0OSC9yMiol3X4l1nK48Gky5ZY
ceyc6nyse3jkRIoyacJOgw1bKlSaxZI6QFG36sS5UeBritIvokgJZ0OUKPvFCUtI
y6Ij/AxAkCjk7EJFERm2P83/unqzXsfdu2LO4sJoOiyQwVRZlKiV2HPdbcj7HyPt
G60Mtq4A3BJb224SMuM53zmbSWLUKCU/QOC6+C0IhDBx3LBNBBcEvg5T+6i1abo+
6Aj1pM7ge/XFR1mpqUtwg43L+hGITW5DgGVw2ifdCPa2H/j1WD/fO8GAEN1NnEgg
SHVe/+dFlhavGg/Zhf419AuDEopmzN54PfGSVvsf0WzGfjMf8raZg+PMchjI72j3
E9YWsdFJdISNani6Su9GlgbRFCRw3zTZobIHTBI6zYW+/8ICnJvUwzsHHLKnnmrH
FfofpDLCcC2MAFI2PHbg1NSNotEJiEyka4vZw6CXJrjdeUegCGQF19Zpu2nStXWP
Y1KKZ9CKl/fN0aOaBUto/kbWZK2ubpLDYfOTpo66+ir5EumRaScaHxPbdJHkBSuQ
3309GHnQzG0ayBQPQYq9D4aMY2HIHOdvsAVmFtuaxAAkOwgn522t4E15nOb+nKc0
xmGuMbLl2RWcgztvmOdprblBF3q+TgaE+hqU/orYIIZcNUM251I6VEHy4mK6Jk4p
T6XemM6RmW6s8VE+Yr5Swfxj6KZ3sJbvgkPxQb7dvLYWclGf1XeVJfSkJt7SPY12
TA3njw2oZCZ5zBqVaDu8iOtzV7ECQkOgfqGiwNzwC6kpicgxloDH3QDM1zI3GS5R
+vI1Bqp7cwtPjNuv7+wQ10KcQ73HXDV4JbRJfgPC18GmX0f8csxSFB/8TpDY1o4Q
AufMplXPriPYLIGDusu2AbI/N5omJAi4TrwOrwVb4gM5iBKaynaRGswYvEiuG6MH
jiEcXQFPfFWGSwgm/XtbvwfyEQB9NwVjlXA+VgqLZXEwQPoKVUnK7A5ROSML3m5V
LvJQrNYTpo1U5iZt70RTbjHP/we51bdjZhfjWdmmVY+n0po5vkSsskd7N2ai48ie
AMWmSHWGwp1KQQj6Km5bfcI+atZ6LInLAIWavk4CNC62m/3pSU3wD3ufSUGgOFjT
r499UFbAxO29N4sk5323fv1YIsHqmW4Fbv6n+7hjU2gHYPYebJsSmWEE/+956xnU
JycYTyTNgrHQhEgnAInJ7aHnYpLGPtwOPwrreuVmzhygWmqeGDFa2rgrVw9zg1EC
P90ME/iDifv4kERmvo0r0MbuXL8kCa9WINjvVIrNtGA0gQGxDLLaZhYbTtu3niNe
tR1F+9OE8VomHTNEw7DpjXWR08DMzgeho6pKx4U970LhHRSVRzC5trcBkxg/JzF6
MO5V3gMY5PZv8cj6Q8f496xyJebjpwWK4MDkXlPuLynOtsaBoeUUuTl7ANgb1yQL
l4P1LyRM+JU5iYlhBlF4czfxrOPllvXVHBttor+L704nnFiJc3I8Azp7OzvXNGqC
518Y7xOQDCMMEQcXlmQPzffWGB2x1NUKzRb9kMjk1g2mTVsfHbdS5w0S+iKBUR02
qmYl6++KTVThJ7hWDhASGQUjYfl2u8lIatCfL/kkYGk5C7vREGzjhbC2RpknLKiu
LVjtUlBtKSd+GF2hSKBvy/hHer85HLMEjKEG0HpUE7HT7Gi3AgEumP9Uxds5GENZ
K7H8N++GfMCmzDrc+RVa/841IUVcKg4rDhZJI/nL0AiGT6CYqdlcgOqq7oYxzDfn
OhegxvaEvpFhYNeunTWc2fSaOgNpxUaaC+Tw+dh3qb/a63JZJ997V0qT8EAoK5m3
8hHkfC+D0AsD/CUUebEpzyLSOJm/B5paL42tWTST5r1uEjebIOHFrKGbcV7D+PjY
BSC0vbUI0hthY2erlbUOJYgwM9zVHgmDgFCBcYbOHrSjZDTM8PRiTDGFuWSSWypT
M32DNl8JSMRhGRmvos+WvQDVyfc70WSg9xYuBsoIdtH3ZHXQzBpmTlcfkrXYiQmL
Q3kM6yaYraH3jlUbGBwJ+ALfBi79f7ejNv105iGQcn1+s06UrlLDg2MqeHH0JPED
8Gei5siz0XWS+PNGvn3Pq9uYbF5e2R0BAw4aNlYM2hcF3++jFCPTCSJeNqRUH+KR
dMI8XYUxT0rn9rap+io4W+2pvubOGV4/lou3z+7NniriP52/zgV6ItSsAwIQeJiO
40rrwHBAUi4zhJ9c2a9QJvEoKChhnsvAbO7PjyVntMu1TbB2ibPE1w/JH8mctDDG
LeOToij343v4/asz0ZkdluGZrk2ANUflDMqJ/nCEWrdqFYhlzAWmLvOBPI7o94pD
25ap0Di16EjxB8+8UzLaatHMONRIc92g8X4n4q8mMzRhkOnundwteiGZMOOWugN8
pYe0wX3m4qxZcoaAj+2i3lc56vBxTTItZaJ726P5kNCJ9js71mbcxnVdNnQdKZ9J
25yru8eU2iiK5/BxCCjhBdyd02Fx0PP3ASmfIJ7h24R69dAgZlSq2d1s46FsmaNk
671DOQ8VDYGVIGwpkThNnSe3WgvXQOAK4HBTW+oHZTnC29tO1bWpWT+yOyBCAMm3
F7hNT934/Znds2CogEfAModZnWgrAgyp0fIW6yj1ZiKofV/LWWTLq+zGNSqxZSlX
XCGsUJvep0Z4RPMHC1aJs3ryxskPgkQZOXqSw1Idzb2nRi/zrjqWQx/a7gRKEKqL
KXLiL/JZQfm+3c0KYJzn4r5mEXVexmfmzKAK60IiufwV6jijbaB7/qZyTvwkVlXC
aFQlPUglsk7nCwVO0w6rXlTC6nPScnGS0Pvr+VhgForZdflESFxyrDGrLUNxhx3I
NJwYHLXPbw3YUvXMVlBF5/1aSxGz6UnCBGBYVSwyncatFYCBGYnw37ixJdhbc2/H
6BqE5qX5s82mkzFFBdKZX4p7uQi5kR+sdBQLOEjDed2D6r572geMQDyShxNpfVGN
8h9d2dRDq6BABtDCTT464EN7hZdZIYBG36iU1SJflbmck4ryi1nG65Lk/I3FuiLN
vHaAtzwFOtDYDXhP8FpGNtproKLIqz6zP7bvC9nsplVgu3uuAGQkOsg/n+ACYPSx
f3KP0LGRA4f2Cuh6iYeaiMksIdAte3P4G6d6EsKM1l80o8sgDqpALWGrJszsyzvU
NKGo/C4r0/TTZNbhif+LwOgEVlb11lnvt10TwDh3TxVculm7uD99fMC1EGgY/NYf
T+FkUT3quefarZR4e8j619QgaubR91Xei9l9s60J1SQvfordrrHbZhCDlaeE3rvt
+iIjoY5AGu6J1E3iaUnz4XRa723qZWd01+QANuYKuZeIXsXF2lb797a7GubaobmB
XxWqCzQ1/phpwc7r8VZNr9UJpfNu0GX19j4P2S6SRaA/U7cPyt5RvckJ2+R3Dh3p
qdre3EaWOtuS/b1SoP5BmJvtasno2KgbXluipRR6+ONNnXfa6MsWKav43Trf0luo
AGVf17CCk718qP9lmpVaqCN0JrpZA8Xt50807Z5crxlB99u7GAKj00DpITw373eP
EU9iSZVWGIKt9ow7IjlrHpDSxUjbva4bB2+0rvsf1JSEOHa5mb+ZbinQf6ne2QHt
F4kRkVvTEmrKNf+2XmE4bBMBzGnD1Pp8HoAs4gtux+v/yRYWcEZRURrkjt14cvJW
WLqbUg+HBjElpBHFy8L2YJJmgUXkmGcDs1ugcAdzAh39xTCyhhyg+ONNkFAQAQyT
Nv+TFgdIZ7TTKI0ceMDuTqmkYtDrJ8bCU4jd/uevZhg1+LVVnFnA6MqKDp5IdMsa
r0tRkW29Vgo5QbbcNYTmvLOQDlkyDP4fZCLlpYY+I5s69joQ07V1JsGsEVHPIo7r
Qbb9ndMN0wJSHxV7W+Zq8lhSTUeoR5BevX8mG0ylAw/COSCS5jsiZ5Xona/DyLSO
YFUbvfgFsRA/XQZCrOsyU8EKq2DuoB8mQIK1hUWh1hVyTwiAyqclpI9nAB1gOn6E
8312Hf+IJbVwuKj/mnqbsDN/gqCulcEosbmw4qJ1Ffk8o9/TR30kGgPUZSIgAMOd
2xOdcncsDfsHEXYmJOVPRfgShxrAIkMcQCN+wnMXKkIPOYhNcVLnErIMV9/Cg8/J
xNvE/e0hDeR2VaIgwIOFOspt5WKzXckm3tmTbgxrqr7C07N7/MuzsAvE0Qw+iUgT
EO1OkbrEfpNn2mGPIIH6obipPuHGpkRWDc+BzMqdmIRZ0ur+LsWUzRTji6oEPz0t
u+Xm0Tzut25tNilnlSmQi2/0UnmwPQArko3zEpX9LPDJJk44f1bCdNxZW7odmQ+F
WyDOQ3KjJX7GnstBwUWFnN3epKXnGDWam8BBqSRiIg9UhBxB0JtH+WrkP5xUQ5s4
sCh19L6275rrv3+z+MZkcdy12yJToVTqSXEWNPOWuhXwO4j5SQrNIgUrWKGc8oaZ
QZGN9h+vgLSHzIX0sJl8NnhLswbin13bvf4o7gR1yD4lUDNe6RV54+NOaVd6jt5I
G/cj5DauAL+sTPGDpnbpSgSke0VK0VpgaeDLJBemGRlh2tbixJwnsVAmsIwZzZhT
HspvdOJG63duAAhMSurx7weBpT2diWImmJtyu9/MZ/GimnAchJ3TKvQMh9uqOAX3
YjKk1zMhC2s5jRuofm2rPQjYy+4YOFFl/oJWYjPXlCYXllSlc3D2V4NUBoxm9yA2
1Tr68VTKrEDz5FbvoT7aMwJwMOaVZ1gDUqWGpZsU6YwCMuC7S+tFWDHqpif1uf68
Ne0OklV6+8gBIlXPpCLJC7TFasyXDFiREPV6gsQ6SvFj2Yv9KK8p24522VBcP4Dn
+Q4zfAW1/QMVxbWo4AYpHKk8EHLPS/IQKDBU/k2DwX1/XFCBVbdo4RwgKmhVDi+T
1RpB0Rad+b9P+BgqlAWDcspVYW/PCIqZe4wE6+h+8KjSJgt78smwFors0QS0l0qh
SkjeR6cwXLSoBDj0a7BaN/Ml5P9SKvUi9BFVakURG+TJ/ZE+3soGj6DGNHxl6XEA
dkWgdGiaq2uZkVNNFkfcCfPgfRIC7VwHaHcrV8YQdGlNRJEYLzSsoA+AEpiDlqLP
3IO5O29aByqoFyBSzvWaf3XkuVw0dTLrzoJSeedVKQA+uH6AE9wJU6nG9Un2Zux5
PENovzOU9bBC3Fj1X2lJGPAKqmH9kvN6K7Y8rIjp1f0xkRacyhpmrxqM12dwHM7U
3XLozECf3PN+5R/EuG2K3/CnJeoMNzeFike5ld/KuQ/S54rir3d1FAf5uLflATp6
0lpOUs3gfner1EpLFy8lkp1I3XK8B5OUqhF6d5+qELJLLexVuVqoxsSSjUdS4bny
73OXx7BB6eqKX9AliDS2UwmwwzENFiBqQCOgarPxYaTzZqKa0kwHJImEOvz+tVv0
EC9ZYNbXx+T1GAV9NyNq+ht7xG5qDMjt0HZstcTEAVOdZgNDrubJy91HeRfMuAP8
pIORUdEj9ANMiPVOSSeYgplCiVKEuLEfEZPT87zV1dSiYciu5nC+xPyxfRKR9sIv
Dbl+u0SiciwNlss7/7Q4huG+52JBeIxAAMhKWHqy2d6c1ox1j6WiPz4BuE2TvQNp
7FE12NRJBx9zphajWUipvcQY7YAfLwtvzm8+N37qcSUiKBcOMIAOsaemp89EszMX
V5spXvrmrt1KA79hyyU0PJP1TyEhUc8LEaNSPz8Z2uNyxI1grofWmB0V+Jq4VI/g
JOUOBXF2f3eQG7aMmSKlO/38x8eZm/M7SzwCCGpG8ZHvlKUsyZaEJJbIUJEsRUyZ
htG4BYl7f/3+QKzow4MaSEu1nJ7RZx2fAbUzNr/mlQ9wJbWhvJmrVz8waB0PbhNf
+29zTHpXIvNBxtcUSE4qzOxAJ7AjxS2B6H0QagXX2MK2yw0BXIUksKG3NOUy2PCo
iowXG0mY3w7StS9YPaJvd7lWoCFtljFM/WgVusTwyOZ6AmTRGWba2MzzG5/4bcan
1x0Nq5mM216FRqymKj3EqsmqM/Bp4IH2jBc524vfwufVYHF2mV6wKqrlqJW9XORT
cIyty9melVP/IxSWd8vOBFaCl7DjwOafVDOd1E2/hAcX8Es97USb/Cm9tFwf9pt8
QP3GuUV3iaBKp+Et74jYThxd6jmpVeoG1EFlCjzMrI09058wQYAjGbAKjVGzjTx5
rHlsvHZE+MhGXwU2HJgOMlp+Bqrui9IGsuJHE849gBeK9mS7tOc6xl+g9e0LMwCU
YwEEaOpS3DqeNKpAjvu3QrMF79VsSQdA+mC2zYW8Z9/Y3FXLgrZ+Y5gcSF4I1WQu
5WlkhUv42JQBmHYLhqc+45xM98LxUhNnPCwL79+hClMW9s5Nb0ggbCHizFHjYj70
TLCeiJR6ocEC/HP8mzMaLP9y05sDlGxiELSlqeu2/S/6LcYi/VXmzSBZF5O3hlKe
M99sFiLR5B3M63DG58J6ZU97F6u0dSSK7bJZaTBOpP2maIyhC6wqIh64zUlIeD5E
JD7aBxX4LyOOfaxdF9zjTtA0eZfgEAQXSwvUwslZ+NgFU7cKOT7iXsjmtoEjj7vL
nFP7ZNfn4PipN4FZRvHR6ynfrNFdbQmPZVZoAeVD5TOn6UA5wL4Bpx6mrP3x44Fi
GBcIs1/DIvq/MOSsRuZr51i/h25mBT2f8awSwXzYu9wj4OufuQ3YeNgRIHh1/wgW
ByU7Ovlk1RYwQ7UpEH2PGKnOmi6Ew4s06/fiWzjDS+RagQlQuRpJ9/4Qlpl2u5yI
DQW6H0oOLmtxdh2zfpNi1e+kfUPTkxDhFOv0hSi0NNL5nEFP3cChWSX6gtjr8tnh
srPLh6gAiJBBs79oB5lw32bXZcCyyRX5Zn3RNyUYF2wHb0XK9HkjbOJiP8oFMV+U
M9jun3pLjg8VllshXVTZApbDfHi8MugBFBfhpBmR5ID925Bulfh0PcmkwrD5jWdJ
2IGvHXj2CLgwTr2fC/0x4D1QnMdCs3Cu/EuNWEXlDa6L9BQYf2a+b0ogP9cO1ZBU
l1DD631IOwoahpmo4cdOIoAbIQ3S21pCX6PxsQVC/4XU+XLt3dhYN6XJoYsCaovH
8nG8JhIkQ82ja1LJWj2OZ7HH3IHnribN+Gs1Qt7RPdhcJvBLZEQqbu6vXzRpJOsD
W2+NIKrOOSjUPr2ww4GSk5zUHtNkmZYTEMQxiNj47GNyMu13OwvkS3ttIwVrHKus
LgUEl2uym3FE8DSzeqeC3xnrdHxK3k38XFnwmITUZC0Tb9jZsE3YyOxXIPDF6WRI
ekpiyFERnAIrWhddUkysYvYU4uX3DtNO99GMi/MywdH9PLhitBYykJEh/Ja06dJO
GugdOgPZhfjJKlxt4R3z+BMWy9HpIDKhiyEhxIxF3rMieByeKWmYXJAW0WOTM9p6
yjfYRlu4CGAiQ7dspTanKE1Htrk7zJeCIPpfgr2EMnkZybBINq/NiYnLRcNtB7Qr
i4ksQCU5q81WJ3JRGRFJDZtz4GmHL9U/fdvGY4OyYoWlneT6+b6teowF7PSIcoS9
lnzoAlp7G/ZFguJIKNm2S9V+9HSNLt/1c7LCP6jyh9+S2ODxlU86LxgE8rPfKwgf
ntCpzlctC/2hzqkNf2ma6yPTkuip03CUDySCeBlc8zi41xr2XDw6g0cPd/tXOrOp
EKA4bpxjGcobuYq+uUu95gUabM/pxG3t1VM23AxJDBanNMTCdtpJz7j48Jw5NB2o
Zz11FgquZ+mVQvRCpzqW9BJglbw5RHU+1/3Fm5qi0laAPcCMT4l2ZHOgWYgpjX2c
sbf7iiz5v4P30kfJ4i31gMRl8h5mO8rscI+O0zp8Rtj3ihXK0TNlIS/0ziswACo4
s9IFM0w05E/081lhupW0pduWYE1+61OdqxEe8BQ9OfyJQroRZ8AbVvO/BwcNoh+I
eQMQD/rCePcrm5TPAoYug8y6GQVyOE0DzDrES5uZ5oEXFX/c65eqX/HJOD0iVQpv
KbWrMpCi+3vljjKIApvokdGP2TbROFiBbjgCrOh+ZBIeLezr1zFx3uCBxyZOhY56
WuBOOZ5D9wBv0fsZQ/Pe8D0jRMx9Pd64tH/cB9JAT+zG4o45fsABWSxp0M5rBvKo
T2hjOHdL3RUhNzHbmelvHOL7ECVjCi0WPYMBAtWAzeu2S9ZuWe7cdDtzcla0LN6B
PzZLV4r+V80/hzeIVOMb3eBgYWoHpXk2eq/2Cn1umtYubNp1iR6umO4W0P80Cv+O
rFSpXPnPUoe/rPH9ZffypJmpp3GDNmhGUfx1iMArInfpuiDGZi64bXWzBxn6WYOL
2s8V5fVDNikFKEoIQxVYi9yfRn+QQAy1uXuuOgrVMYNH0omYjUg7DDJKRCZOmG4n
eCaK4haAuMqPcFxvuP6d1VsOH7G88xzWLSpxQqnLtMEGeOP4ZJ62i9oFRQXDd83n
JJObEAkoAufd0alOOJnIMhulP7BFR2HZr0Kt78/huly7TlABXT8HQz3QHpMrzIsb
R4AG6tUQMo5pRnEyuKNpDzeIl6twPDf0uIekLlYDnG66H/KVwQo1x/f//+oTtCB9
spJU8nruNZxcnYm50n5yx2U6FshJu7vSwi7q0rQOUab6oetSrSc7yM7VtNZPc901
HVcfYE+21+ECkEV8m41I4A5TeLiOzjYq3sQeoTSsDbBVDryfQEPi89iMMAxXDHKS
p86hMaIF5/EmC9GRXWmElZ+GEZQcqzNDVC8JgpIw12pMQXJtdmwzNqVtjcVW7fN5
QCuf3OTeU2ojaqCttrGANAmnVjSDuX3nX8OWrLOdEdM6vZJMbV/VtnFbuKZB6B8K
3uIGGItha1u6ehwqMmHJfdZ3ITHNTooPxpKLBV92Yxneteqgr9NaXE8wU5yGdQ2s
vJAMOhFb5QoFaCeUNYWOvpcgxG/m3Ad23iAc/O3RI8Gi/MnL9/0IFQUlAmtdkFyO
jM6+iA4lAltm7EizU7KwzopykWTvss2V1QPr+CgDxRATV9fQTIqj5jHdaeWJ281j
2TjuBN6cF0rm+MTmE24g3fqZ7ivxEIKMWsYvvtd+R8pylLeuFI4R5eI6OU/XVs48
b5PKEzPx5O1iUMW6bd4EXkpUTrq0b45/LrP4neG6Qv9dGlwN/GO3KSSZhHNubR/a
zgVlZnj+AyifmNEVZOcK425UW407z2T8UFu3boDiw4Avy75Jsw3xBhPCuCRHIJB/
YAES/Qa12ErRCAckbRwf20tBBoPCHMSNsdmGoEyrsy6z/0jU/NoQpm2hRuQVUGWE
udiU+mV/rlwiCygmSY9fKeqGwq6ESutDDRB9gnXXH7ANRuk85DOoKWZOrAavc7n/
RlIm5UOwX07A+JWSe89XHWViSkdvkkBpEOJQRtV2g9G/c4IIBPVuhlTmaaLAHyaC
3z60ugPqucJrE6CGfJUvyO9yuZg48IKXnPkhCNLO6w1fA8M4wywxeCwZfd0Hp0rh
s31RlZ2MgOWx9acF3XDpxl1+zywx55dPR0t102NQqw2eZmK4YEhrocUUiuJE8u4j
v4tvBNjYyxaFeSyxxwVGciX3rFC0hEOF+JBnRB6kvM1JLm0aHBHH2sWoBuLCFceJ
HC3YaUCXTqD2Pe9UgiZ228grvsR1CFVZdy6XhDlHjEIbfdaWkKWdIbNeUv5EWz8i
+CqqM9rSa+IreRYVZtq3U42K1qNkNLMuV0+9ysNvVXGjjkwe9sy1m4nh1VTpi9Xn
8MsalVGtmL/Wiik+bk2F1QRPOtZCj7m9XsG/36LRAzqwtc067fsRLWUftZuHIdZv
mx/iIc3NSG419dtwbl61KHzGN5pM22F4eNPysPfqSSSN7pAYBwsf5R71bZdu6Qfe
X+sfd8CvayMpqOf3sC5HewO50O+Vmy/I3Mqd1qkbCJbyrw3eVpAEJHCcNxRRtnjF
XC5DBXx3vuLeHE1fSQfqYBwiFABhqk7wyI31KgLNqGCXgv10OCIKLbcqYDzuasym
0XtZUZMtR4yX+sWvPcn346hbiJ6APDvLAm/1H7LGTxf2QzDhHenD3ITNXxixr1iB
WccygjKyMNqEvOBt+CL7egIWfRPl06LHvJm+k/53P2LIey830UYL1a3DlxgCSyFC
CeiKUkaYZ9ukyLSUv/dKtP23gvwyBUf3eLcCNhTKxrHlUVbJkuV1dMsrvN9Dmwnv
TSg/Lveeu8QXz7FlWZSdiBb1llgsyliDaJjXrAtvq7O3xTrqGCdKMI8rQmTD2bHV
fSIjrHdJg4QRKVfFhpA9t2g5LoCsrPudxxCeVnuRGWy7hTKpk+9Nz75gwGFj81M1
ohl/W7UPg8coJmCZH38MIlhq4cZ1LzQbn9KmrrTNubIJxXGQ9CUv35WqhbBPYddb
4kJjNkVzZlM7865Y7VZsTySQkeFbL7ansW8A1PpmwNcMsDPL12/Y0JSyYgmx4pdM
7bheo6vjwhtK8/4+C3Hg//KOP4nBkFfw8sWlnYFCgIeZaTjctcmYjOBFdkY/p8Uy
HiB4Z4hJyn1t7bELJ8DeX+9qkA3/2GGcvgRhWclzXplbQe2BPMoQa9IUScmEYaim
cCcTA84YGKUc4AxAsllYiKUZF8oBVHSSKKQ6u5qafJ6w61VdfXkougM3QSBS1kbK
IvDumrAA8noKa+zEq/a+6Jj2/1/kdj/kN311LXPNrRjklQ3xkB3bks0sJPPTJJSK
YmN5ZTqWHZK0AEzjxZBpY5kQb+zILp2iclI/SYj5n0+WJtR83XYr/NBmPTNMQjf1
7q3KLWCpj3uKp4m9hHe8vbox7Ul5uVt/+D/jFwKOmEq2hSpePC/SNrBetQglDH7A
nzsvj1MJrfLjVFnZ7oa45cduGd6Wkzu05tiz4X6uML+Dm+I44RV71WenGaF+s3vo
oalEPClhcxX26vE09VlNUNA9+zGEHcGa/rbOEj/xTJm3BNtzLYhmUBm58fAEN+mU
HVVjd04VLt+pdxhu4Fl2krTwOvjLT9SCBjT4O4lhKAiexsMBfWL4q8T7QPU4TD0l
gSEeEv8QrMPCXXzyjQHFGUAHuJUn0h/7nLZy3/RM3SFc4XPV7Q/d6V+5bClYe8vV
NGSQ4izpF20p4MZiOtSLZqn/66IKRCQPQfoqtItAVtDzhLVHhxKhHBEi/MWE4hg+
ac6HbgjJiEjBIM6A3Sc/73MOYb90MyBFeIaVnBo3PDJYL1W5MUCQoH/5lpHZ7NIW
qvt19t5PDC7lX3JEOkNkvgk/c7AjQKLq+0vTYHjLrmM2Nb9jePf6VP++7PfRdfWv
PkEXleV7Xwo6F+4paLqTPSeybG25NrfC0fGiexJBcmEz83iGIiEH7jrRMoIDdHMT
c2afgOHP5hPgldzW0Zr93qqGHsYqfuueg3pkoYNStvDf5fXx5nl6wpT9PE+zZEMh
nDvxdhK3CQzi50MTLZ0JnkgoDai/dto7C5n6sSS49vgmIm3/mwS5F0KzIIjguirD
Of84EicFxr7hcOfcYFX51LHawb/WuimkSiOoejGL0zTKI221kEx/tlYnC80Imi2o
cJVUdHmtHuIyNWJm17+bP7kuws2gC+rqHMlafU7hNNEJPVZkhUTphPfbR0L0uWgV
TSGHjFcmk6T2M5znD0fc1ukBXxrj7ouKuzCRUyVzX8i3/5Kb0InuGE3r5LO+KYc2
oSS0OUjYJyh9CeVlZuvB41Q6LmHlrgDo20USBElw6PXmKO9hoHQZqLGuuaILQNYA
S2XxpuC/2TUQjDFW3KASgPBa1wEamNF96NTQGI+l/FTmyv6O4KJsBmynaohMVClB
z+gGBU3p3xpPqn7p0zexE/rpdnEH82PBIeS31t8QAMU0HBa63Z3z/EkEkl51IBAc
Fk72dnLqG3GLMKqD9+AI9P+HNPgv5ntp0xFIr4oLvYDG8y60LJuqvDdXr94Jnb7i
1CwUr28yb26Sj9Dq7c0wM2IauumdnWpZalLEj86SGALXr4NZ2+H2MpSZLb963xea
rFt0+a5JI+2t02PAhZK8vfI0vKEIQHA1M38Quk8wG6QxbuGZCkd/fahuCPOtEM+H
fccTSD3X6Mn/3u4TmRTFvQszqQlLebrBumZYz4lqT6busz9r86Xfcdwpf5muPetj
bXoBwPRHIrpg9gcYPCmOJnrAjKqobEc1Tb5JsfBMnpwErsvC+NZlRBOEYdDq0V3O
qmWWc1aXuQn7vjgl2J11QyNmGKuggjOKE0VSL9f1vsKICtLUu1yl0p8BCoqJ+r7Z
11Kb7LL+ALf0y1ZuRQ88TITlZ/1lILVIHgxjxDvgwL17mDMPkwH3LRG/E2dgWwYS
eGAijVZkuztxTux3bpnB+LlcVrYK8B9vHukvXvrxAmZRH2+KogA6M3kDTawfvOmX
rj+6M2JlRUzAEKmLtkoUtUvqy4xww7h9Iy87NSf6HFCE80OIEFlA0bvmkCnpdFd9
2q9SN/2wiDV5C7k/XeTKmipJiG5VTNKm6JtGvjYLFL+gsLk8RHrv869fgIUBOxGv
9qF+9WxrUB7HZdgcKdQPbv5KwIJA8CVTCH6hS+WbWY3vp2HCMV0RhZFJzraiN59X
Uhz2flFV2w8WQ3v6YFikUQ61E/QVf7iw/owoJq5oILUvZ8i/gmfAJSa8dACq7QAp
VngWD1XXweweRtHsZEybbTwhXVu3/GKIPhqDXsVa7sji1P6juusY4sL840ZwJ17A
ZZVppm1A8Rfu0W0I4fnb2+7O8jK+d/4qClmyA+3giA3I0MS10beRb8/MBdM6u8Qi
FljTVlgVGAjAN3H1EaVB1iR0LGigQcYkc5D3ahut7ao0hkOr6+81eetzosRizfCr
g0Yu819/DJp64h92L0C+7uDNqO41HKON0cgyd1DiZQsk6a+14ydSfQlyghfNZVRO
RSjOHhDwQ7+QPGekEY4LfA5v4pHcZ04XP6MnxIFW1M2e18ZHq+1fG/ZuHrYLVq++
dqvC73+vDsrKyYTii6Bo7rjMnomfgJbjW094rnKGGOji4t2/rcnvw7thWKH6o1LF
Uaak8tfEaLDtfGePyrVd9DCRYj44hWKZre8OVxloOCO0TFX3U0aFdqTWlCyAMrp0
fILOf/7blgko0ob3UWM2BCCac71YRnQpeftJpWmk5/B7yYY6TslcwW7Ch17kpOcc
GBbqnar0YmE8Ypa3elD4S+OnosTFxzg5bKSn64MxSC+6YWmohB3+tJS73Vilggww
yvlPVhJV2KkTzmzGYFTSOcS1AitVWtpDsKGWji/1B6Jxrpr/IE73zKllpRDzob7C
KUVLEkJVXK+c3yllVvMXLhiTlZhOeRa1LUH7I3tI6MGCdPGObpQ0OiIIsrYUDbeH
rfu4285dOziTJ8okWvPvVbLJ1nd03w9jYQHC2rrunlzZVWWe/mU13O5gmxyHyVhM
D0nwguVDuhj63ZqaakBuwzfZTRZbA43CVQ9Z62+rjUZ8sPMQDzb/17Bl+E+lU+C+
lYnQYvYR+CU65LpiQUhvvSsx2PTFQPd0XHOCHOpDWvavkNBntkXPeC1Ewmk1NnXD
fGF6Sjg2nvMn291UQ/5s0g8WAqbNiOWHG/vx1bT+57XPdwSAhQACkoOOWa3289fM
0J3y9f6ZFXaXu+7X759mjmRUVEdcMkkYMZmFb8HYBeHaYNtxLc2UtjEyNbBlvPVS
Ze0KEIaByFVN9I2EDUhJRLwp3o5i1J++HKRsHaOvL+I5YfSombTNVcnkoK2PeTyB
TLndyn7I2OonTlQGexUiEbLX3VBj7njfJbTSs2dDWxOyYeOrpvFTyTaGpp3VX0xo
9Vs27Vp4YpP8EBhkg02BkFzEAzg3AET2nrCFUErL2pipKoO+QxUBbb/YNczW3g1s
PGn+mRfdpEoa33Kep99d8mJB5Rw2VV3X3z3f4VtFVn1PjreRbGi7s2KTa/kq5qFF
VJF3sW5mJo5nCmIkbXKqYtMD8RlLE9rmVbmsHmjm44DgmYD8aos4x39AnAkzvBwV
9Tsf0xBm0khU9uPFEKrxK07MX9mn5zMsNBSO5RUGBJZtr7TI3OIBg+NgbZEjM14d
pXcaM/YeTezsujMR68Sefe2ZZ8AvoAWT8yCdMOQrZnqa4yBNjlaD11DOe6ZLzeF3
9YPrf1ZXEvcLnpNJaXg88s0+AjsodRLU06aFEGXjUus7zWRYHUidacnSDGaPaX8s
r2pWaT6IRBCTXb/EvlxjhQpoqHERixnQykdokkOK2FYVKETn27KOv9eABumZc3py
aVrk3Z/UlZ+WhkV6zte6uaLgMXrhZvxM4aY7lskEXZvypYEAU0A+Xal9gHOLR0eA
SgzIq0oY+VyJCOcj664BQ1DZeZu6f0YlP9UXpOY3zQWYTHyFw5DIblCIXSBwcmf8
F67Tw39wyJ6OO7esTLANjIVaCP4tbhVRXBAPMY2E6dKfnjLnS/mI6FOdrtKPYi/5
5RQzY64gpdJ1be0iostCaKuBbzoFV/z1zv8XnJDsEYXL9kM5Tt7LJhoExKb49+1Z
9FgOHekgjV4fx4KXjsu5/UjOH50+JOPiZ9Gs/AbkTcrEyRac86eWqpZ3pBINa6Xv
KzxOfipUMIl5PTpPqTqqCpYHKiICGy6cwPB0F1HLcPLcesccHem1N3ZAF5yKU1Xb
cjwTYI5/Uh+HdYD7GUkO/I8JjQcu6wSDhNPwvnEL6R2DEnlhMVXdHS9wkAnUorYF
g8gKM4P3qImSjE81e40I22lH7AECaQK2nrvPfagu93QrjXzgGfYjfhN5ZfRpxNJx
4w++e177D7ZyPWM43oS0pr9kS+2/5gxZTmAA4KjfNGzdJS5uJubUgnZ7STRyIIgP
aA6Z4R9wzVyneJUkHrx/KSB554YfVLJMMAya0wj/+wGlXWee13HO9oQY2lDGd5fb
lDoAozNbrJYv1//Zi4UmvcKWXmzgyci1TyEzz/0WxPkCY98vcuOU12LsFmsjU7Qt
+foFEoXkZfGOIjdRJqKXosbJbHexM8SPLw35lqlYYGFjGKsRbCTEMmDcNAbAKHPC
YnOPfD39+uJ6hPmCOrWGPZGFNgJ4AeWCOqaDhyLpleZByETxg9VyZyhVEAwFz2j2
5hDgmvnYlb+z5owaCXqfB5ohkn7e2/NPFkyLBTdrTCf0RTMZKbjHyuWYcv7j0RF5
nOQZa8tUvKEti+Eh6481WsVHv8+Iqtvdpvv7XP0q3qCuU0cuJonOhgE0PptAhndT
uHTT7ckoemghOL94yRBUA+RQtOIOd297U9cnICNIwXkshae4mGDsjQntJ9oiWNpK
RctlEq6JciXduhpLI7BsrSHBHVjj1AcSxPkQMoHQa8TExGZdLdpklLwKz0OffEDx
gaatqeq+h+lMgpfLrLeeUoe0RMp3LVuTfbRQuO/3NXdJiN0clsJTPYf6gG0KzzXX
4JGF34tBusj9vhONVBZh/Fe76lcyR6DaIrFn/8wZKPJMBV2wkllKQKwEQWTauBKL
YmgGAzoPQPDlFAo7Cm7ljBqhu5uHYqjyeledRd/ZCbmhxJD/LkXR5uTMZDG20Shb
KAqu/sQdTA34Y+d6hAYvsIFzQ5xJ5vAtgZO2889kVln1aFfTO8/CrRxJno2g7dHK
jaSLumupCBFTY+0PzNhmufWOrJFPXXf9+bonougBoIJipBu04iUnjkPlEDQJyOV2
xMMcQv/YizEQxNBv7yKkHFFpKvPLaMuXLOCPCLks26d5zb559AoEhgOG4k4hkKD5
OZ6mxuMSIfmrUPLj3SHnWkvwTTyNuW4AZMlg1nF6ZeyvopV9FwO2ANu+7sRH4YS/
sTn3k8q/3CGo1q03v5y7NW5ocgMLuGERBaqFmGdwBM5kZf62vl+bRrez1dvdToqg
wKCOtAz28NyN4wMJ7TsG3FhfXTI4T/BslKMYjYq2KA9v5I0gamHp98qnvfO90ait
T/dISZ7hgDZ+GKtP2oCKnF0l36UxxhPUtjyfTQGG6GxRFDDvEg58sv7TRXWo3jz8
W+42xfPIO34iaK9wgCT0KNS5NigK+Rq743/aP8WzvMS//U/IPUGIl2s889aGVJmd
FceFPmUZFnOW3fNRXiMBHimwcpUXbB2DGz0JqnpnGVUMKrWNGgaRlvHXVVWLcCVa
C9H1OHCFYxYBFlIec2rmywkU8O40mBrmN2XY/v2KF6pGTluEUvsaswFDOnTH/6am
UQoJBvPPzsfHufYu19OuJj/+sV+7VcVEqwj+IclM+SAOPQNwUHvf31/FDTVWjBz4
DzpxcWFGegbWrelgjit1IZ4wUQjzpUP5ekHD9lVMsELwpEr66eeQ7If9Lo4pt54T
scOXapvZoRyiGVNvRnZMr8zBJutUbthik3v0Q4f1pQvLLqKTWkr9GINlMVvH42li
w9PbtTC+6LWvTW6EepHgTyntnEpsrFVj8Pqi6K4TCQ0IE382VHgep5pv9jpfcPBh
V2l6Vks7ovXUmyfm3ehNXfooqIhdVro6U/l7LydP8syAhuvLlJcW3tnKNkXIAJx2
m63XiQM+6ThI8tRS/ekSl4fhyS3ViJXsSXA5qU7EIG4QojfTBOJk47C58Ikwhj2b
GecPcmdrgeqQ5+7gNvVivdggxqjk5qXkmBQ1gFz8qPRkkazmKkuVCwxcf4exehp+
Xa+bGvX/E2frA7NI5MMvoyXxP1FpNbBl31QEZOeeoN8bcmJ1Wp5Y6cY9uQQm4cRw
PIJLHXk0V1ZwUcGmJZz27XvcodRdRYo30bBUrZ1z2VXY0X97OgaC8zrsl98X2IaF
zoy5HU1e4VM9jTwdB1aq1iDfJRTQkk9yB1X3n3eAmsrmc2Ffq+Sb2e+3XxGUIqHy
xpvcCcq2KSG2zMcMMpMPOxDS9NTgGOvsHvQ6C4lf/Y8Y3Kc/b0mB1G7hXHZQMNxu
CvuyO/wjBVwkE94mPdAdjP4jN7wsHTNwUInJk0t5wVJZXoroR5SpT78GJqiYRD0o
8uhg+QF4r4kzKuhjM0SVxwZ+fDhWc64ERNbVoYa7rN9olau/Bvx3ea3h5hK5pGV3
XqI/CvWcLQ6TMLeAL9r8jpInqIlQ7eIL5DIFv96/P4ia2oM+AS4VdMAY++NQv1pG
hGGpWQ8sqcDgSSRh8+jb6JUFVeI3i/D4RT8NWVjb0vKgB0VN9/HsXuxHcqpBDAh5
zWJvP87hhwzm0VY8QE5j+93ho8IanRHJ+Elk0Ag7hve5+w1Lg6lLKl/7GiMQcbbR
iVrPx7lJDq+TJezvOQbz2/qnP2ubZEzYpHq69vG0sGL9Zcfs5g7g4t/yce0P8z7i
7j13bD+waMQuTK8StV7KrHq/ZL4sHrBBxKiU8pa4IChu7fgdHg3Os5cSheP1dZRX
gcz5vpXbEg3hrYTb6X8FqotDkFiIe/9Ke0g9Qr/UjEG70mi+WNHS2TeVm3X8AO0G
riwEZaI3vGQkI8JNUy9eTBsjI6XlVjNgDBpKZluKi/CJxzdcHS2441DFEPYFCC88
zWlvliTp0zj/m6RRQYeRBozdnNc7Br1u5pvpNTETnawpsKmDNCe5y3XWX3Ur9phB
EkVCdu0wBdzyEzMNRmKK75ri1PSpTc1m8Q8iAN0jx7PjQWQh2CC80y7e971oZWm+
ZRayylngLtpZUQZ7ClhIAiWC45/4v4QJz+706TSey/dUE/q2PfxeXd8K1Tensr2g
BT8zVv7Gpg8WhK5npdzwgVV/uRY6K4P4HMGVxg/MKReVAevtklWxRG4EqqL2sWC/
+kwoJoeoRLt5Rd/j8g5e36Nb+WpE3M1wBDgpO6YCT0PEipBqWExh9VMOa/m2RIe7
DXGoprnJyUHgsCztjjOnsYSCAinNDcXXZurSHouusFRAqLfkbQLgPzWaqlNFI6Ke
NQJ9HJ2JxAy0Mz/DKSuml1nHjvhzDjICwIMzos19TwCxkmJtjWh1yxgqh6dk1Lwa
C6QFpmKNx6rdLwgrIfLBrdpH4y9QDynDpaQZ9jkwKS/Y+HChanIVkOkn9pusbitc
TBTgRG68BGf2R/5LOsKTVjepYgONuL4afEzh7VibnRdpye+aFn6nRebnl0XNrE4j
FJpX4CZiflwe05M1/kYP+1p8DJnOaUJ1wMUsZDlPkNzZb/wswvVnrs1R+Fxf0ygY
a8f1er19gk1kZBUVsW7jENfn/64bzrBSQHAI7Ogd6vvQ67aBUoMAodJ5GRC0xP1V
pr6aqkx+FpMKeedpFO0+7Ej+ZIt9MCl6Ty1CIOb8plCXu1XSMunjm4Yy3UJP/QG5
YM+X51NFpp1HFo6dg2BkYmJdXRBH1mKz5MgNyi54HSbptfzCJZS8yXta4Ct6zwwq
E0FJC76DMJYP+Ht9Vtr5/ghkpJYoPZY9Pdywo+GgW3eMXXRo3PoOJYyJkpO3GInv
8rDe5yPY26I4NA2kRCTwL9/Ufpp4zFKdlCg+cvr44zGbgS50rxl1+K4MSVKgY4w+
zpZWPQaODUNK9vKp3pNaXGHA770MpOPJ2Q4tovMJ3OjSSqj4QTf5mEqzJSl/Yyin
wr+GJLL4BIxwb0el1ITB2L5DtB9+N/vQwTJ6B9VS8fLb+NjQQ6g0lyf78OBURqEO
4tKNAGK3OtKbv/leVKp3IztIuF7Km/b/TsikdlcJDt4IIWcJpHgIMdU5tAKQdvoB
uvqkcz0Di2Uvo0LRWJ8rtwmMNq4GhblNthOh5H6bH8073c/3YF/pvC8MakuqN9IT
IRVHn4wJBmqkF1Q0vZolwvlaMoF9Ot7pb+XkF36+2BqcfMYm5GQXfGQmcGfAYgD2
RDHziyycthIS355RrXiBa+xV25nKZE0ODL1lSh7GYXammnQJh1OyJt98WWwvWSWj
HB56N6OuWdLb/7EdXDR6nBgERrFs+zAUgdNDQt07EH5Yd0LyFnpgtYxP2/8t6EPF
t7UliAbonECbUSZ80/UDIgL335G2oZmRmtIOQA4J97mbYhtL+LMqR/EW65n5v/zm
RzZTttLStJUG1WGam1qN9sGId6yBv/C7+Y/WEitvsE5XqgOSShSA9gebV0w7wXYI
jT/lci9GdKowai408/hRGTzXgsz/9pFQ1VvQQdtayCA2BThbVjgUpMAyXZr6Buko
Ren9seFBG12IWgWazgMRDqsAgfxL/ycHGRHHZLW9Wr6SMimCbMxYwYrLl/HBQoI1
fZ8CawB+fR8THnX4VIpHX5mvNZqd+WIsEI/5P5djVK5VC3hBG0S0JgfdfsIGefhk
AAUIzis0nZA7PueE5cfTqh66j+M/4AExNSO5xqZ5ykeaPT8Nn5WzhOuUCnT3wmXY
VbeYRMLSUyWnii6YxYAD0ElQPIyPBpILg74gCsy5Qnzg/kJVmMn+G26FafLBMA4t
Mvziwz3xvJyiEk5Vt5Noh5rK4cfhpBbnBOpd6OeNy9mtgQ7w7s6XZw7DMLbR40T9
rARKWkwfIdfoTLR+OPs9KxYY0QDDiyRKDyjESQYz6Tuoh6pT4cq7DsGvGcvcYn4Y
kdpkR2u24HZS32ZZW8/KaNEPV+Ub5T00vloFYCQXBsqlFx47A/jj+LTU1zP8Ptq5
YlFIaOlGMJDkPHxUZOEwhO+D4UmXxg8OR3nn9Jg12wkfEf3HwWOVU1Pcxw988YG4
2a2td5L79SbnbibzKvxXFJqja2xehAhGt6zPJZf+X6LkMi8jmte0x2HpLFwwK2L6
iMl+h9BT+4em+7IFMQjIyyUhlXCMCUaAfZT1XvKT3W69JJhibRNlbyXRREtf9wc+
o2LhSOD3tfNDvgaPPYd/+BbUAD2RIKvyec+nGE/QjRad9E2F1qK5EY2rwDvyriaf
EUUWax9FEdDg4Z4Fjq5aaisvFC7f0WKdEeCzyJ207Li6CH+omeOkUQ3TYgmyYm2R
cAMBjIdEBW5vt6DGzPAfV+APlYoq+N6uQOjHkJk9P/i9+HTmWjxY/zpJDpQsH0Jo
sqKCSRppOxjZRtFu5lj5R4sBhxcTeF8HdZ2uyefxNvfidYeT+vFyWDz55uj9med4
+R0xgjxoJXeb9Klwk00x0gqGkfP+LDG7ughjTMVp2q0BaDgZjRxb1ekb/042IHei
t58RPrFoOCs5c3SrtdLNS2cYwynCF9nQwjwyIC36w3xyNxUwTW7wd/ZqIeoQwt3H
o0DIJnRiMwnaBd5zJM3YLaNoZhMpxGfBFD2alWW1wWa+qLNtHeO8CuUBBNa6yV04
/GCsam3HJjU4QNN39wE0zd1NpVmXsm9BpOEgN0LqwDdlEnaSJjKx+WIE2Ua4WdY1
Ojnz38m687R/2XhVwiBOIVGAv4lxEYxsDVi6zQx6S1sLUjgVtjCtnPu1CfGCISh9
ASFFKMoLvg5c2QKkVEnZ8RF8UfQTiHzF+rJf8BOotAmd3l42i9922oubRbEWjjg2
VQ4zrFIZWB3qQ9S/ffKBUztu33S0/wnBN4NRd0Cke398kjpPSFlPZT6/rvYLmJm7
dUU4l4EC7PXp1AcpBQP7llRzA64tIrcEkc84Ge2tb01o7mhz9gLEGQhSK6DMaaW/
Ux1kSTqr6mMPw1nVaIxBks+Dbcgea8s+zJmxfelX1JJSndQf94KJEpsWkV1KxNs4
Lgalt4IbAKuFKx+DS3RjFLYWtRlNstxBxRiM3jDI9KDIQSWkXmNn1/fp+11HJ+9i
f73X3BMTtyHCM70QFVgKhyDX89NzN8DC4DMPfJjNKQn78uJ9xg8r65brviHL/SdK
KaKlZN+aY+olO2B4iabrsAp4DQ7J6JSHsSTo49jWfnfLLGQIHkqLX0KlrGKaVGXp
TzwIuAX5naE/fsM5f930qORI0S1Z3MAyr9y+UDL4EohEDirMACBW6MMn7Ovss3fk
6F6DXNxhgyx9vOfzWpnjdshLEfR8ddJ146tCSJHlKrGibVPR2uVlsYyhoIHlZZ6b
m105oD+vX9ZSSU0CNYIOHMNZPGSIzxUcchIxAwNC2ILp05LTTV8oLe5TKWqWfdTO
RXitC86Kz+Ojkjk1mvnOkrknx7AmFE1UPWelJVwr2R9vzlp5rijVwYJDBLVtvkYK
si5iXaMExur0Y89aAUmOURPbYTC+4jlt3HQG1tHLn4DfNohN5sBjWZaYHzxV4xBq
/nnWMYUMndQsCB99C8QCtV7W4LQ8p4sXAFhDRTU4S4GHvV29z/ot0lPlAw49eP6M
dAktBFtVF+4vejDpu/T7QY3iUxKChDnPSKiycTH6mMxwCTOUdRe78WCU8/IY94DX
QomH5mZVV++TnQDVhNKEfTXnhTGNHjzSyoBxIss+hPugiPhQb/jslxZpBxgIi9Fs
fZem28m4fYKL06OQOCMw4o3tOgWcnDpqAGY/ajcQdA7BeDqgWUJV3dHgZkcjaxBf
IXQEHYy393lA/ziUoHmJVySmtkQJOTZBEn5rI2urZkX9FsKx4yUYLcT81h1xeqqR
y4x0HByqZAS/h1sZBOBDcdaGEemmEhbYCO39/dNHbUTMPfbylihWhdGPAo417i2A
H+yZNGPqHZzta3GGE5JXP1gU6twdaoMobK5SI4CoQlDU/gGERtWZnthKQO2f4tD/
eeFwiK6/6WXUztwWGLmO9SoQ+PY8axhLPfYMgogul11rVjWvQVWHVg+aXwPXpg/6
23wLICLZ8UXHGukn8Cx1dOZSUoi2eM5KRuG98OBlC5rgYH7cWkQGsTJ8EHD9roDK
Bgc4HiAA/5FqSUuJu9Boq2sDdNRZy2Gs9C6P59rbUstLAeRVQr5eRTDneHoD1jNq
QDq+clK9we/VUNa6LVvqJchvPyHWksExI5XhuJVmX2pjrBQRseTEMTNcwgrS42UA
PEGOphurFFlIFkeZhe0PEtPGFVtxpL7fxeaWbYwHNKP9lRlNb+Bt9tnCU2nqK8Fz
ZCksr689AUAiD3woy9EUAvVb0+CcbCp23Uzdy4kaM7Ua96BLCj0id6TbBOHBepDU
leaJJ/maYcRq2/Xg+6Fo7npHGrnh0SAw75f1t8Q1ouQWYde/gfRenIo89a/7RsoH
tiwYoXMs3v7jWJTM9NHGrU5JWp+L2Vp44BUuWn49Xxbw8A0GN+J83m52cULMUuoG
AOag0w9+BclLnwJ062pwIh/c9ThI0pxC9GDPHD7QzpBeGinBccTD9lxeVrNX0ZlI
Zn9Agv5vSFS6WXXuSeIUfU5zqDEu2hxdVTQd2Gnstih6K73g0Ql8rYdbBz4JQUA/
lA4anl4iuwaWk2uzdSJ5O+iBDiqaPdRZQoRL5oZGVQ/Q/fdKNOooAEqFQS+oqPwj
+TbS3zEbNagoe9N7HnLQua6G4uzUYYYp7sPb1x5NICGAez6SefRngPjpCgu/kI9C
FzzsTx97+DTy/2+Ig10L/UUHvZSnILAsMmXJatoxgVE/nHZPH+1n3x6I7jdOap07
Yfmeye1HtlpFxOnZ3+hNx993sVGodsxRUiDYl4sWKJ2OjYoYuCpUVbHZAhjR5jYA
ZN3kV3mT5+f/k4WocUu7VleCUw9pUd/c18+3k/1BiUh/UnC5AxXSgy9myaQmrPvn
iq1G7gg7yEMEBJ8wjOa2JRC8khavVE2rRSIfst/JQzR9+TF7pdkQYfpw19fb9Gzh
2H2KRqGdFnJP0AWxFHDiOiSgZ/nubUyBW2DWhBNtxRe4LJeH3pyUjrRmmWoRVyEM
mXupNelATwcnO0ATe4rjKh5+SGSyj3VuIsQFoaZlW8GgVT9pAReljEQOQOmBRvrR
PA/Rpp69ztyBh2kCte3faNKD0ZnbFZyow7CoyjX0+W6b5Bh9pZNWi5LM2DpfF1zx
q+JHxyS4ys046fHSRcan9zU5DrhIZ37TbUTnCih2l/ME1xwRYe4jJn0Gden5Zpum
fkOMOc4i2ditjh0SL73kQEgUUqEibEwSw1Fa7qdbr0eve0A/XrMOfUB2Gd2AvHyd
b4ce2LtRQhfpvmfsSDU2PGNCDskuj6QGZJFOnfxYlP5Ps4QU+x2PmoqD5B2Zpy5b
W24w589m80cR9AX/de6rLS9WJLPHq6swMcl89OZ+qUHcSt4i67N+ZS2YyjNihiQr
5foTuJ/Eqk6CN4XEGLoWJRFB1cyGMGKPIkQHUdiDVNXMnBLbuHvUGLOWVyioWWVF
MdqIv2WjGz4xikyt9Jvu5y5a4AdIgE+xlzKKRedr0GxNzWIWd2E0yO1Oxz/RF9RH
vylFDUw6rTz9PFmtD/ZmKvgblfhBemXUSKgjIyy1HpiFX8Pb2OS9GqjYMU5cjvfx
NnRjboXJc2ypOX4djbspi/wMVnx/8xmrv1+TLl7iwSfCLhLDyNnHBRRQs83clHXl
bI0Wch64SsN/5xBUheA4L0rrK8dq4HsewAp6RyMcfcNCPE75XiW3Gqrl5lTVDJ5Q
RiddY52EeMS8gTTV1AkKIvllTL44spBnuLfzDyBW/n4oOZhxkFPlwWKvBzMw5mZ1
CH62P4S4odmmOL4jXlWTB7xZXZXeMrLH2ulXvljzvgo6sfkyGnI0HzeGm82tk+bg
WpxOpGn/D0fSi8A+fT5X1bkr+ULtP/6LAf2cAkrz7Q5V/kQxwLCl5uSI235wFetV
jHFDqklcuzO+Y2I30zWh9Pqktgx8sW/uopSiMYt19LZzmtacC2bQSBiJUMFjDI/T
VFnoFpsjpV2DXRysA1rtQJdHvvjUcZsVpGxvC6mV3zx1Q/1+yxE+38oYyxlJUE7g
42igA3E2uukvCC66mIShBZEugNZhKRvjsTITYhdgDCgPCMKy40o98CHv0YYEc7DP
/m46ELcUYvHya1UQWnv0+Ky+ZDfkRTyn7sRY+1dqtp2wRknwjQf4MPsbI/KN14r3
rVP/u6JfP4zYldKwmuxSRE7YcPtFxuAga1CQTbFNxMKGU1A+1oMcNOiftRUxrqcY
b8CCkqxqDkvRPL4AYGM5z68z4pKHxB2pwCdo/ip8kSlmRPMNUViUdrwWNbtBjrXd
k9epcSgZBn8NmPJjX/1f+YEeHjay9fi8tdKhUFRUo4dyzM+qM2soNg02NjToPG3U
U7OhabDI7CU1r1LxtReBH1j03O8NHN7vg8ecnwVRFgV5YikRslTzQjR1asT4424h
hU0xa6LiNa5C6hQcbgWRWMJ5/dRbtNZdA+tG8YALknEZ2o3BSGdZ56rbGtlopn1u
4ttUw15GcMFwyLawDkRcevhZwB31EyJj32s5h4eIFkP6CTBTfumWBjjlA0PveaAy
TR68+whxy4BSvtVdITItgptxiKoIM63+/7B8S4vrnDAWrvNRf2RibVi3t/vbC9LJ
SBUbIPyEHWO4qvzYMEcBkbJTf/IJhet9o2xr9+Vk9zolMx7D7elMrB9hGCsJY5E9
/1Vy1D0SNozXolOvS5c1YAYAm5rFr9AshAEImp0B4H2iSsaAp6dVgjtFUgUMnFoG
S1h57LF3tUBWWc6Z1F4YaF8/qXht3O+XAU1D4df9ZlvZeA31tgXJSwHY/Nv9TlxM
+PALKh2aZ8HZb0fmMyT0tOQtvEpinyGfJBNS78WNl9dSDC7ARCTWHkb49rMmIbvw
Yz5apEEmaoHdsaAiRe7EYNdrhJ9qT6MDFf77hLDJaoB2PjrTXmH4YSLOlAgsBsKr
T/xmh2IfIgsT/4+VR620yISwkPb98RFFKHC7azJH1aBgJrJRMGiKVHQIYxNl+sbv
A34kaPT1e68maMs5x0rwuXzWLCmScj6e6tuXjcTelniMHf9dLtdCY7VAA9jKafxm
G2nNmrG0fbzYdFzztsUe9JdsapGqRwPf0XBg7Z0EHW9NA43JyVNuiKL6WptSPIEM
8FXo3w4hV1UNmSsPD7xgAgjk8gq2H2RASm7bNpCA8hXc8SUcV8K2XRvvy8EAypyd
t7BOllJdpwzB2W0IMkZtSVWYWFW/dgVEmgAyM85Pcpcesitw4xqNV46dnsLFh6sp
B3Epkzb7kUhmt2mxVvE7j4EaYB7W2M7w5sJalA3NQLHvc9gIP3sV5ifuAuIzkxK2
z1pJVT3pviAFEjC8NTAxUCv1ycQ9wAS8vWevSm3AK4TuiYhprc2NkBKZ07P4viXD
USH6LJiZC7yE38qUVRi+ZPhebHbq6YK4dCLzKZdrJrbMqPIH6w9LqPtlPc2O5VUi
AuqgUihcI7ChdS0F7UDrL4P49UVSaT6W2b3KmK5FRZj0N+VV5P6PhJKyzSXJYMHT
xYzeBls9Y15b76ADIGKD1x41jEWYcMlTRGg2u1PpmlwSKrAM3lKqFaLZb5VbxKIy
W6AUer3N46sI3Pq64xj5LEtVOoWBaLnjYgnSL6gqiOSV8uadN3QhSFtxhYg7L5R+
CQJRdJvx1ItwuohMAlV8rhqCVxxG9vPZLFklQctqsNYepR/3DaO/A+r/I+vEme1/
LAWo4c3SpWpb6qH7z4HGXV/VAnC522nOfkGvbKRUsm4Y+A0Cs5Vj45hi1UE6kthQ
TJphPlG2YTwZr8/9FKLja+6yQGtPhvDjPz3R7O+FSmB9ssVATLg8oS3a87SJGQ0V
BMyHeywWNCW04qNKGRfRlF2tMyyh2PB82RjZiN68R2f+GLksKnoNEBAFdhaJ3Ilh
mld33Nelo38NClHX3TBzAgZPTX01IRabOk2aMtt3ornHoMw0PmEb0/5GIS1ogzeR
y19JI3PAQBr7nK5WJEBXXrsRb5Yw7KvTcmqMPlCJsyoi7bMNNieIzMlgYLiOMnPV
RRHDNKNu/xter3CY24jCrAvR6N+znTvveSt3Dxsl9DOHaeofc8kJx7Ffw/2qjeaK
LgwmTlzEP1HDIR3ZLW4SQ0eC8JdA2Zxn0Jh7tv39YaqPNQex8sLcbHkhpaN5BE3G
nG7OmcIHQ5JSa1o9GLuFB07kh16uGJ64mn3AZU8+W4OCD1Y0ADQxFRzY4udva5RF
xKh0R5C4zVLPap5ZbDen9xvikT6VyPfVCcaT0OpBp7ryejl9Eznn7xd8ZM1zZ7Hi
mwXCKpWyg6t3OdOhCtlICwcgc3EhtuW/jsgqJmHcKZWAaNuF4o22OUOmrEvO+6/6
RqyTrQs+LpWjn54xOER3ny/9REmpXQsb+yF76aX0m5xsbGaf+YcWLlEY7Nj5cNxo
kKIuR37jKbvuhoxZwkFZB3a39Lr2uZ5znDcJBkSVdp7Hhj7/8cTYVXvaIWcoUoZB
gRKzVicBzxebiPfWDjh+otWias1XqxqzeWb2hvd/u1nXigYnRv+wMemZKzF/Qs3f
Le430RE/PtPN+gYpohyNqh07i76oKZ0Rd2sewcvba9zB3W7EAoV6AsyumK45F+s6
oY6dQ0ALQdmapQilTl0Kx4hJSFRpfH5YBAi+Z9PMgsBDGzHV7CjvfHtD8vmAHTxJ
k18OdGPIYaZmqijFKRinQwTnKYS1IOO92bvDMaNc8X2r3Wq34FdJN7q65Nz2rY9X
NWB6f58QudyGoKRYDB4hHsXK7HGA0NopJxqM1fMf0TeZWr8eZcFajrqMZX3XKO6v
tmUJpXwOh7PgZTrbRVPbykrbUrqv37Uqbls5UMvQSQVNXVWBTQDMSbyrgIeg2wGF
lmxQvcCQGDKTvbK2TpQ5ooN28Sh2//qBIT/KXoOD7/QOmRbWf56ktRneIoLxTCa4
ix5lnYlLCaJrfpAc7JGytW5La6BW3IHkKaTfVzQKLjuGDR+MaWDWK51sr+ZrCK79
68NY9pKTovKaEvFNqRZhVZF06JI5Nv8M45xFwq4ToxMvOWh0V9iaSiVNfCWWJ6Pk
FvYBbJce2PhkPiEnGk0YrGoV1F0+sS6O/t9pltTr08De2xJHfqbz7c6bX7/H762N
Q/mV50HA00Gk7j55Fq2NigMVMcSkD4uIHtyW3/O7ljLNR+d4In4FpOslmDjH8wj9
phf5mEu9RIRpEUXv5SWKNIc+hjFawREhpTdZrAuiyZRaM+AZ9itaabFiMsSeFu5i
br/aVK0F8g/PXTwJ8fKuH7OWPmzovvp0KzSS3CeZiuwfQ4USGOIyV9vBKYg2xFRq
RJIZD110bajEOaJ02nXdOKaA+EpvgmLHcuQ4Mi4GIvLapBXRNiWiRj2P0eKix9o4
ptt8N2X16pVK6a/5aG4nMiLQqdX75BnxkXCc0Mhf/X0re30odgDvL4aVpnNu6Dhm
7gFX2ipr3d23RRCc/+Mu7d62ILD1AXpmaAogsRz4tIHm1hWJanrnkPkWcredPPzp
BCHM8VLPXVGjM2jXv29GVDlK7WjXX2Gks9SooPYQfK7yDabYW6qBaLGUhuDwQvmI
k2xj1lqsSoDp52fdERa+zjcEpjAwIC9GK0RwVqGLnD66/2acRMb4nvbknYNmfNXe
v4aJqA8AvLUBP45X8+sjG+pSsP48v1TRt/9bcLOJlonrc4OWh1pu5vnLrnEXaTFf
3owe6usiG7gObUvj3vquzA1HABCxw6pJRqV00S88Y+468XyhI93rVi/0ng+Olt/B
hHj/naDoTx+RwRwZaYOW06mnAPWPbSnsk++094B6IXvWt5J1k8/L3zoK9i5VGO4w
4obqXejmmcF5FpUQrPBDnFx6MBfJbbcznwOAlKr3oU1j+CMEX0VhfAIgLIpIIPwC
VawxWgz/rH+m9zyyTfWQ29gCRrFuvADmoV017gurOjsI+L9+ELrD6m5if5dNKTk5
eZIEqjrYGMqEtQWNY14bYF6bct55m/NbF8paGc297obXA0a5BZlm6KM5c32Ws5o1
TIN+Pv4O+116H+PGXFv4M04vUcqaQwDUOTUexb8VDuSKsztK7dyd52YF7IejnOC4
+d2ScM3KPlPsd7ZN8O73FFHXWV46XQtiFK/gP9h02WctYUFQGYXYkjNvKqOM/yi1
2shoiUHI+i6KdZ/MMH/oWz2lcS6u/emteC1L63GX07EahjeLX8XuJZQzwxZdc/l1
6gNg5JptZvo6OcbnYiEJPKe6Cf7Hk8x3QqGj3Q1ZMT9sSfM8ISInPujEYmcJva8j
6ZNz+QtcL0NLPtxTZ/JUx5lUYRDBmuLxBKXG7Zl0JF+3FlvXAzlozAN+BdRCR5uL
N6Z6uHpKLZGNtMhfW2NpMd0sPauFW00u+QtusofM6spROHsrtKNmQJ5VbzpLEWan
tbXdX5sdf4wVKsJM9kDM5xgsv2vNJ0WiY6RFxAORUBCU3ALrygO8NpKg7/zAfoQp
/p7J9dtoVViwNsr9ppH2UisW0K4Iwnb0UclUAF09JEHIaGZFpcM7h4QE2a+LsEKz
9AHxOypGJ0rqOJGgdftJ/9+juxG66EhXCRcP6UsoMOmHvWayUcejVJTyjDqP1ckb
TZYBu+ff23jDQsL5wCVjiJJbx/VH4whSg2QQfA4xZNzyk+RZgCAHNNBMVEOBaHh7
i6cCeN9gCWsXU4wLrYQoLkiKkjO+N2Tw40u4SijpHgM6XTgwGLRwn1K2n/F8xw4Q
6Fle3MrhFKPlGxmAFwxO5b0cZK+MgyKF10mUEfAGDB29cxKcQIgA/ot+8rCoirG8
8/fp5L3WtOYpgY+YnU014wz16S5X23S0DDGNlpcEx8ksN7bUaGIxhQZcPj+7Pkse
/gVqV65pUDZq+HnvrNtpJAbX2syB5iFWPpJzY/IfovH150zuPA16MMK3LP3ARNXc
x3oOGW7IPfH/G/mFS0W9yZB1guW/hfLJWFvnFp0kC+bIcCTDDAFOq98EE2xr3ANN
cNqMMPguCzkykxLzvDHSaQX4JWGtVFeykwQQr22/QFnIrB7XJ9ApZ9LssINdol/z
Vg01m7XsgYyY8RoInle6LfIgJTk1xRtRC+4+mzphrp1gLkxgoUqGnfaLvU6+/QVo
MdtZNwHkPHU0HRlhP62pV5RD0me0vnnDSxY0wYJ07dxhK7bYwGJ6dJPhZQ6vbbJ1
YRXfWxS4+XyJNxcT8u8Mf0iuVrL3jT4IDQCFR60O0lwxud71JaGiYICjVgRyc3TF
/OepvQPvnPu8/6Ed6VuY+fAlKV7IiMEVOAVWPQW7V4DqHo+EZd1KAskbkYepAhhH
28f/bsZpgt62oH/mcpHPbDC/vM++dgkpB2KUA399vh5hz9RCQEvjKmRLrDaLV1Qb
U2THOqVMyQxVchskM/nh0attHrVl6xzjRn1E6bmEKe9nrY5BGToIaisePd8ju0SS
YkfBssOWWToPqIlWW5YBFtx8LK4Sryk5Gvm2d6c61Rs8bsvOoau2I/2bqrBiq5LK
Dw2siJchZPH5zcN8QJhKtktve673p9b9kBfJ34+HWR7GDIsn5bUhYO3iAqvlstcg
w+VYPu1WIqraaWoALhkeXKu5wbd0/mELWVfNwF/jhz49doQWAQL25ulJcYkIKVHZ
gP+1BCLYmgIgyxfvlKz8FnVnuenyjXREBT7peUCImaZD6tN6jTlC7xR6QEmVOWHO
pIdr4Qau/6wJ47Wmx/BUUHeDgSYrdLCSAa2s01IianB7T1yh5OvgHagOpmMVc3tO
yqObCp/SSHz2EkVwa0jN03dqr19VsxXgTTcG9+0300Lf1/dpluI+1TTveKc0XWB6
5OEep5K0yc+ic4DHS4s9IyD6m0B3CHi5YS3Q5WBs0VrXMCsDGVQoPlCQh76HLxsJ
BJmXpPoDl/BSrek1/057p/Ct4a4roDK7QVTdm4s4owPJQ68FfLqAafLnlTVd/cBe
qmxw4CJ2v6HNQnxb/ZKNlIT3zMI+9l9G8jenXK1pskxfmWUfabBDFXFkFsG424Xs
TuScxuJC5pTOHCWTqIBsSKRrn6NfPv/a8lAuc/145yT9dvLGFsu1FEfRC7MP/44W
kKjPUnog7/J/lnLt9yrp9BFfeXwTyhgUpg1Xpl6Al7o7ppM+ZyWHznLDuvIr2RDg
yHitpECD3ZUo8R48BC2nWlJFhluXLE3QPfa2E0bOn+YPOMr1XLvmbZyh2pv14cKl
5UV8yDUsAe0ZsKwme5DYi8bNkV73HuIxQhlC8CXc+eh/lCd6oqv4C0IPFO2IZPtT
dvdOiz6LacSLf6L7ut3OnD36s0vyPKkvpvneglw8GTIMj1QQVOr654gxQKJRjrkZ
KRTd8HyrmPf/gkGg7t48TT9v3mqsx/Tb8LBMKDwqiUtPyvZ3Nr8/PGHPRQcC5TEM
4ON4IL1sxdHmRtWV+JO/oY5wkEr/qA7rN6Sl0TsadmQYG9Jx1tW2vNRVdP+/QEtq
jsEIDE4IcVJFDkW0Z1t+DfiWK1PyjIJfe6iM3AoyObIqMV4nkUW/nV6b01mXmrlZ
9pOLU7MiAxP94Q1nnc6viSgHxV6UrXZO6rUfKz2nO3FSd4YiU4O2ctQYsOpeq+vp
tYHJtU08npd3O7w18GPFds6qUfl0AK9CqH5ZePnZh7Ja9DYLWjP1crFUMSN9Xtg9
yEUNkVOW5AsRIjatH93hekorS1EHDZ8Tb9cbW+tc7OEW1Hw2pLg76sKqYeo5SrJo
jKO/Yk/dTxWDK+p70qQ+5M1cpNgGjnDT16QYBgHTyOF2/bmsJYLMWMglpiwUtqSc
w+uLJTlQYg8jZ2GV9oryCGk2spN3Ka2o+TMq4Z+jxB9+aBrpYsTgYed2mO5IyyRI
AUMysaHIdIT31ZhRzXpxCykcrKjdPjKMIKrRSjoemjqEzDmr2j0jD38Ur8I9P6AS
x1M4wlf29uzUeNPOA2WSe3KNS8dnXztiCcDJrd2CyH/a2dpxnrbBaWmwdbpoydTV
tFowu5KZuNpl7uGDSwXLHQZuWpUgV9XYPG6aG05w3xNDKBExlj8dyOEIusHrb6Mq
nPQc6VLHv8UE0dhVqOtKEMm2yXQAg9UTACTMaMTuYFvwkgxRukYHJslLoTCPiTOd
ksTMmEWI+gRyyTMVTJ4l3kwEqZOkKyTXlZMgvC4g+bZNgrieXrtO25owxJFx0Dg3
27uXFoxU/mlEb4ooc/WmwgMTRt16fAYREnY0yzjRa227haGw5plRPWJMJJv3Uqjg
wTMKxYdPBpYb/9BswOXL4HDFl1jkgAz0XNAXJXNJ9VE+vz0P1iLIFz4NITYUXXcG
gzg1J8CFI7Fe5noPejxh66HP7B9ogOcAIlbS6d8gw8eidXZWQ9AxSnFIckNYYtT/
UwU088sxAS+UGaLComVxLO5B3ZanNCzTn/n6Ja8jNT8GbY+8ZH/ovBdQwCJhhWei
KtYwFkFrxzNQYsvCQ4hAwc4J93MWjnyjft8LwqCInp69HVP/uobfrjk5atj8PDJG
Ei6IBqj8ulH+qhPCNcwpJZxS5REMQVvVDrCB6r1IR/fs0swMQ2RjKx18Fj8GxlAW
6xqZoKj8LhpBAFxp7n/HhKpuJNjdOGsvTH/Iv72byLUPCoqrL9UBLiKR3zOJMIqz
1EGZwRlecZWqGm1fR2mCts7DKUgQQkBy05bHIfSaBYgtrnkTzIEJKd65sj2vJvZv
LctbtudEHtbGEZbPf3z30dlmfBqccvvKhjuahGv0WdH6B+OvTzbJyMnmkx9uYFeB
Gf8/4wEjTbpQMeZAWJJuiThHCrgBygaAxEilGYaiZ6+SUoeTiGAAxkBZcxEyU2Fu
v+cVuHbK1c64kdWQ8P4/6xmUq3TbhhVU8Rx6mIDmuaMEFr97zgRNQs4HJf1pZJlH
B4OMqnEB8RpWW/7E5dut7GA8s4lXSHzrHUskdvdPSXcAh9OR6CTHQX4G0nP9JcZW
8GFW/NSo+fw5oE56xjiFiE8J69HlnGBhidMdf9CCBTNTTejzgZXkYwqmdPaN5VNg
HQ9olfoOq9/ZPwTb27nmB+cxCRuuRCFTwHtB9oUvWA94V6MxOU0y7hXrbVoW2AZK
drAspoy2aJwb9RoOI4a26ArSXk2g1+rz7X2ZUsqPWIaxgEeG4PsC+qMO4y8zRpSR
OsYroXmOSpJCV+RZ96UfimdyOhdtAJ1SJJI9Fqu3Gcpcv6/xGZ2niAFYGqWwIAwQ
UerAIaPBQ30aQNZeqyIcXViasJlDffK45cH8LvDzQvgwh38mZmVdH5AgpH09nyL6
AMhNDMT0X7wZiqRX+BZCVfVX/OV+G+iwZrzA69mv32UxByrzFrQxLx0yrwxN7Vvs
3tTpF8ES/j1tXODfe7ne6EeSDuF3xA+6n+rtwvDWR6lVVikwphVhNEGNVy0xHhQM
OobV+bYZKLRcYAKhLGdQvciXxQqwwtCo0j1qchb7Lun0pM33mHoajDnwzg38OBZj
vnD7MD19LochSu4KpcprKCtUrsspMyX0aoNbhlHzT5RXtGymmF+KsoWY1iHRrHbS
yUQ3brqoFSEpng+cVWvrxHLnayv3FOesvUsfPzQxfyJpRuhcnQ5s6ZXePbHfoJ0z
Me9oLryb/NSeFRZQHeOzvS7Fh2rzj08maG3Otrz5FvBN1sAw9ISH65dhM159nuNB
`pragma protect end_protected
