// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:28 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DJADmh+zvXC63r3cEkf7IMT/81ZocKkM68LU3+ybdEJ0qv+Pl96kb8gRKc2sHl2G
hX6e7elSAl4S3fk46XjCxvXITKpmFzoHNWsIEgANwflclh1ns7kwG03qJeYo5rwl
lQa1vuwgY8bsL/F+grp1QY9pl20pGkG70zXcRX9ZEU8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5568)
TepDYqhvpgbMjhQob7oDuE1twP90owefP/pvFiovJM+MWrCI/bbO3voP+LmfEAId
yngTQWiX+63Yaa1kbMp69ZOcPcoVYrnlfKjdjYiIgixmLAHD+uWB+jGFj/M6Mat7
UJxImqVEb/Ao0/KJT97STx38ZrG5PhZoF3v6L+eMY1djEYnFoN4mIV1N/2mzQOV2
qCdTC0Iccl/RsRZclRCo2uYolMwRU0laDntScPuYM0iR0PWi/KZR8XHXHeYsYDqR
nJQM90PZTMXxtrY4Gqfw1KbGxJE6kv6klYPxv6/OqafQkOzNFiJDy9tOfgiXDr+K
y2M0LZE0fjLaLFPLJexiPWuY2vneCtqkPARI0DFCXspw9iYn9TMym8xmv2J3FVzV
fQde+4xwqMn2KUOqSWZsKQgVm+AxzDPQpVnciCk1OZz8FI43eKBG0zM3gCR34Upp
z5X30R8lf/tFNCOITRrLlWJPIu3dCOeyjaM/c7jAIgXrBqViiX4d0wNd/0Dstb7X
Rz4Y735eF2xS7/ghPTvS6aqN+A/9IB+U39blsdpm5/8yXjzT8uJCz16H1vUa/Gms
2o0Yb2GQYhcQ5t5TG5eFfJKDA5oDvF1ZBYiPA1e1jIN7uWqrMxyHN3jbyqInEOu1
c8Vvlbg/gfKecmjVgsnhRIhsW/KaspYAYGmCfPVnQ0EQEju5vxE9t0cut1Ls+XuD
8YzOnilC0C3wn4ElkUBMx3BZ7YoX3DcvvrF6w6iQQJYh3Vz02VBJZsjD2wlU7rFG
DEndZ6Twl6seInWlg6S7bi7s1c77Ha/3Wt2JMfx75CEqD/PEoGBYXYPxQbT7fuxx
AV2H1YSpzuVAcSILXlAhBB0kE/YSQBR1mNoc+BrUrpmOQTYeIdJ69XbM788uAfgm
9/GjHf1ADrZWBQygbkFQuQ3Nws5C3/Jjd/RFXEEDNSl52woPGZ2b48QeDdc4tfs5
g5JVWxhCypxHlZEtrPb2cmNLgfwJEhRz/HhtTKMHbXufUnZ4oNP90pJtG5UVpuR7
yucSdubsrbp4z4V0V4qny/VkIrD1gmuhS20yRw+LlbGL626raNh9UJ/yo1kOUfN+
E6B1YFaSifsTo3zmkWnpt0fjfQeB4GB02eEDASi2ZBXp6lysLs7TvwTiqj7389j0
00rZcBnrx9R9F8RNRlUFjy2PcM4y4YdVdqERwmKsxE84HpxIh9QqWcug+SeRnHvR
gBV+yGV0123V44Cf39CZ7IgSwNDmGE07hEH4h373XglRXvjyEt7pO9orRSnxJVmt
sUsNouKKsKziCVVKwEYUPneO6iNfwEzPXdgqQK7lwmpksrHBVEaQ6jX/nFPj/ROQ
SOjuBDN62BVN40s4ztVXTB8ZJ5nyNIwIGbA3+o3LoUjj+x2gqUoF6wxmcHJlXViT
kuRc/dry27y/hqtc//naYn35xeucYz7ZGABHaw8tkLgHo7J7ZFt+HUOeKsm6rl3i
EiLtIu+Da5lwlYMhFQPTUYNBpMLn34PBePc+tQiTWBUFTw5lnDgyJxrQAQRHryAA
qj2k9C2lwPTRSqFIpxzuXSmJGSQO38dbnmkYmcHHI9rTgcLQG7M9fcFr4EkAX38S
aCxEFTkS8eikgsj6KDY1AnxzvrdFGEbTQrYNMrzeWN+kyWTZsXvorCxda/qjZHqS
8PqZl4FCVfMe6QJT1LpUS6z5qI1R2T8b9MFdhdproRp3g5kQ9aPL9YqAWfKtuM+n
lM9l+TrUPxGFR/7dvpofrR06EFnfvq8KYamXa7QakUIKEL5cfadw+hVVqw3ceQAc
aomypQdwhVk84tPlrxw5oSQKtTq53YBbYiux6VGJPIlyUsLL9IRvVr42oclXv3eY
rxxKMxtfINmihYcho+NYv3IHIVIEk69wjfXULYCoADOKdwo7zTYTEQ9R+pZNyAkO
TbrvpbDggoXtGr+03sLw6S8eV96/YG8QzvBTTiKKMpqc73tCzlwOXU6Qpvlc8gvp
8sFuzB+CXQ2nvRMqYengGko3N0tiKrSVbu0rXicB+x/nCZJXgt9zH5XBdFMvwuq+
KYBpuUg9Alaycs1gHzMperNnN+FLSumRccFJoTIO2bR8TRXW6GAvJhYvXXMMHoM5
KJMZfYtdKH2PLFqzF2GpgsD+j89KZIpowVJkS+hED1hQzGJashfYyZYm5pgYmkin
p4c/WU+TgBHRmLXryLedWTvzC0ab/6rc2rTcKbCrDdRdPID/WnSPYkOyqHT6QV42
tbbrRSzFc7C7kQ0G8swmE+BrTlDbbBHGC/l/hnW987Y4mCxV6UCPnB5/oVXC5dHD
gNUM8Ao3k7Ep2o20Xa9LVM27tFVW53zFt+8SdqS2Sx/2imHkAU6xVLR+kcDUzeMS
q/siZ2aEZ5KwKsJ+moKjexdah9/nHv5tBqjLYi/sU23Ns5KF1Q5iH23hMf8JHtZ6
30ezckIsyNVdZE3en9AWN5WPJ8JsmCtOtOvhSP1eKWvVeesgXjxwGzuQ3B9LEKCo
UDHWebKTD2b6wMZ2FN4QqnQH5Vm+a7/brDOa3emZGnUUQMz+ro1RVt41YKVpADs2
GJ8X3WBcFWrW99aZIjRFF9Yo5IMSSMpWbAYmiIj5fC8mtpPlrxODtK4IXFAv2WXy
4KcGSLLOEfQy+wf0p4GvWiN7eCbZNLmVe6BYXTtcoItN6nhjm2fuRuPusa1zTE7F
1+gYyUNjGV8EQyj5QmIvCmX3E4YnYWl4g+9G3lxBwfgTJ6t8vYFi5Gs3x67hDAui
9f887WCwWHBO+Ll/bTLNfYkuDLnQ6EBm1Z33ikGBKAmwbs74bqdrsjJNmmiL+WlV
Zo/7/GQkjmbFZ9E9NxE28UHqSPfHtVuCPS0T8fZL/vI4kPYgHTEMX5MZF4iAR9VV
R3jMook40EYk1ffa3wq6F9pn6wDqDryumDK1duHViQ8wojstk1uzyR/fhgN/i20l
/YpKqd15BSQuan6V2hSFNH6TYwZUniLi8R6quomWiRSH8gvW34JJhdu+ZjFPUMb1
NuTte+ztw8KiCEawBxDLaHi+oC9oY8RuAbro6FogL5eIdKRi+rpPC4X8Ln+JRYWT
On1H7Uw//PoaEaiYIJrToT5emJwBDcS6Cbd+j/ND/9cZmGd4emJVjx1l0so+WWwD
2FuN2HLgObTOaSgX1SvPqU4KjmjlGZnuoCvCD1O8wHsA/10doAZc5D2lwy5BcA4g
VKa+/Y+32TPBuZSzuLztiZN8OWaubbbPfiXOqhpHot5jM6zIut+IuMUDTDtRzscC
qmYZhH+U/RoPMYf0qA4wtGdFsKFGpdIcfVs5cdR6pIpYYtXUZ7hElIfOJYBk00kX
0wLefbUJac6M14ZWpR/m/Npjy2CGfdHPN36QCDu+J2fZj43g5poGvet3MN73TZFb
61rHOHjP7mtJZGXPTN67CW44SEWbPE6T8tawzrO1JLROUnhc6aKxTJK/PS2i2KPm
UJSnO0t46kT/7h9P9w9KGqSCOllYTDYzKK0VizwaOUwf23cQF2l1FrE3UwAMvnei
R2xU5G7Tw+3Iwg8EbrOv0sEmTeCbR99mKcf0707fqt9xNn0k2IvKDBMnN0JJLAMn
Ix8ouHRtPOwH1Xseq/IB6GR6gjhKnEvgV+AqAli1tciyVM16Jt6+lqntl6xsvNps
SQrm5GP3xiayMgQeGBTM4AIEzMQQ+Vm37Qte1EpB2OcgojpLbGxDI+ESs6ZbTmED
MlQ5DrxmxoS8l8uQkQFHAAWnkGTbx6Rx+X6IlWRq1QoQrkv+hKXng2s1nGAc4euZ
NOFOYnh7xmDsSGdpk2RAYLMgNqLOwXJc/msjfpwkHhu5GPBm/gwrPdUWcEB+k/5a
GcVsinn2hem/uVoGqUsy5tGdtudEXPuwmaTGagK9OfJ9UWvz08seesbuK3z61wPz
XSyMTKBwcTlIFRQ/Isikn+1e0hv+tuEvbUNPmchp824UjhFWOac5aFfi/EJHkyEy
p4zv2C83uGA/gN8nU7hkySx11SXxgNJQOu1nGkOT2w5wJHF+bylNTUqMTZmBIkg9
rdFpB/Y190qSvlTJFM1kUncjXqMOSrXT8jNJGjX1FsLvbe6RvwHuXQdmrJnCuTJS
7ePAKOaFeCS1zTLqGOWVbCKtcPbOjEfMMpjfH5E6WKZW/sclpJJtDToSEmf5zfum
W5jLfXwu1kjscuXU2UblDuNQqvfEg9aCxyxuxgaTAe3oEIf77WYE6EVwH+L8gJFl
SoGlZKlU11zr9ljntI5I2vY+X6FqCQJpanI44hlWlu8gBldf/YOIkF3L5qEdQRyH
FOZjlx9jxezmViaf/ll+7D/rS+lxn2/3qqav27QPIh84EzWTqLthbGYBgRkIsyz8
OTGQuv8AgKCWJAnAYZkr3HtZGxPm1ejUfznsG9ac8QbNTdrcBf/Z14pKzrZfShh8
bmpse8ng1vZcPw08qv09e/c4JtxPKHVSvGRE48ijUpMx5YfvZeLhW8Ytm6oBmJNN
UbVqolW2/Vv7dKhN+bwWFS/sGTYHh59UymCihPLAw0wQ6O0dV5IIDXahu/yxd3Vc
AKu7ziavbFW/R9IUEIbnifB2WxCw9a6nAWPorGcDuAGeVo3ndTO40+AGrhHUAkFc
igs3VQ+YuZiGYJL0pK+KJHoPo7T248HHtuIWXK19jAWsDlfWMvS5zHaO/WfGKaVF
E+F+AjBZfGTbjplsj1YJqAha6qgDi5jU1ruMh7PV2bfkTLXsHkviJdlghC/IQeMr
AbprD2VT3kJ5DTOfqg6o3QDifDAWSum1ULE6QPVAq/z1xP8sWcCCBCaryIYN91AJ
HBG/7H7Sb0Kyrd3nDDoE3sopLqHH+qUScgZN78WXhIIjvCX68x8lj1w8xCAfBtrb
hsiARPeLM4IYuXrQESCgH+yZlQ1SAVSEJWrI5HPPnW3P1b+0MVu1Cdga/Ch3rEz+
jkCKMdieWWZ2n6Y9GuJ2XbBEDv43YBxOMpuG6KwKxvCurYrtTJqjwwvsYqO2igLL
94x8xE10RmhkYst+W3n4dXwwnWHATQOsPP12GeFtpqi58r0rJfkXtmG4PBn+NUDz
Mge9ey2/HK/5k/+DtUEqdPiTQIH7A17vNscTdmDul44JBTpth0u6yjPq4aAhjPwM
iTauzs3w1ZBBveAEr3LiKZDTpt0I51zGtqqMv1F+khTSUPHPg+PCtC7+nykMFW3B
cmyFPEOnM1AQOtjBEbOe68dx2XrMqs1zaw1/9e94TksJajwoxAU3ujqMslLiZwx2
25A8Ldc0RZ/w8UP+dSh49vABebSa5YLqya7WLDtyc6LuxYCoM5ohVwzP1XJeJHFR
XzZFc/QhFOO2UTnsChvpHlXsdigd2DJ6A9czWxA2v/TjV/nOvVQazBjpVF+f6zyn
cmLJzTy2jOgBRx1F++Sy/GvQuRjMCld4CXrAhF28djSWoqbeBLZs8a8+PUEyY+tR
lnACYeD2vAk0mKkP62E/0DPqnkfslNrwODUx97lXMZ0ulTXHR1byt00a6L3/6jID
TwE/PmlUCFlF9Y/GMvp+k2jGBouqv6RbK6lSAociEIn2/qtfcuAMR1BMeOHu6uyg
1lX/TInFu67hqZtkuwMObdkw6Oyc3/t4NzDgI2Ffplj9GFxtZ5+W4z6SV+6Bdiqq
KisOWyE9cFWMLJZNiFMCVbP0mqUj7cSPOvfQuNqipTarNyP2b+dXQpSIpoGkGbp3
4aP3DDiZv2NpNdD+ClHo/h2j8f7og4aEscFu9BbWW/Vl9Yw0P6pnwgCXd4JpbLg7
bGAdC7Y5J0f8f2QeWH9MLPNNxwnMYsCnH3xhm1fwQ5ctrp791eDphihP2ZAaM5ZF
Z3r5qGY0CnmcgebOVtFw8TAn70mo6jGChzb1CFC+UIhgWMmmSvzc78d9PZclBHij
gfuvVjiOy+1n1awnU0119/2+NqBud4JFjLdGA8l3UBPW8U7fuaY9Ieg4dQPOBgJN
fc01pUkbSg+VGmmIhaq+xbvHNLOURuWK+AabcAqZk22QkA1h08OWQtJgrxffRjn6
ywKQ+3YRIYwzP1YZF5Fyxrm0JWLlJ0xyg6VG0KwlQX//X0rPebmbL7+Ud8O9NoxM
InFNyY8xxkwffmvg0NFKTa/BJ7sGlR3PGbz9l98x1jftlOwqqUaBOj+FhRD3BiDp
Xq3cXvQTzxIxnSyiRNuB4pKDRu3a4gb9ZbvCiXCJMFRbcMsUhDgH1f34bB/2g0tO
eYV1s2TMm4o2jlTmOtk26Y8+mDMkwCV7hZI+WnI78O5XeaPv16OMZYjcuz+25ROP
hKayVwI1BywYj1c9uj6Qidt7h9cLfc/fLJgRaxjJ+M09ydsWSoNa48Hq07N0fVVZ
jLSWv/15h4+oDrs1t7datn3uUBK2fAzS/NgyQHBnOFk9Y6QR7Hszox8d+Z/Cs/1f
FUfhkJtUSunJUv0AlOih2ka3u8eMePcekIwHkklUUXTYrhusa+JB9FEXlQQRRQmn
hy4w53kWr4IPYe0dhrKFH5z/ADcBc4eSqlkzcDFgLU/7EnxE0IjuIyQbiQx5Hdy5
EcEqeGLv8Jo9lTDH5tHI2ybxn/hOFK+YgQnj+k+pPiCyPzQoXrTPgf4QKsc8YjuV
UUPVOMy3a55oRCd6U/ecKzJmNvgSA/JwEZyl+AGZ/qAn2gPA6PZGmI457oGYooDX
yPi1WGjr6nXNqg1p0pPTypcFXhvmJUy4iMFDSgvazCKuHfnKhtBuvM+WNjdJYcvN
Sg3i6wcT9GkSe1WSUw5+33Zdd6a8kEq/sLnJtSVDYWAEL86Y3nfs+QMPVSHJiJ7d
NhzgMYAOYSTmUviiY6Rk4gJwWLVc1v3fV8mvRHPGePbJQIXcxAvf+kJ+dKgMAFpo
xaxo+BJxUDoOfhQEUXYzgbGEayVj69THhjJC+uwpctVHecOUDgwybq6ywQMoB02F
y5BLoGX1aw3WGFMBeVXTvHYY7A77ugFcZq2aLH2/fQAArs2faDnj5xiMXJvGr73u
YDnK/nYB1yiNUOG1+zgnfIjrw0C3gW2pmN315A6JehqftZAaAtRxpgtD4YDBqwLM
5AanzVXYYX74BXPjzS9rKnb94xze7x+ncpfYmOuk3BBTxLrESR9/VnNIGkH32H2M
GJaobHQy2vJ1QNOBhHuslypVDyZ1cumb85/oyjb/83dKV8jYEaRFZIQFMeWtUNVe
gr807DyAPwXQ8pFZCDHfenqPKmZWTH0KF5xKTpSb92MudGxgButqLbDDfE/0swKD
yNQ9OOlu2fDpcKUlrygmpGQKiPvW31lq+QbzRGNvPsm+ofN0oqDZG6LbSOQ0mILL
OFXPOIuDh0X/PmqIGVJj9alKHuV5GJrMhUt5Lv7ogpIMKsmQaK+DtiQqbUwZFfRs
uR8/7hh4Um1afp7TY64MkrDDnD463rsCKoAYVUIqY40t5UdgfaZz8NBxQ32Wjahn
`pragma protect end_protected
