-- CICU.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity CICU is
	port (
		in_error  : in  std_logic_vector(1 downto 0)  := (others => '0'); --  av_st_in.error
		in_valid  : in  std_logic                     := '0';             --          .valid
		in_ready  : out std_logic;                                        --          .ready
		in_data   : in  std_logic_vector(7 downto 0)  := (others => '0'); --          .in_data
		out_data  : out std_logic_vector(17 downto 0);                    -- av_st_out.out_data
		out_error : out std_logic_vector(1 downto 0);                     --          .error
		out_valid : out std_logic;                                        --          .valid
		out_ready : in  std_logic                     := '0';             --          .ready
		clk       : in  std_logic                     := '0';             --     clock.clk
		reset_n   : in  std_logic                     := '0'              --     reset.reset_n
	);
end entity CICU;

architecture rtl of CICU is
	component CICU_cic_ii_0 is
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset_n   : in  std_logic                     := 'X';             -- reset_n
			in_error  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			in_valid  : in  std_logic                     := 'X';             -- valid
			in_ready  : out std_logic;                                        -- ready
			in_data   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- in_data
			out_data  : out std_logic_vector(17 downto 0);                    -- out_data
			out_error : out std_logic_vector(1 downto 0);                     -- error
			out_valid : out std_logic;                                        -- valid
			out_ready : in  std_logic                     := 'X';             -- ready
			clken     : in  std_logic                     := 'X'              -- clken
		);
	end component CICU_cic_ii_0;

begin

	cic_ii_0 : component CICU_cic_ii_0
		port map (
			clk       => clk,       --     clock.clk
			reset_n   => reset_n,   --     reset.reset_n
			in_error  => in_error,  --  av_st_in.error
			in_valid  => in_valid,  --          .valid
			in_ready  => in_ready,  --          .ready
			in_data   => in_data,   --          .in_data
			out_data  => out_data,  -- av_st_out.out_data
			out_error => out_error, --          .error
			out_valid => out_valid, --          .valid
			out_ready => out_ready, --          .ready
			clken     => '1'        -- (terminated)
		);

end architecture rtl; -- of CICU
