// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:46 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Txm1XmwtdHnQWYot3FE4ypt54WDAMs3I+an+6N9XnkuDTahT/nt6sEV9Im0FGRWy
B7HutK0NhB6+PTbbkP49M3Zl6jE+sb7KSGX9g/3eKz/NLtxRMCsEgmdjUf6ln3yV
In4EGuPeMSStC0TxfNdTvXHzUBBmAw9QlaOP4U254nM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
heanGWvjtWdMi4AEG5DS6XIWvs36swdiH6gH6bg494aVTlhOJlQym+swFEei3rsH
zAC6wiDDtJGi6KUvadUYegHeVaWQOAtPsYwOczdevw68y5bUo1kA7nDs4xX99aoF
vxydtli8ckuEvaLjjF7OO0PRitE6Pc9Hhr3R1f4+vNoqjD8AH3HMhur0tGb/gkVh
qRjE0Ur3TpZGjxI+lnfVgkgShzcrEAvGa1S8u8rTJ+jOR6EC03VrqKD9NRcSKsLX
TP8jME6P4r10zBx7UOuC5mublCG1JT39EzHjGIk/adm29QsHWcXgKDMptN5HjIQk
Yy7ytkE8BiG82Qr4Z3fffNgRi9GO/X3egro9pv9983atqoi+bNf4c9vOyyx+IWE6
WfOBY8kM6lXiYr/XKER+Gsek4eG/1ZxW/LinzXaRrQw4sR0oI7gB2yOnPWgWS0Pf
Kh+j5Yn4b3kFMtxQuBxyYNl4OzbdMdbKFjjkyzT62C9uvm0SqZqyJ0pK/ODmCBOE
kLACu6pvV5j63XTqiNHWEaJ7D0z22Qw4NwERY7noHMDXp7KWHwSaUVRQMLvc5gO1
gYNg1fjkeilC1zKJBAxBGCdlg3Al5LJ9K8H/wO1YdKTxK9mCDjMF14lP7hsXIbez
tw7HKtD8ToDODaAzWyFPfvtrKVwdyyUD07tYL3wymu2ntaX5xjHaJjCnM51GVeDo
TVepGJsBOm7i5pb2wcY1oYrj5myqNxDV6icbrj+mfPrghs1jf2ljjV+CdX4x06+l
KXHp5epWT50iXv8crlHxIzlttiTsW6Dt2hPBnviKdLfvzolMJHHR196rmhqkXoyB
PfAxRGanLBt7P5g2KFFFOGlbWGf9ojx10ggO+HNQUpFTtdiQQORES3IoAL9xakUT
46yhSB/9DI4z/O+3ovghPuU3qt0fLPL7D1OYbj/G+F9lT9yMM1mJ1bd20CLv8xkx
/C4LFW0Px3SFXbmgPOzN0Cz+/QThg/by/9AaaPrz/fvoHtup7kBDkYjoDAChEp1B
hmjcdLewDE6qKVkg1/Od64naYht+I9dkcfivsT6efK2muH27pgr1t6wvkz++TFuh
BRjH7DQ+8GtgFk8/t99RozPFAAHTd2AtZn6f6rBQxInLa4AfXbRZW1cnEKInGzqT
N/hG+wgS/9tBEi+ghgQUuwrMl8lGr3GQbogLUgjPdD9Uo1Rp6EO7n59GstzhVwth
5DeP20+9c5iiX4YNVGH/mH/vDGoi//sZ1AiEmFHEOPUtTbspJSqzu0eNfn2L44F6
QoPTiobH1lHMKCQDUFmg/IuzH+/SxmPdxlAMVs7LdNeSMrQpWN9XT4mYhS43JBWy
Svo5oIC3CfUxPOuGz+bW67hpnRmTGMuQwIZTqLaxoRBx7DdPSWPbjbfXOdXfUz2l
yp2okm5tpq+uq+hyJvJdZLx5kbl2cW12+8C3DymNh0xhpgpUHZtKYm6st7L0Obq7
n0FaADXSm/W0RRrbrBUp+ixuAmMKbYd3SwCTubV5Vj52o/PzXE66j98Ht7xkZ0WP
s8shq6cLFpyn8QDk3dk91tOonB9rYiX96MpcMDwgSm6G2caI0GoPnnzcNgcgboTj
/7NhTKehms87AYa3P7pdmF1xHVNUdWnjYLgiQQuFncfQ1wYE8fb55pEy2CVyQxnA
hsPEgn7HDQh7/J/Do37F2T/vdJUqruIxp0FElDdkY/yutMBk6Vy5cfyVyH471jY7
WrgRLhI8uiPT0M0al69rZqFvUbuWBXwwrsAj6GEzRADkaJRdYSs6y69FCZQ0ubrt
FzNYLeKLVSBcW+8SH6Vb+7f7/q/u/nGh32Wujt8BE6w8s6bYJkKVoJWX+UN9Add1
VY21CrY16IjiDSRqGL2loMT7gsOq38Ym2jZpKs8ZhuRnt6axpposDQ0aRkP42TmZ
1JqXc4EGjBdD3MSbGlYQeTaNWqZTD38+zFLcgYkkyzWXkkb9U5Q/6bDfKiptTEt0
0zTid0lD+tSSZlwYZDDBGjYE63Ihe3QGRzsQtDtREAeULkXZRI4Pl2IHeTTd5FlH
2iflBy5sUq2beK+qtNm6GIHD0tG9ragYL+1PVPAkTq10v7h/MsUSxU57WIaKQxPa
QuN29HmPWaifjYCcqNEp9jV/p6bKmbxBQy4LDQmNaWF8qjxUA+vm99yyRdEQHTMm
1k6AYSGyYAMejq84AzubnTUhS7C7zSeVE6VUI7ps8XhIX72fB0kAdz91av8yZYVM
m9w2yVNynay8J/7YxcsuYqEzohwoU47pb409Lhip7UA/qD5Br+0urK9AzZdmUZzo
TaPW3MR6jxK8es9W+SVfIWER5thGwxaqY2/uG6v2DEaOU75DEBOE1HaCvs3Wiajh
5YVPJ5d8VO+vwr2UBq3HLVWRukdFpI5JBWFBerP1nvXPJdpLzNk00kHFVn7SPSVI
Hl/welAUdiDAaGv8/NoJk125+xacgSuOLuQ1WeqmXd3dC/xFX6PDmhVahR2c+Nab
jv0xWKi7IsSoq+ml76JvzLjuAZtjRq2Gaa5re+cUh6BivwM07MjvO2keguJ2Cpry
XLumIVOn2JuBgt7NHge00miYhsMtYkpslddFIgyGLXhZ0LHx3R0S3HDu3IjgSbt7
MHyoITbiGwkDAjZFjUarj6WpWvdnVC6IH/6pHzmdEoQlRPCn48/7yWOmOZmrYAkk
22tWKOX2UhlhQeJshlsvUlN8eKjN+oQ4Ki52lApuFpBwfxWt4B233RP2q4YPoKFq
dzSpa9bkjzSRfP/cvTj1+hO4aheyMps0fKim8e/TZsRHfbuZL5dsM3mHDm4ldbib
sCIqSUyTLFkWrCEfLVvZD61b/H+hCwPGaRAYqA4w+hUy7+tqcjWIYT+SMQoY97TD
LPFrWvNtsUT2zZEkSWcpFuYFNLMZWnrOo7SIo51jpA5dxBZ8jDTnSXZwlJqYcJv+
8sjpEGdOFaarUZ1MqREuTOczqRS5ZR6AU2EkmNQ1MA9ToS/KmxtaVvUhFYjesa/X
YJYQAi5C/9el5owU2cHUZdmsVOwt/hlq1EbOsSZHTNN0vCZraEQZ98DUry5ZyOe/
5PrOlHk5hlJ5AHj1oNYIgx0mNu7SJk1pCFoxvwfpIvG60B6oaDONcldkDUvYhcE/
2S9mFgyV6M7bRq7ksmFA+CLGzsObY95UF+rxjrZB+SReL30MS7X2Kq6MgbrEj6zh
wdVckvzVO6iLiVpuv0EuRAQTYvbaexZZ1G4f5Z6Bkaev79ZbBksaNeBnynJEvhTC
XLrzqIxPenG/lOwFGl8HfJW9ZcfiAyagIHp7UcUJ/k/moraOxq5OhgJe1eWcOHQu
obAQDoTyj9l5xukefs0y491C+Z9DSiXmmCyeYmqtDQkLHzOble4Qq5zNM/+/oApM
B9pVXBUYnDfdNRT5G6DXjEyeDbeOC77n8xqJIEryG0NBZBtK4lFVxy0aBwBOBu5i
xgJ3nH2OwVDsN+9Li++KcUZN4nkdWrmXCRN65csCXZsa4L3L+CbZcBKiJwaSNDkt
KdlsrO5nurtfMWve+mByxbHZGgd3Xr6YME3OqPrm57r9Ln+rzxhpW26Y8hSg1yXW
vGN92EUmbNL6ywTqEihFlD7Wbo1eG9kDESCwg/SB4qhaAADgFsvHK6kdBnuQ9XGR
oJUvuumdbMQVojEnkcSYH7MjjpRh4z8DP81i4fTUq6fnon4b+dhNIK/I09KiGu4T
GkVG4pWRjqvlrKDyqvAy036kU7L45Yij/t4Jt3z6cqQoCYzL6Wws9QFmahn8Kwq+
NoiDFwuHCvBlbs0IMuj23JR70rka8/bGAlTqaOCW0iv4SApS5/R5bQLKzPktY6pX
Qwdx38UnvcueLLI0Ts6nG8MiHq6hZ9b+u3asOhh691pjIUcnDKXc1f4ZIwm9vZI3
bl3E4NLHCFnpexNk5lv2/DpoyFpXoqnkF0zf3vbMWrjCRw7n9A0Hp/AyaStu7M2k
1jkcTzykF2nQ9sU8Ep1SqTBXJrqO7AR0w8q/sgZS6Dfy1CY9oc5uxPPncRrlhclw
XWwSVzTd4niVRzu73AgoK25mYT3rXmduBsnP9ncJaw4qSIcKwxkCpJb73W41CMZa
PzCfdG7bQl7zgDtIw7AVfb5bDhbDTU2+O8pi6lxYQ7dOeUzzzFzAgJyDkSJ+NDNx
ceJGlevzve6UHm8ZjTeSvrZaAhQM1lAbA+DpjFlfeSOhS57Yh+gOSzSWmVQUAy2e
bnUVqtkTu2ZqIRWc9pk/JEP/gudZXdeKoSWrrYxKKBS/fj1ZCz/G+j1T0YSTPj/X
uK3RzBJ8LSH+0C/nDhTEwfJaLx6TXB+XGKm5K2HunIqF2Cm+w8FSchz9fk5KxNMo
19A/dxvwAIoetyU3ok9xrntOWV+wpCGPghIfhZCgWS30lEhKLY4mxSqRzAV+Jjmp
0ZOSZ8gH/sDb4CcGiY5wZLZsFyoNAi2KzZZLMpP1r3XTna8CVVvmbPGBIPcEypHU
j4ccXpPSkJVrb3XLSJbcSn+SbUzN74Qcm0+4fxYxbw/p5FyTDc7SAhSyyWUYQ1Ea
gVBiu2J92CErwWVFjAM8qJGMhTIXS15wqDmtx+mMhDhEStuEqHSQa+FLkz9jIqmI
6hoAbjJ/+j8zWKwr88DiS9kd5uOANaEZBzTBGnI7F/HqBNwkFfntGVY3DeUfx+GK
STiUap85Dbzk8A2rQB8CAa24t6m7BIbCxN6fzWLcbEaCd84/Dz90ECP1CPbXAoMm
jJVIk7AVlMfTKbTF0ys/8vYtGMnaOO/ViZr4stQRpW1c70GFz7AbExKPFB/9fjsK
d6e8uTB3WsbiCM3ERiLiaThbR/KJ/y17iCaFs0boYxkcaSgdZgeOCZaluzYSzy64
9xZsQ2o6l5z74doYynYgOibS3s+m6ngB7KaSN/DRxX1AizUK/QabVob4Sht5WRGR
xn25RDdShH/3ulFWl95KFami51HN1t3NiVj4OQCKbvR7BcyAn1kocQzt6r775YbA
2fmuDmvY/3IAFagoCn3cClzIN1lIigAArMGT0vGlN24q82aKFyq4gxjN7ULOC2pr
H6pLMH7vBgAJ9CkRTbghQbbWOFTdkvccPG2Ng7QpGsUJ+PolqTCHt+AlY1FiKa3L
uizBDEFrXZsqLGx3kVfnAQNl3OmKLBGmA1O5Xz6zpwunVrpskGiWwTZ9MxQs/K4P
uYSEjap7bJb+wzoJ38//iT+jb45cgdRI1yB5A9IQOAXqkxt4fWDDSRJyHfDWunki
UcIN6/3d2SS/EfOE2eVVSgMydGmDuS8zMtqr5Ci46Pr4V7PlBznZGhxc0/ov4l5E
qkke15gQUq+e8h7X3EahZLQCsM/192nlPw6vHYnDv3iOy1rNSZZEYidC/tjAb5yL
GkOOcPe+pyBdnebc09nC5WJ4p3DnlcrNCvCHsxhlufAIjmDXUefbErQhkRBccnJ0
QYNNodoyhrwgcmiw1V9NA/jVSuc3HrMdpi7PsiocW5hOggkMRjkJETyuH2rJXWXU
hMw5NQ1/DSQKkB9z0Iquld1a+dcBCcXxKDj3rSiT8hWn+sxQG7zlJcbJ4xijDLp9
Nww0VTrkF9AAbFts1twKq1u3n4MkpYAjBUgWx8VwUgaIi6u45IO0huCF+KnUgct5
u9gdEycSt2x0N0Z9vLRp9hDmlPqoxS/u6aRNNhedWxDY+Kwzhtmpce0DkR9bNqc4
BDr/Fslj03L2ZoUhphFe8wMYHwZ6vH1qumrHpejH1LKG4AsgEq8E4N3OAv7Y2I61
QOc0RoWcJ9pM/ATph8Xxel5lY7PU+cw2HMREYlqGPXC0Sn3plAvAeMq/CxD1YYPG
ICDcJOyaPzw92R0Yj4m3bKJVRQA+b0UTdOXdolIWkyce4qA8bGt/hmoLeNz/SuRc
S+ihf9ZUAbx8CO3NesRJedkp8r4E7eZrRWcfmDoibH6ne/MEVYUng4/2/ttK8cSS
qWUvUZAjC8pwRbDEQGWnZ5LoAzjf+AIGUxFvuiaK99SltgpZDf3j6smiaYuUZKHk
v8hZx+4f+t2VkxBK2UsYIspgFoMR1NXx9yAGqOQwY4dQGE/t6F8w2OzU693JEKWg
/42cxAWp/GMYVdnLWzcu+TOTePzdzcN96GKLv4BFjEYQeEQ0OsyOjwRBN3nmdRuz
HhNYZ9om7qQbW33MuQNpzyaEkJlLd7Jr8QIpI7bVCCHBKRNO0ito0iqDS3+HFnwe
OQpV2SmSldvOb5YuUcPiyz5NsQdmSNiaVrno92f1navhS38HgdG+++CKpThnaK78
4M5c26CYir/1dItnTP6n+hcFaDI5UXUuMZiD9YlbEyYvLl34PeAQB7BrS2fXqgxD
mEjMPnCbGI4hpmREw7hwjxMqbo1V5X62xhe2czw83dopn9jdx3ENOPKfclhgT35m
EGdmf/TBgPKbzpDF/SYOe8sNPJgPQsNzTnZEmqn+hKbY0IBYMFJDdzN1GqzY2HMH
2ZOOmc34ZqAduOS7tn+Nulj3DeKEy/PKm9rm8oTrz/csDwDUjElw4ZVwxcMNLiKH
xZQItQjmEtSgrr680/A4tWjfYrAm0RKNGn0Wi4uJ8nMzusJNKZILf0UQzjpDpmvA
8Hk0gFdG+/bkltLYCkuPKqfdg6OLKeWa8LaocEBC/6R39MqW/hK1sIGDXRrPLyFF
e3ShoEHHsCjG7r/YhI9POr7axxxp68ooMk+3+wwTyJmOUQ2CszjvDfCgWSfimnq8
lW1bY5lJKTHdIZww4x8PZGQKLFrL8oogbNStxtJFw0U35KXMKZHU81lK37wzDRam
VkY6X15UGafkUso9YH8pNorueXQst2kTRfmj0ezmjwQykNhPSiIT08/Qy8fDnqi1
1w10T7OY2GxtApiUZ1lHEBsE49rQCZxSwIK73SoJWB/JAQ/cbGDJ5UsygIMwi2dM
hF+H4jKele9mM2jKqk+0lGYHKr3LpT84hbh6o2ymsQEbMVrxr2mLMhmnWEQx7cZr
hk+4wL5z5+zo/rVgNjbcaDw5ZCCJ3QrmQlH4iLRrP7GhPpw4GSrywqkGrDMnfyBW
FeJpfYPoCOXsHgNHuh2cy1MjYyUa990tYkoogyq/jq8r1DNiYGj9tLx+m1bibaoz
o7NC3ZpoVzahK3qC1DrVg13nR/ydh343CJ/0OPAPeFlLJoXbrZviyW98m4pzLmzE
aulxZfDqILpI5+ExHYQ7r16EV8YmaD3dSb8niYrN8SrejnZoWYsZTDxF/Ti+syCj
Z0HluFISHXuN+KiSUWFH4A3oxk26rFYD9L2fShcYzTQe5Gk666cGi/mwQEvvUYpy
Sa6RP67ChzTk0ZdmKoghhTPn7lC7mDkVwqSky1Vd2Vsok6aVjTP63NBW7f9f3bAb
bf0CVCyC9VtX4LQ0cJlpgG/PdsUndH8rJbRLXJr8H7/b0Clg53ZxzjqfS5X0d12B
bg0yeZRseJCz6Y7gDaXFUMO7D/JxOGOx+Xu7UQq84gw=
`pragma protect end_protected
