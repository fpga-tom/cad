// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:45 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GE9Rx8JDZpXHUOXfZmimUPAl7RsEfKbHj8ESfNgnGabaygcAr/RtsvwT7g32F7RF
xZ1SqLn3HUs4MAQEg/NchvnH2CgFqlv8HHizlaMd0gK8ndjI/pUgizp7uRIK54DF
H/idP8rqxOIUOnfcNlm0O86TT/K2FyQLs/mblDw4Jew=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15616)
ACxxFhnmiX0B+tbnWvso0jQ+uKzqu5OJSH5eUqD1eJqoWd57ayNiPuTYwVWdMuLV
4qQLAqOonRD2IvNwxEbA2RZZdCJAchF1Dr+Vc5s/bWVOu/l0P2ABrmVAaRklunmL
7kzEddSEBajrFX9WmBkR/fu1GCLwMxzWll/b0YbADI8VEOLleh+GKmw6Hb0HS8Mk
CBYi/oj3NcHzeTxBP2/WZDAutfi/38cQ0I899SR8mxG6eL37iDinYagJOpqMnkwZ
nZupbAVsjXh6RisWzvcm1ex+OpDGBtRPT/fxSEVOqZkM0h2cDcpO6bufjM/1Uv91
EsvLB/GTbxEyIhUUis+pvF4cSEpmQF+Gt4Y6CwuKuRDzCtf7gKZViSw1ci0CMM/c
yye7CmWWDPRfxdTfEdv8LawbAe44EOzbHToG5vUXljGhYCqYr7C5BvDcpxISLFIC
buw7qHXTpgoluby2NgJKFKQHjldGe1OSPmrvearJV/DlIGxnL/EnVeLOaiu98Mr1
RCuUi8df4Wp0PKlB+Se584VkV7XvaCx4TS/8s43qlM5vWxQaVlfui4DV58s6vfI+
Ql/Dg20/CaxDaS9bLmJcY5mURRtV9MHkCRHSF07CnvBcxkCTGq2e0IM24MBoJiH3
m60MfjyO+ZPF9Qh2UlNw+S+OVeVxkrvqPeVSDdquH4Tf1jxm3x1hmbdt13l9vwZ4
SIOHgmT1tIT20I1gZQtO8iDHBXDmvRhPirLDtqzOU9sG0itqrmFjAb8PVZgdJSDz
DTFM5mVg4GVPmibO1QQ3YeZSz1uLTfVpHAuOTgW8t17+N3MbuO9OK8gs9XeY1gsx
HqMI2LNAE72HIvYKiTX1U8v3FcBpbCJozBFkq4R0S/0CJgh1p+YLumiQ574+QPn1
3qwgPEq7FGH/PlwegCFX7uQCs/gl6Nc1Sx8ZqvfiU+nksZmvH213BNsNbe5NEzBR
jxtvU/KVixo1Utqk3819nfeClw6xUrVf1gMmO1HN80vSYu2kCpawiYq1E/twPMIk
dq1fXVgrTb9Sj4gLSkawjq7vExnBICFheQxWkjOeRDe4v8mVshaDThhmAazDq3Rb
38gxMiG7DyRoBkKhRfF2ERAJ+AJoILiH10vjSnmB6CDBRlGkmPLHVOCuUcEkPxQr
VhjmGLvTiSLFbHDQ7h6ewCIVR/z1HxP/xRRCkPgn8VIFz78TDXgiGvcFTqK4NorE
rMhKBubJoSfn0tBJiSNiBgG6efdfQJk/hWOGk/4YTgN8baX3pIKq3xLdn2tsxddi
0k87x5ygr4ND673G/pKjUFMsZA3f+wClAOgwhyRhNxkv9OCXU0H5jZJG9MoaeHQX
koUp3pXuheTRnrQgNa/bSfZkzT4KW2d9zAL+yjyLhYc2TwjdpGNVbFmPxE4/08Uo
G0h6zWys1McVVhB4IbL4QH4DtC59XsMV+DhKOWc8qzEDgPQiBddBmDhz5lW7bbvs
g2iegEWFS3+AVnRHtK692/A3hwAhhtfhjIhOUxnSXQ9JOjXGI/zR7k1lBQsaDENx
ouKTyP60Nc7zD/XR8Y9DC9Ph2eOoxs8VbyNtyQkHhuqb8jGmnJv6WF/+bYyEKefW
gCsnTnJZHAKeci04RKJVzCx96tPW3wn5YG7JdIRtYRJbPZG+LzmRIuD3CGPuIRvi
u72RhrjATbxI3Do0QZaaZqFVbmJpGzX7gOEOVfhjsDij9MPH1j/p4YqdWNUXnZoi
VUbv1bcvVhPPJ2t3LJ5dNB7uMxfLa9qT3Wv9P14RF+WS3MEPFPYTGGRiNEas+vAB
LdHzblabK8Xptd0LrcVSiN4hgi1n0e1K4bAFjqArhqRuBFiNKpwq35eCxLXN0YHG
GBvM775NdYTKDPkpSPSMsxHAD617qq2Qq5eaBXzuLneUHMeaRh+Pe7G2TSwfZlNk
sWv15RSf4QzOUZvDIi/3F1HXoPWkC3kB+bMePtCpJ1o5aLXDSC6hv5YggeRI4/oe
6abxTOuP2px3SZbnjsCV3CM2MrXEEWgPxwkPeW28UgwzH0LzHRXd+hopoiQ1y8VX
u+JjSa+xnKSll6LYQ4yxX0Hegxtrqm7z/UZ0nBpPFPFwa09KwF3gRB3xlvL2KiNW
1xtpW3boHyyaGjkUqMdcxK/D1PA749SLNZgRhyqreQC0Q+cn1a2LU/o+oMp2L4PV
L3TuaouzaKvFpWXL5bLRjiNqPEvxfT1JbNvHmWCvaV6gui4SWcw2IxtCcFCcr4q/
Pis2dFVfdjOqxcoMiKLvWaIwYUyyEPDREQDdy7SVOjUPSDkPJ7Q2LjDtMEPgfyeN
QSgmyuUmjFyDEm4CZT7KR2o36uNL7tIsNPPjlgJznE2L02v94CQhejmsoJPP5Www
q6XA0HaBE1SPUpiDXuUEOuBMMqmUEwiLdxIeGDbltFhWvcGELBr0CJ/Y5IfbPNVu
+EH0x7/RhHOvSX7EUKy4wJVWl21d83Dtg+Pz4Pz6JBb/nQiW5Es4AsyaQZ+fGtSs
Dp9WCmabFaA0mNsTiQMF91jd2YzHTVQnSk89yBUwGz/5XPiKo2LPlY1bOva2axX5
dz3NAT2OsHmGmTqgz0cKGkaoDfOh94jkp81OIevWv6reabdnNrdP5e86n/XvtCrk
lfOEsBTIUo1Y6E81xyq2FaAEzlv1jcIyXmOZdyvwKrYftSFRALwX6DZidDc7VEDX
syadfahXBlsxCjx7carGHntpvRgKN0DG7+qiHlF75go+bkHhNtdnvH0gcJzjlNvn
ekLU5DyQeg5z24lPZqFQnZusOSoexjuhsJhBW9CTCjCpyK1AWFMkcKuYTLp0t7Lp
JPMNz6+lwM3KtleYk1PC49lE8Ifdv6w90rOe9VUrkPOoehLBnZOjSHRfFbCGsdlp
Y7KCM3Qf8gQcgQ9dWrR/0TpXb75b1DdB66wm+cwNwUDbUb9dAgjHFBfuGQA6Or96
YOhQajGjLCHUUKcRDLJ0YSwNUpufHOjDgGUO47Fh9f2BzAA6U/5xcrgDNS2mGAdZ
wb+g86BOeMEQiHIA9gPwZ7IFMI9bFV+/56P8srijvmFJvAcuvlF6vaVQ9Z4Xxn4S
d6aFjLvsGhz2NW8wn6ZMw5ftW9pctKnBWaU8IBETkp0acT/H0+3N2bqw+YR04jZl
h5lqlzQTxCWSBvl+ajHJd2KLONmNYIZjif29K/ExQPIt7mCZKWIrEZhN3fQsrkWe
q03SxPDk8qhospdvUArRhGB0ke8awvGsfyJVq/RVtw225PYVdlNkKRiHIi19Bck8
wNuV+aZ481iZ55mxGy+FGOiIwvYX7V3oEfzzeTvbhpgjXZFJKzlEAslHCX1OngOl
GDLzpCcakZoVA+H7LsD7Z8Ge74jtK+gJfFPbIL2it0GFbBUWbLm4gJkmHOi6jc2R
0KClMz0xmHOhdM7bPUBUfqA1+3q7B+Dv6gSCY9k/an69VuQpO1N7VR5UijkjzSXU
pOcDEN626bHYO2mL8NurNFCI0Spq+aZ6Or9qf+fh4AzdnPNQdju5VqYGnpjGVNlC
c7QlxeHVzw40zykj7hgIKYmgYBOouKAUGaiedjdXDJgbz1I1sV8F2B0HN6V+Njp9
tQxpwXOBHqLol4eL4QOU3LRVg8NNeSQcOgqw4GAT1WLbJOIqwKSyPy7RDuhjEV5I
P7ZSEKCraZfSUv+7pGhuEYRO7CqWnI3Dt9/XdchgWYdFnx6KyzREn32ZPZHgF3Mz
M4KeG0rRtSsH+bHvqRG1TmxbcI8mwtuf6wqeW0qyMF2RVVySneP9S8+LczzIxlxU
6SeI6MWK77ybHJnD83SKtmJ0I8dIVhFgGIPP5FPQKzmzIs0c2A9KzufvR72CVYPV
ji0CQQ0YWPykw9K6RTeUXkH8hkT6bav1JPbm65ICGhe9wsbUykzZgBUaSKVox/hZ
QiFkul194wR19F5flgrZP6u9mIy82rdO96ijqaB86kXVkS94vwusXndf00vLVRy7
GGaDDBohDZyJ7txhbOkfOXuDW7nM8BBn6UOLFjwzyXNbLmF6c3EELwozz44b7qVy
Ui/fe+18XnSgc+/3x8L2ceXrANUdGhZhdylLrhsvYhGE9QFhuozGFUyDzmZeEc0A
II8LH6x14HlpHo3QvLBM7AJJYmZ03aj91HKceGc1Pe4YT/sBxVfytO+nN7ErNC4y
XXz2iSifiyA2lg4+vrTaM37Qfl2Shyk6HUtskto1WEG9yhrek3JWRwoFXBwTlMfb
VnEjXUyQER4iGuzIgJulQGBOVruTWIQBF/0UZCTEbZNTuSeMF8r+uzvCAS1oVpN/
spI5PS8Dko1KH3uetQVl0y2uw7EaTsttPwtwyvWiEtGzoFC4h882VbKCcEqaFwt1
vS3VPbhMFfWTlFnBW922N0r3T99S4owTY1VtxlcQ+H2NokovpKxdDa71qSKA8G3C
DMffV46jjstoTCyqCDrttVtaaRR6ZGOGFDzUKNKV96E8M9dRLgjmMfrvblFTyc6S
NKkLMkALR9CVg4VdH4XP50OKCtAaLt1NIX3khv5Sb6tuZyZVCUWGS1ndgO1mE58H
kiSKXjNstnLl61EdPO5JUHPHTnVoHnP6AIW1iOpL7N6Uaq+YzzU4kDOUTIb3idkq
bM19aD4B44dx25a4eYpupY3WbzZb8V/r6if4OULInXZEltyLFRfEfnikQLvX96VT
fFxZHNqs7d+J7SeN1xkEHTlkZnOsrv6tnHCc0gcAw79+9h6YTPkFq3ZHTnEkehon
iqMlTEdtzK2T9eminCCJpKD9sN2xLwuEPP1fy9Hqj4cgainh5DwixddgGedHXYC1
TknZXv4ndLmkIk90rVwKSfqvonhu1vigl/eQ0Dzctq9PpPGWwJqynieKLVCx4feD
0qKb6S6igX4ci0mQsw2EV5GFI/lxNrUjGjdhb70lG9MYKVsnmilcFv3lCq2K3Bet
m14YpaotY1Bz3zT6Te1TL26q7kBFnhSg0UlzFShjoILLjYcAQ+YAyabFz6iMQgmZ
kDzSiiGKZQ934almqka+H00Uk49H6ph23TJtAOtDrjAOiFt/Oeiquv/0YpbLK+AS
AMKGHP7QRdcyfDYswRv2Kmo8OsVdB1+PHYOaAtzy93A6ullLVPKdE3+bx3pOzk/D
+Ep4GydpwyMYlDgiPbjDUpk5D6CgwQQwCuDDerdu2XwIIC5jP0P6v03X4fVHFR6Q
oLc/XegBCFhTb2ntVC39Sgc5pjQlJx4pZLiwEFmZPGrOvBh019JVr+CSNhsjUgXe
QeHYSVMMxl2sGrz5XoOx9j8WLK94C6Rw+J9Y6gyq8Oe5ZoxP0AkW8V0ToIWG/qlr
WPsku5DapTOHNpR10g0YA+il/82eMGJHA4V+Id0ANrQ520EAUrKPXnWsTexeX+zg
Zd0zhkGff8KBCsT/ZdnIHkRY0hJcXis1szEc3iSDxG+Gw4u9ircKRE/qBI9NyO4q
rWH/3td2+h/t2NH7jjs5tiNSn/6uWOY6vmKQV5Lnxld04YbEivqt7/qfHGeHJ96K
9pcNnHtFBljZN36jj9h8AW7h9H7dekkZqHiw86o2QNcnL5Kr1ZS9Pvh7y+HLoBZo
/I4rz26sIO+b4A2u8xBxo10szHeUXIuomyfjSNVgTV9MNBPG/jTOOyKIp+yY9xGZ
jLhAI+gaOmvitR1dJjf9RmjMgsMhycnrOI49SqcrbKsDeICXEtvEUnBozcxhCwMT
Nc0eJe/4MBGH5eDTGVZDHa/8Kn0fjH0Oy9W2xCOrFCcr+IsQiUsSKhRkT4jTC411
djEGszxju7bDTNdDS5XQ/53KXD6qCrYHtIcTqej2vBlw7VvsiEy9FHlzSdRove/T
gsctr2Y9L8o+ryJTv5LS0R41Q+Jo2dcm3RTXmmidtBH1TquNGqwvtQ9gafGohToj
zQJ4YG158/shi4yHAzQ2fdZCO6WJGoVasp6ODMezBg2SToEbzyaYJos6SkUVFueC
asODvMqHnrAAzXKH0RmRl1kK3NCiXKtb+nDA1cRMGucwUWCUnOphQXtVG9bbymeg
89Ay8WiQeRmGdl/yMOeUbUzvTSLiD6UjiocwPSUDKUe9j/F1LmTN/37eQnkuU8vk
Huv6MnqR91UKLPLSbwB6VhPMdid0UUaYa6/rPZ+YNxZbmwIlE1JPzEk1KSzxZ8wS
jrK54jmV/r1a0/P1zOqkcCjf3EjgV180Yv0jrpNqDoqrzWfB+xVa8DH/GXJcYzv/
9223GDNfBeU4iH/VACmUkfOUhiFVLJrzgqCS+hKKJMuDzFpHsuXcDcySka3sKrNQ
QBI9gcZ16coKvOxb50ST8VEAHYX3u/6yt7xTJxqyZCWFif0Y6qQjVCwp0xfzjCYL
GzVUwwBLQEi4RtNIm1KBFZnlFgr3gg/wXYnThUXb8Ugmi+NiZwOAJJ4oh8BnxoaA
9wJdnRSi3ppZ3VZNHvI1SjAxvkch0lWt4ZvrC0UvT52xTKcBv16xeFNB+vxIVW5f
RBJnRBNFeP/jIujG/wE6Khe2+AawWVIwPb/UUppKZG2uA4hKX+V3aAqr1mhd6CEZ
mmFE/FoIMhgDwIABhKtpmZ5jtKbtE8ty0Zsz7/B5pTiMIfW5YCagm8Bj5mT7ijhE
teURyirt/29w9RcWUhxt45gImFYD5ih+p1bUVGSyC0Es14Ivw3IpFNTBThl4T01Q
GivSo0ClrA5bCTPGQKzqVXes/fHh3WlMWpZpMxp+E+q/fv9cveqQU/Zvg/l4sUTd
IUudxKTweLGDoL+zZBbtDJdqi5nUAbzSSzRDIojwX21y2fA0+ElhG79EAVpWQA1f
IhaMFO8lHxtGWCQbRWtj+mEFJX9RtF0YPUBLqstBKMVooMpaQxQLvw7Be7t05HKy
ry2Xom1rSwTwM4uqxrRsixdP75fw4Du+L66S/X8s5BjJPexlook+7x+eKy7aMEvQ
ZUXi/g8Q0jOtgSenSLJxSypK502lBOwn7jge/lkyO0poD6Dg4o6Sj7lSGIP5R71I
nXMbEANVl1/AnTz01epbj6pm2SbDdGDgnAD3abveX1NGqWtRQ8ndmrm68Lt02+AX
XrOFSM/kaar4cdC1tDnADkUIaKdlzS5aWHrb7Z9cUB421B8yu9ulgCrlK8/Ury+A
kwM0BYCmbDtEQpt6fr7EroqvscQ3pplPol2/60vS+jViL8FVc/vT/bdLUv2VVDTa
RLEnYQS/3bAHbYY9I7FCFu7IEC6UgSRljKrTe+nWcsGe0EGETKuFbrHuvbjazyYz
xVIUTidirsEhcR50bdJ20ebxxog8k7Lk2oUf98jAtz8YDMK1JnxcGx0ET3SULWTl
owjX93Vy2Chlzq4BoSwbzSzHLJNxI1csTS97sVSQ5w69q4s5K9yz6mCXpAdyX6X9
AET9D6/htj1quiqxOqdp92xpp0T73IW7crIYotS7HkgIr/tfsjhYNzw24vO8NErr
+JR5NC1Wk/GL8HwdbgA/M1mUn4+/c6tOu45YAxfrFLeKenIqK6QLIk2coV3ROPwZ
waEjlukbh83uymr6w8WHowIESJlCOUI1xu/p8davFt0G0ip5Zc6D4ThnbEHZT1JQ
cx6KKeOBj5Jkt5JoRBHn6YtkjIRkP1yD4G/jVtIHbz1ojD+0eqIGlIJ1HSfREx+w
tegMW1ARpgurkPApP3ksnq5dXGJZFbugFpEsg/Hc1w9AE6Y2KYD+zUKpgQVN7SC1
3cZxgjjYYlxMcZlCGj5atVhXysTPs3dsbLhYLwxcQi5wvkrZN0BEiqf+tkpdEyz0
Jy9qbMyvJ5zeMWjMipDizk3h05wGK8io7SWPQ4i1jpe3lYybVt2w23QKOs1Ow0TG
5FkUUqKn8lhXiJ9008v0dHNxgn4opEpOMMeh4kYkCKTlWUKdrtCnVmFuShPjdAC1
hW1HJGNibFkwpEUzj+L7A6jqkHn1z3z05+CElBYvzfxFbHNPcXubxX301iSJJrmR
iHwgq7XUN77Jp1r5UFpddkLFduVO1t3fIekVkgAsy10n7hBEPj7bU95+nywjSymZ
6HjZjyRB2xLRQeOyd/YV/7W8mb233O7qhXTYd3ptMVo0ENSzprM5OL3mYEvICHn2
oP7ty6ihTKUdGiZ2tjUwqYtmw5fk6yQDPq7Cc77162L910hDOmXOJT0ncTx5ZtTd
+omwT4U6om1cx3KmGruBZZrECSQt7um/njEEKs+jaSz8J24A1uWdn7T3uLx4s5y2
cJ3gpvFwYUUFFOwek3jtdichWmi0QiqcMUdSHFjGqNVPmqUEB+dI+lXIkskL56rm
koFI6llERdbp/bWcVLLFB3Iv1Snu8A4hJs2ekpe0bC52sdesp2eCKsOqtKA7t+yb
dvHv/PYk20ciXuQPEMjiif86ysVGT9fRRtExVKmnLYLs3GFz9oqKvcmfBy7gRh89
pYG0dVNtrCGY0DexyUt0YOCukyn90HY1/kAtCHVeXPtikrJotsuVQtvdM1dfjF7n
mZR9TdIa2DrCaMjKjC1HWtOKTcn9Ujbmc+JCqZpvf7VlB/N6wRbezRyYgsV7WnsV
FDjGBbBJaSLA7UUvWpDB0ANhICcWn8vmNp+Tos+jA6ls0v3F8Nmx7Atbw9Tt1MfC
MBg+C7iUakVnRTw2qsemMCS+bxc01FMm6ScYOXv8oH8HB7tHNcuE0Azq4bL2kH3t
GXKuYdbBhBp/SU709aEkQa92dgvQC/4Sx/lHhepI++vv5UyTHcuqdvWkEUvIMKes
KdH5Bivvgi9dCr7+ddQeXQFJAohZoVxPt8dylOiVwpVmPYGtrG9fiU9CUeB9sScU
Lv29PQtd5zAWQJFmX8Aei+UcgjzT+sJ2JsnajQUrLdd2jshPeqW7gwiPzmoqExjv
T5I5PnNb+Rf71z7cnsodTNd3wBrA7CKT1vqAUxhGFjWi4QD0nWN7AbZPa6vdmRQq
+GE7iJXwEXAj8tMGSm+/Uj2z3rqpxB9Mei8buWCJZNO7J6aRpCyxZLAN8YGTX2/S
U787hGk2Le2JXI02gZxRwLmtg6igMs3cgNqO18yfTKPEXHn2362Bo7UdGnZ7oWll
t5z0T9ymnFrpo6IARd6ct66I/WAIy/CWtkLMRy9RDXNg6uYGNRFBOXYzE2mXyd6W
GUV3p1Uu8TDj9J16LvarpDso7ikTb/M0V1GeW+pnbNX2TogxyoP9B8OlpYWyp9bC
4KeqGCj3IkyJ9sX9VeNhDrVetnypYg1vj+h2O+b0Mudlzugl6UsSEr6g68VsGtRy
C9DhQiHp0J6pfOXXJDWoHZznHYnl8kniw0rkm2PhWcbdjET62pLvjN7UCB6KZHiq
gej9FSGi6yiJWlieF7SVoIMq7SyyQmIs4Xjwa5FaYfwoIo6VwgawRlkq2Mm1zU+L
74+c85SE5bkRQ+5f/1dT/vrysAP3ggPxIIOgPfn2vrpL28YzHoEBETuF161u9/pn
odOgPUXFoxSN/Nc6fOifCiE9782g8pfJcuso28EwO0/7muFx3G/j3nZ2kVH5sgNk
A8qBz9iTSJHJx7nu21+gLNq/7k8xQcfHBvBYFu+OAzLaDJxQvNBQjHrHCtXdOr2+
Y3/nwDodVDnQLOVwi4mj5PTUsYIdIIW9gTi0U80KET7SgzkZdupjXrOHPNjz0uJD
AgHkkxLN9ElqQE0RaTsjWmPe78nKNBw5BHJSVECEul01zzVuReF/2HgejXw8OvSm
iKuuOtHTLhXUaNJkqOPOBjeVJ33S16q3Lh0FWHpL6Afyi0xiBPZWE8gn3/5BmP3f
/RPHnkKf77Ve5V+seWNEDhE5ZJY1YmrlY0YduTp8QR4A8AYj4IzytKvWqH8+Dqhu
hSIut3gQrIsArutVHZfqHUwOoTkL4adLsU0QZZ/gEXUlvh4hcSQHgC20PSc4HvAO
m1nx0F3Kyt4vvZu57EsS0O5wKAEJR+o6c71oDPr4SWYjiZVlQl2rG28GX2kiS6ST
9dqRlpplb5fZNDLiOoJuqtpUYdxYkGWxsajhgjOel3oala/pu0Ubnchne4hGUrM4
XRLZ5W7wfaO0g02/zN6flX1S1fucwGcSbLGKoePnBSoY7Z9ud3W03T1BcGbDmwBt
5Aw70DThWfLLO0RXJmrV5v5vhva8w9s0cOsHZH85nEgtF5WjT//ySJqsD4+YvpqV
TroyrbyXZiyMArTR5nyuA82qM2hqGxnmes2Q8ztl+khTd06eBT1NXH1D1s9w/KA1
U2+aU3T6z/ijkZGZ/NmG6xdKKICaDKOeWWD2ecGI1WctAO0DpH3Cu8gBUzISunO3
Gm3PqS+JGwRIHHVfWtTZQGQ9R0e4KuEybk5w/XbiRJmEsz3C6C7C51AEPXwKoYsN
U6yfpPtkyqmjI1de+ZOWfudIdlFmP5Wj5sZLDoK2OOzs3vnbfSlzTAmLm4zbW0qT
PkLQklYflinusOq3EM5TsK7O4PlycDNVOmxXeSTODhFV5iithIjlRGd0mOcssqV0
LAPynwJIzuHqbwUxQvuImAcbjch3w+zAR64ZVpnReqU9OPiYLNuQvMAoMULFYVcr
/9WfkKyE9axgWiIotrCjAPae46QtqIWC3//7YA07vHhF0tb3Y4eQoWMMyiCgUJcd
SJMtXrxMWqJnuwvzLl5KeW01JxqCpIwVupBnmNVNW8+DEcrjbSsZVyBr2uE4iV2m
bn0goFdL9ha71QP++ksiYcU8+PaRnep3gcg1YHUO1Sujma3A4ErxLaeAkr5ZJsGj
QbTT/1VfWp8561OfY3/+5aa2Sjwh7Cz063C/QpBMEJjglqNannpcDH9OmQm1qY11
T1rx8wwwhE7TOw2SJTWpNHZ97nAPDZffU1sDRU9MT1j4R5mYEHZ64rI8ZLodkfHC
tqFVb1k7HBMLM5W3avY57hqScBl+SpHtLGSI/uo6VW5jjE+g2/TIyCleuEX4kQCP
UtDT8aOc/7eNeIlz43YyEF7N/oReNp8w5NwPcW9PXQwSLA9ArMEDnG7eakLtBroo
GxhXcJw5iGmj25pJYoBmbDLQty1ZpCQaeBXVuwWQN5dweNbPWULBF/rxIfo+AaMe
VFa1A0IrbIefS2kUw2qyYg83rppFo6SXgFMagTzdLWcrkF+6nw05/SSvik+plvfe
fk2rFqZ6AvXT+P5IWTbMkSHM3f6wOYerUL/e2855D0i4T0O7OW0FfX4moHHEzUzW
s8Iftpo4lzZoj2XDgpv+2NOA8GGGKUaay4X+qcYDU5ZgOqRd8j9Z+CsFSvRPu1LU
YvY8s0IZIj0aWHtMzZ9a/bmCm/83GZoO/TlMkbMZSCOPe1MJV2mFaEcNeABdl9JH
Fo1KkuBU0uDK8x2rZGFgwn3C6w7rpHSaZDYbxcdxSgM3btoDNMEVvCfKBiOaE5vT
ri1Cc5WdzTdozdxiFgx+7Klr1uLJWGQIIH9bc+UXbI8SeHmjbmwq5H17fyXq4y93
Z3lTQpubfyXw7AWEfBKPhYzt2SWvSiRER9twXbHzJf3DCFvBKYcFCdN4/Bwb7aNl
fY0DDojKSC6X4VRitTQIbRjX7Z0kmGoaPdeNvs91n5EE55sZDSDbFbi1IXEKsy8B
KrXvJCgw7zXaVHL1czDc59I4IlI3Izu/LmZXbZS7B/ipVxkaUWhL8Z6twRDiS0zt
kOQvWhAOxcsjuxBXBJNK7ALEockPvWvvyecjKzIHgu6IYjYGCdM5O31hU1l6o5bL
3iKRRwRW86xlFo6Z4V4Ey7t5koM3EZZQUXpBTx0FBbmTHUDuJhKpnwI8qEMoi7I9
AUfZARnGrtu8q3FJ/cdncbPQ80kqYMlWcJTnlp1n+38ewMWspEn68wq1KtAqybtP
cLa/bc3yGHiLp/xSntVBPL32fomuAzANOOtN/J4XL7BF+1h6eQZS8riB7wS4PMln
6ZQslfXU6Fd6RYgLMO9BHwXFI4e3HsW5dtOumHkF4fJC+qlrNRqW4e+7C5n+d9YH
ReK3YGkO7IsCy5lqbj9YSsraIR/4mMkAjQ3dKYfpe8G2tHV8YxBmTuXUGZQxG4ay
1YFPRlAb6GDl7VAaZasOB3/E+iiJ0vodlv6TIH0SSHxhKe3EHOj1pGtvGkqpoIU7
k699r+dBZVcbp1leUl6VVSLYpJjTUqsG8talDQ5X7ZOcv7XGb/kwNeJSFGcEiUKV
fOgiOHl5Pn2H50vqCMUBy58bUJEje6qpDK9EfHPDlmt82kfzafuhDPNTmcJGdeXI
ppnMHmPxGhr0GiiN6jpHPPL+kL0/EO0ppIdtCTnN7SH78wfEYe4xa8o0/CUYv2d3
RtHzn8rKCd2UFBA92aVMcbeq+P0yYApFKd1789l4SQeGypsM3HzPEGkwea3jy9ql
F0bcDD1ZsezFjbvCqLj3oyy52tnj6ykE3r5vNNJqUaNuxPoo/Eke/Y8aFDuPngnR
cWAUqWikJXnXuTOqu41nGCBz283b4Tpjicjcromxb9aLaQpCVZjRaOcu/ubOhTvq
ls/MWupFJAQ9GvbCPu4bnxqFl5LPL9qzMzU/HtSaZHsr8R2I7ZNS7cBFyI4hZcrV
XddGDncJ+4Uya4ernTwH8b4SjGTifr0BEHjq0uUyouIeaLWmYYf0oZB4Pu6q0xXI
IzCitUGYuUg9VbF0eGDVXnXFN/1GGOpHw6Zg/aIV0P3Ps1f3Uf97lHpKf3VRrfkw
6TTsPl1GgvFIqXC8t+mOzGXu+Ir83fxH1j9HuytvaSZ01+752ajJkptrMWUtGQMj
/BIJjaY6bVKpHB0LMv6G1Vg7qkFRkbstrWR4oanEeB6oW6soy86ur9DofDAGx2F2
7BuoqG8C8GpcLLV0WeoBSfOI5xWXE+8qjvI+gzNctF154AZRHxqHVx1pi0WoRq5N
2BajK549fM4ErffHZ0hqQn7z8tF2ml6QFiIKO9y8Q5YpAPTxXrKxzHit1jUQ7MQI
RQZaYXnXPhX7FcInm80AM7qznhR9m98vXtGSBmgcu3lkzZu4R00n+igewUGFFyCN
SexnOcVhKfBZMas9YRXmg/cPxL2U5iYJBXKl44uLkVGLnZVMlosKLd8rdZ5fb4Vg
mRGd5Bxy78pnRRcExp8bl2T6IasdRl5Hzbl1oQNsZkWkXajS+AAz7HUL1OODg1l9
oQjHtax4Go7d0fNkAyl49kfE/oL3X9+t9gFLZoItJQr0izItpF0/iKHFGzZuvZ5M
pHULKZMEgpieefhEeOzD2kGvJtAaITw+YyiyQDV3YOOHhmu7VEbCuuHUWviYde13
Nqf2yd7yNHg7CFMcXi6dzK9uwNTX0L6ddcM/739wPmifTTmF+4SCZvvnWTXr4la7
CMeITlAavsXD2w/OD/Bc61xKTJ4EGVmV/QmBJIsV/JjB+FApMfIgQA+c6GuRR7hy
MQRC9ctPj7AJt1MF/zx0biTGbwUGdla7K43Gxdol0oJsGKs02wfzdhLuKXmOKQxH
S0SBmgbRwFPxS0e6MucgH5l9JVciXgFFs3pdj5rmx65H91bhEEQHOC/4BgA9Rvzk
c0f4M8HezQ8SdsdkLXnfGGLeyQZcyv/Ivvw7zoK/zOly7zJT8t9F/kO4LY4sdbIz
YAibrmVKMhiP2pQwB7YzAK9HJQF5S0xfnsAOa3ky7flzgRicetezksy66RF2RUE6
oMiR2+j3hQpvEqLOQ6FD3l2AmjzkxJSJA9iDBuKkfnrcKSRqCn16eznAAzaW/rdD
8uRgoC5/ZcPkCERwKUvaEpDw0Uvzaf1Ty7Nzi7cenTzjHnc7Ss9DDRljwDqiPTr+
jCdC0/BgCJJTyXzOLF+g4zRbNnRQmQ/nkYctZAzbQHApz8a987IKGvzPOMbQwT1x
vTlB3hvo2r082IXLGMS3TImISulPuD/ARM+sIU+Ogn7xkw/zQNcYPPP4gll285sp
kIN94dvdYOUi8G7nDZAEysXF8ei1fm1H3uEaPhE6n3Waibjpdbh4EJ92YRZh3OSe
naJteNChV9aJZsPSxTc2V4iQxLagqAr4NgxdaY2UQlxiRRnLtu3wAx93x7WciP1T
rh/PEWDE7UDN/41V76gidreixAnOKMZIcWNZ+JTE9bQcEMfcZK3MXFge1asEocL1
1SiH7Pc7382wEoIsAINmKs/iLoXYB6A2wifiVyr12H34PKcEAEktZWpJsrPZiT11
CaXnAh+2KPCCB7Yz1JV2HRu4UnnNdU0zqc/zi601e9CBjH5aqdx7eSCa+kEKI41k
2iRdo75NYNGtyhEG7api6L6iu21vDwbGRPlfXra2Pgp16pPV5ZPV/UcuaYnFdZvP
3Waulu2E3IWFlAtTqUcW38NaACED1JU/idkyZIAsIHr3PtPZzTyC3xlqyisqJGEK
c1RIG3JAJZOo6aHTkYRUNNTHR2qd+tYm/5daVxFub3vvfR5XUhn8DIIgX72SsUiR
GUtMfjGfadQUuiu2bYN3FscyoYefJ0fQp+LebG/Ui0HzlUf1n8MoiR7iaXzGgOpn
lwAi0VuJJCFXCK7zJfP72aJ3Q8lj7EGQIdRNDobjPAFgC22tosQrZYrWWtJjmqIL
7axUmvJBY4/KiA8eoWGd7eNp05tr9zgcHwWObv3iExqLkqEULasR2QPM5Hdkyjgo
y7a1SDQmiatkcoC6DgIe8IUdKZS5PwoGrqGWpn4bxXc5NlXl9SiQMG2Cixp51s7c
5MG+EphAjpyNIUaE7VR38WPimKjRZI5yrZB8umCLWx9JT7Dc2912jEZnC44ajzQ1
ESRDY/j9wT4OReMuMnvxPTweUyxhGn86uRlpYudhRmdSydlVtnilQVxBlqud1Dm0
9qd8BSxITbb+ZtmxK/XwXsBW/K1j25+50GHIn/uNxHLF503uHs8sJTnKWUyL/Bf4
JBDm9M/dNAIj3H/ABvpJDCzn8MYq7SVpe01DiH2mos0OmNW98KKZxfduJ9j4+P+r
nYfNU3Qp5VpMWi6KvsXetMmDxdSr1cf9vbeK+MIdf/TVnrMUGizPED0iTdfJJrw1
N6C5QAbje3aTcG9HFuSo55v/t4h8zqxaQA/03CDXxQ4LDx/WxnUn1mLJ00q21lRe
f6cIPHqAIWRnhrrM7aZBJbvvMx51DkXXOBH1FvsM3KR9tGcbogu0162afgMfZlbY
8hn4Hcp2BFgB2skPgiJYyljgqXH6vFiYDg8iD/ATFVmWSGt3QJ3CljWvcgvIxe09
v062OdYT/MjXoNUG4zmaY31PoonA7xXn8FLA2Y7KI+yLcC0vizJufVH/iP5Get4B
reA5X0IAXG6hJ753BiBmZ+hmjXZyx6sHXReFiXIBeNfJ5ewnTjuPqZXhl9VkwomF
nE2MkVK4VEw0KeTVNaQ5Zbys32F1Ns8jrFkKGUT2g4+wOQOztPUEFSR1h+BKwdPU
Fh9kqLD7vLUPNr/tShPh/4DnU4JBVUcnN1f06J1Zmjm1tOAcc8ZekIE/GHUFLDc6
ZCSgE9fEPMRoE4wrIvjj21v16YArkp2WrDLoX2o4K+pLL7OTU6mf/4A0cclZ1Dal
To/BhLmZor+TsDulAHfCsyI1XDgZdAJQDm+njMMAW9tigzzpNbyIJpbzbv1DUjm3
tfUo5iVqAAp3F54M3XKFCRF8E2izILnTid+/eHwSnOryBxB/Ykyp0Y8jVFz2Ag6N
gADzgG5kjrM/58yjCAhVZMHMcly8Cw8/6ysef0dAZ3NgRjKpDy9tTtAcgyVGS9JQ
tdFK9HrKsU0OWeS0Ta+8Bf4Z3Bf9NqzYcA5Mj8w0vnaWvU5g7c0hMgGxZ9i5IIFp
0cTxnqLTvq1JwM+pcpIUlfjMB1nlU7coiZK2S+XdYZWEI9Ukd0x8odJUfUyeD44P
QUL+O08pfjvPTVJkD+0HjZ7NEMb/Aa3k4srIatZ6jFOYvkj771KYg/gzSJVrXbtW
YNRqLL6BVaUfNrUBoahIuOVuctdlkYWabmQIRkXVG2pOwAcCEbmVxctmOWIzlLhW
aQGZvebtV/EhRr8ynXVltdccMJFBeSxUHEnv1MEdVlMAYanv1NU1Ndnn7WPHG5NZ
2xOUM2sswZ8HmsT+WeukuU+pLnYXOV/EiCNSEI7DakpMdVKp5c0i5Be9dbIs90AY
Giap6VBeQbOvU6ZoHzF/Xsp0VZHer54CFYS70bm4agkAW+k2cW+DCM5sXPhqDawn
n8oPf6u/Nz9XwLVWQrQZBa5TXWZwY12ku4vpBLkdoEk3yZtLbtpKYACkBjO39gpD
JG1GtQRtrjKYty59RnZeGZuC+JTs+CGo2lLxfRsDqrGPQXkSqIer0PwZ1Ng3Rmt7
GCBPZM4bOm64/05tVrZL8JcK1cISrfwZDQadaFspKrilGg/xY21NiHGHc8DRH2RO
1yXSgAn2NlNH+iAgGF+zqQmdd83PbXVJewVhwCBRdgFXh2G0CeVNfdchx1Een6bm
WiBrEpnjWRJ6Px+kwlqnK1jBam7AKlAby5unBeoeVHEm3mrN92kJ62bGGHFTu/Yf
uYALb3NJFrN+OGlMVwcf/8Bnxx1b+Ggkpmp7dVq5CToVWrg8SatXJSMoes2IenFu
SYMRlg382WTMvshtmDodjBAIVQqgJiFoDpK39X0i/BXQ9D7d6tYBzQTEmfy8jFB3
LkBparLVVAGxGUL4wZ46IlQ22tmcNgT2RkWU7mrkidj3QGJAM0QfdwveVS+oIkPr
65U+1em/ryEgdmCglNvmkeB9CkLjqDxPYL6T11e/piapBUNzlnLxZvNwGKmIzQIy
4hVc9kCnewEaDFTbYBnHFRpO2/NgxLtwRADfDCTmrF7IYiM+J1QIvJB96TXWprPx
nbAjgUJVnxRn6lpLOKjAtby0/AWrmtN1urBX/8lj7wcvoQck/SKfVRlVnRY0TIjD
TmRGHkcja432s6xFmxBdVgQPCCDzJteWVPS/XC0/26WVW0S06BqvOxLK57dVeaMe
PMVcuSM/Z4x4tjJZvoiZu8yWCu+etJpA+XS8yibrTcZw2/Py6soxPpt4NfW4EIPM
6Q+JakuaxA22s34Q/vmYNoe72PBENn1D9SjsY2Yq//PKw7o12PYPjpWxOIkJsk+0
NlL2pVwKEC3NUwTEWPv4Sjy8dmlYbbhci7i1+L5RuWV98AJiPhAr5jIdhV5xEk9/
HNLSn6FMdwgD/VrII2933rszTNqVA/D7w+yN/rsq1f4A6O138CgxCI+RlfF3Y+xt
2WEdqXpGxjuDwCu81q3vl8ZW/bH7tJkIDzNUCiXZ430QoMJLRzeQyK6N/EjrVlRL
N168V1s/KtEhXrK6iBxtd0T1pBjh8OFXustMCp6zojHX984VApGOm+PS92tzvmVs
dwPljx49xbNa5s8XojJ5/epuqmd0gW0WCVKF1aVwRfefH7nThn0hH3fce/buwFNR
ZYOZw1J1xHP4Rs+lVbP+VB4PQfXavAoHsiPIyu5kRijlPZJhCphxstg+bcjfnIRl
D/loRfaIhIJcwovVJa5WODrpPhBD1o8NsvO7Ti0BOhSdunlpL+1KPK0MWZT1r2D6
dTcRL+v+sPBZjWqts52WXDLzroW32L/NxNTIY2zU45c5f+JdS3zaAMiCsbGJd3Yx
Yhd43ex0bkJzdWVSxzHXnTq9QI8RrQtmUVd0/FxqLP1SCMqy8dSHBnRlCw/84cFy
wzX6k077lXliFNVOkzvChh/5yyzqYCx3eZPR3aU3SsvXd5T6rZXPDeYGCKNPYeAO
I9LAFG72ZK4tXc7JIv03/eVBmnB10nHoifta1ZWh576bdmpjCMZlvmkAxOvtGpHV
A2t8O2MILS3qK0mp5eNVDYeg1y1wwV8liEUgC3N0Fpy4ldr4vw1Q3p3AU68RLeNJ
qx9245+3aPSIxJx4EBovWciILJSyKJz1LHfyn2i590exXzj7DJQDf1XeaCl0mwG/
mWJmK9g4V3TS4SY7wzkXzFrpyBEvFXrwJcnLmd1o5sCW9f5AiCGQyU0WL8npBv2i
sQPbLU+hOGXhdRguUAx5Yj4sv7pqniSuc5pAdLRDGP/+sPV9vLJR7HVpYsy5zvc5
YECfrcz1ehT/2T7Fje+34SEcTnxnriJoJo/nQoMsnhIM+QKVYeO8+FonHj1eiNnb
RCYDWGGZw2nVzdN2VoeuFQwVbf/tBaut483lXWexrE22GKsKlHlmyKS2ADi5RGhs
pxrgxk5IFaSXJRR4Ur5oask3dn928ya/pgfaCqhgULJQxWBCfqyCqUXaj7NQsXNC
XOIDL/EqqRL3ix+jK28EZjAjTEcwhCWrUZPk5Om3wHFJ4F5iefaKOXTTy1Vz9q5b
uXC16NaDI7t7+ZYH2NZe7Hg98lxhhdA745bhWZGzhsMf33JQIXmL1Y2UMc3t1Hwp
hkXwbckfl2pKX8u7YJuCDB28Zl+ZoIy2Wa7H7EvAElRCpGeHKrShSS/QYp9Iskt+
QAT5mK8w7Gwl7Uj1dAKnt62xbNIlXjBDrskLb6Sn24mvSts7l7vJpeaSOdBz5JEO
Pi1aiWet8+T3+OSOk0EsPtGpbTFwEpnGQYILl1WIbQfLlYVTIBPvoXTu0detA+i1
HDpZ2Bvky+FX3CvF8KxF6PPa2uJXmcwfnE02Kw/foKPydMtO9SQ2ctvyPqJiNqp9
xwrswHe/ljcqQ9JohR4e8tjTlU3icgihRrkhST7i4GTPK4I+ksVKfVKITyV3/ZlV
ZRxCGdmAddlwI5qZizdhE3/zhXsAHuODNJdU9Ry051wOhPv5Y6bN4tV+ZnzDqK66
Aw4L33vPMq7hX9DTFhoFhRCJ29B4yvqhDpRTNL5tgeJFTGZJKo8AYIcbwLXGEhwn
qQfv0mU71YpxrouTrcoumsIl7Ut+ovjMPZyncbjCPQUmMPzt+1qNFPRghi4OIWkq
7V8h7hoe3TiJ4E0QqG5C/AvAef5hj/rjF3uK4xNyZi9WII7/Nl3ZFiMNf+cNRmKC
cpa/Hg8/KzG6ZL58j+Er0assk0M48eChjE3ALJ65pobrqC8hnhLniGRfGdIyT3r9
dq3UVAP7AFvg3l0i6hGxsvKHXc6cOL4oN0y7u9iXG+GXKs6sDkve5/lqxfFerTpP
smAGJVs3hCH2WhDROxtnnplJiUXr4XYejgUJEEf/jzh9abVuv4rWVwI5Mx82y5h+
PiKE3ciC+pmBsgIzJ3uLWttD3ge9vLnO3Q13YxmRz/zC95JBLCIY6bDM1sC/xWln
WUwUCnLQGYzONzENVEc4TOzTiu3WVZg1fLb7E0HcdhIdvZo5p0GnsdpbJTU0PZPn
qXLOf4e/ag+SIXDe/CwrKsMhq2c0fvNVvwIS3Jv4KZ/4pCOjJe7C62MLo2UoitGM
ks58Lp13D55pJ8Glw7xVJWCS/b2DfNWgjNnqWKC3aL1tppwKO/MmpdNjZajdtLsh
RZsQsGWnFY5QdqCydG3DBXeJGt52Mp54jVYhxn2RMurLATle3mhyIzdy2lCqSq9N
gKkrwSu/jgAIiKi4SYjW0qWWUZLayv5/N75doJf5+8s8INL0Sjxbq4aubrT6USKT
6N9X+7+pNUS6C4CpjTbfHk95Sz1KV7w0vt9EBe7TBMWqP+FhL2L9ZFlQCJLQY0zd
N53EQnXb+u0AP5l8eAbH1QQLliiYTG4Rv5POYtaIqdBgwNOA9ut7wMisof+BXK84
6M6lgiFLOcLg+iOTC9/XSM5EadUZEqGEqoikLhzYngXVOIU4fZ2biKgow6LBpg1o
la3fLQ4s/HYaqWm8XSOijmFdbCKW03x51ji4XVUA4N10LdcryuJNrnlXi48xYNci
DRyGW9iljnLRLIpLC4e6wd989s1NKPoakG1I6KaZ4/jMDoNP7lo5gcSl+zKdD5T7
q9lLAC3AR9F8eCDx1y/pf3OWe9Ffrf3XH+O+ltZcaLQY6RQ6F9XEPTZoHZahYFju
LIic0SyM/a3Pg6JhdbCgKZi9iEQT37thVfKXEQ9PwntOvkyDuLAPac4IGK7tmnUv
Kq9cpdtN35QFtt8LxkElKlr2HexEw3yaSr3wMXhfCN/jkSAX//LrVwlHvECG8VHN
PWPiTLusmtaZu5UZjAc6rq1bOPj6io6QnnaAVteHnd9XKzMvtE49nE4z3uHPQUp3
G4+xhG0mxT6NpkA8TmjJ77hXSrkNVpMpR+tLGHB0DhpdYt9Fd/MquZDlNkECO1tM
+vEMbD7+DZ0CfmrUwbwqJMxzDe6+xcSqJIHBmgqJHw7JX8emxMYQkXGpVScrM80b
3cL7u9HRXXowyCLgON6TCEPWN8NUQU3gtjETERNcroVEugak7tJh6INI3oOcPHgy
j8rpqQrA2Q9tNTBhMJU+9OPCzM5mPLiB0gKiP57woaV9tTG5/NkyLFIJuLHhbpGE
3vMDMOPez7MBD93TC0mb4PRWnlAne3lx4RIHQdxiPNnIZ4IcxMqQgHtaYS3jLP3S
GDSaEVaXh+WBRwIF/RIDHXeG7ERD85CuhQNqOxyU/lH9n/f8nswnuKocOPROUqVG
AD1q7kTVTziWKQJj7yED2nDviiFGdroM2p5m7JT3XqIusnmZxU2G4wMdkTWqosU5
RNu1JWjN70Rhl8Ikc71HPlMSgf9YEy4V7O3i2f+bO9G1XXHSklmClse8PuW8C7QQ
o5aeDl29NeZ+k3uGj5o8PitqwTMIiI1fW2umaVDular9tuaKXE8SUkPRt+tqZZax
TtRz9kFecyvGb6l0crxJ9/+rKSPt4lCV65uEig04Rpx1L14ypfrEzLEFtvEoUPOM
5Ipuwiu+uPEGDoU5J7ZRg+afvNeYTZoGdGdkEva1A1F3g2tEwDy/a3cIu4PfeeJd
YczpENNBWPWS7EYn85Gm7Y3eY6T3RylOh2i2hsphhPxPl3rrJ0pjE1Mq1s6u8Y0n
WJJ5EPr1e5wUUMhUBjNQk8ZBnpcMtPse5TnVpmLAaiyE2j1MCYJQNgVyysSDmaRW
Ff6YzZBDgNKfewSRKTBbUQ==
`pragma protect end_protected
