// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:27 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XAUULrUeuWV546lNG4HbffzWzYOw8+6aAbYJT0dILBCiiZrB6yxPFKM2lha4QyjN
+XLh1LWjWhS2mz4hxntwJBYHC63ODleWoKZT3vZp3eYdUU3kyl70n8V7k6UicJsf
+HZ7ksfAKKFPiL/GZQcyzpVaX2fxP7eky0KYCK/Ogsw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46192)
HpHay3+oHC15BjCBxQEAXvXZyPB8VrpwMzrJhEB1tnILHR7rlLaJVRCGrKJgZ3UF
2jq1ySQp7nrOubxiW+y5yt6iqsh51BDqJssPpw27yrNXhdURHUak0OU6VAhPa0Pd
TuvqV1dKQ5W7Ojhc+YSWdw73CDsjbq1ZRpoZOz2SeU4Dkz2fXHgSwK4JHUIthtaS
/c9Z39FHMLwBmeqbvBXWkzbBvoJKVd7W2LvC6nMDz126VA7BcZH4Kf2NrRX0W+IK
hXlUyKH7/37GsA427EJiEm310e40ZyTdf7a5Q5Ue0qXy2/0pRihgbqIjsxGyT1Hh
eHyTU+ehp9YrmXO3oxDiVdCHAK2gf8ZFacKDy5RhBqRfp3ilLqmNWQWBaYJ9LRIV
iT2UCyH7DoLThal+PGZkwtnmOTXuBgYxgszfYKipFqGBuVzQXjmzsUF9P8rf1J95
YOaHPPIV7x/9LIWiCJjXTePoWTP9A5WdOF+cXOR3u8Yg5npijBTfW891urQPB610
dGpfgrY6KCg0zjir7+Zk448zgBqygub8RePpGL4llaAmYKn6fA3edCyUuBIBN/C0
p+DkX1DkwAHEuovPfUE/9bC712KHYwJLmHhrYgGcTMovCEIroIaAe+iSk9I3D134
1VoD2fRwjwgp4XKqzJiX8WlvpnP8BtE9q2c8lxEUrPDW7jYtOXID+ybPzXnC5yZe
/DHS/23KFwtfXufzD3K5SWgrJbwMPjOkIPy6tVRyi6FmVJ8+jakzCSsJBytlN/Kx
OAAwxigSSctZOhSDalujXiUpvwzCov54g3O7WGtq1x3gA3lKbeeDMm0tlI38iF0S
RS9QX4PDQwK2nlZIXzxEoHwH1ihkDGQgWrGjxSmD9efvQVLEZbusBQmF0NbURAsT
PnzjQZObtRf0c/CybQ2uTHBjCrcRKH8lc/+tVxpZA8OF6iuIq2+sXAKKag5p8L/Q
HtQXNJQh+P1jS2CjpGJR8AZe6KvAOtch+AT5w3pSz6zNWitE/rXWB4OEk2KWRfOz
htD8tCeGG2lUbH/xnAXG3pFhzAvpkaOi/2Oq2UzTR64JbOW1a5/Dv4fjqphW9RPr
TfRv6mWX5bWVTTnXb0su3F5a7ld2/z/S46ubKPBO3/EUjdLUImTD7XSRxmopdLdE
WfANGmGx/49R8oGfDhubodEmGd3CiH0GY5w3p6vXeebik3A1WYLKVyhf49AXwbvP
E1D0FPRXOBvDK8A8Zq9L4J+kKpxgHTDuy3mlpw1JKLORAwleFGnMCqyXbrjI9KrJ
/r5XyZXFvLQ4jZWdSK0f2jnuzFU8cf/EGQPCFqVSpRqHha37Bi02qXYc8rvaSdDt
ZHrA8ytZywwI4FFggLuiv51WgGc58Paslu/3SRhhi7rL50abN7hf/ofc7Iv6+0Ej
5Hea0Nu8bAzBAqYMuczrI69YBsvXrg4FgSZ+3ucYIqc1b4lZ1APnEKM/iz4eIRXd
O5EvDAbIAQGNoX83jry8fZrmZrU78ufXGntMgHZVBkjwbBy18+eEqLSEvrC/tmGO
JIKOrvEmFmheiKVEoQKy96Pd5GLjbZGNtLuYdj5TjVEpfP6XCqc8J00iRgDc3OWQ
I1ZCoaqjmXFufOy6qcMFhXQIxZcfna2O1V38VbZ3WSGGAhYa+FZNKGEV9PrenewS
QUGOnKIjL3Z+E6DjJ7qIxCtxYlfPCmxP6J5FUSukeOG4Ov4D30dTykAYWI1w1krm
wyEaxx66UxAQeDVpow2p2Iq27WeM75k5f6GdvfkDcvq9ABiNCsrkBk9AjLAjTD15
47eiH1K9XiiZtAiBNSwj9dud5usaaKPxnIaTfKQ5Z+xUgey5z1Agua3GxjEF4HOy
IqN5BPARJD9xYP8kKg6ELPc9esqGxJ0qHhXaZF4YpXHtBu4+g5lf6QKtjOh/jSGL
dzHJQBLaNbjqQZcfJyAHyNcRoVfhUuaMYmYBCkB7cE7eWDlF4DTW7DMcnvihb3CJ
qbMjcRcLnZHhUjqywlgzE/LZJeT3aLVwwdjMtwbEmuZjrmhoJQKJq/gAoXtkb3p4
Or0im7xAXjNcQU7OlqwIIv+fHi5INlDHDwuCLeXLkNyWUG40iqOcS+dZYjrvT3jj
c3Z1rKYk5EvPRHzeIGtjmEiyR+20bk++9EGzuBBouCQA4UFwxiBbiFYJZqp8NgCe
SCzkjY8k2A4seFvgrQhkrO7rZQRv4mxUEe8JpXIMgJUAl0jdY7+PaUhM49YEEZor
YKzP+ddcUaMGmwGaOFE0WeUpGR0UYj+sgcb1CM8PJC4X1+ug9SuF31UC4amEACWE
L5JrNn91BM98+lXKytYFwQInGIVCRAKFDMeVrOELXDDnRHBjw+PwzbriLAhkucZs
hYckteaXvgfZItTbHaM+cr0WW+idhQpIoyAYIPmfrJy0VJgM03nGwg2Bz1VVIgzV
051ZQi4sLQDPhhQAowT9GpfbaSWlEYQI8fit8wZYYbKeDSab61tyA1AD9Q4ViZH4
mfGJxomJEXzK46qnhSACEhHmZKTOTdPQenFV9T3OSuG3I3cd8UdfdyieKP6RYjDA
5T5XE3A7KJwa7RzLO/CvNrPUK9Y0rVhZ18bAhpB5GyK6vPYrIK6apNFJWjL9SdAx
3bhnuM5cGPy6RgoELTNjcGYx6QRZTa6lx12mHtIrREezTNlryYAC3AMp/Z0MFxVc
XgDVzzrNDWUFaMm7j3Z3DaV7UKrT3U2tqQQJhy3TK4MeC2dB4CSagCBoV5VRgY79
TSNVZty30FTM0t9ezxbL46YfLRQ86cSpj71BZcR/4Qya7wnijyByT56hnA7eQ+lj
p+WstDnhs6Kqe4MNO2X0W1dZQqu+3ci7PAV2vMp2IJCa399BtDQBQEWYK7mwwymw
YuDgaGq2w6/Qyu3eEYUhacsJx7LtNccu66uMCsQA56m08q5JZbfCxcmeaTl5u+3N
a58oCr6YjAVOTeVdMBVgFOeb15EK5UVhVaAsou+wG8SpmqQDH95PJ2OcMNTvxe4d
RY1/6iA4eh4uX004U3haB1ph1q6LLnESl0YeNYFSvOwkZIPNls2qyniuxlFJyr57
FtsVnoBljeN1PAasM0D1arLpdo753S0Ld34BOABq4lPZFq4B8yWug7gCvexTURJO
NSJfkwesDVsdZoV7J498IPHmhc9Mf8eUsxvOndNRG43WSYmx+PieLgKYE8ijpjxq
lbH+tykrPNVsq2SmJNd0jK3KIYmYXrHwSSQOA1SHTT9kqJzoTT4/fFrO0y7KY3UY
vk3+FxuUV3HLAlMpN3iT4kbKovrZ8PiJg+07jJ5ZO8tj6scbK/SxMRXFIaqd1mjZ
j1PY1BF9jELfvk/BahJHbp9AQCPYiMI1xAa+zJZ925VQ9BycPGGtLT6rJQhlKZKJ
hESA2XvtdzJZ6f2xTI2TZ19xyjNOReO0wQqr6W2uP8SGbynYeX9+9q28gckTqB+R
zpLXjryRHGYTJM+EVF9GkcUPsCq3bgvs6PcLValLeDTOsQhRKQDBwcfhwyX9u6Ig
N/atCT/nDBdEc5CvBY4e0WiGopgc5EjKKDj0ytQcvBm/2unnAYKUIpXs1+83SSbt
8EsFDj1XdLuKPkzknpiiw1qdfqYN1HPKcEWvYyaWwopT56EVrnhYDNdkHuRqx0/v
nhpmL/6Opd8yEnPVSTxHobarCZb5J5Juay8wxIBbAl10onqU8Ws1xuWMCxt740xs
uSlBseXsVAPFIf0Rtj6BhlUp5bXzG2x0dJekwPwIYtQVdfHraBdTIhI6rHcxl+xs
VQ7aeEWvPRgDgFyzZzDx7zQb63wxjUmRpFw3Z1Jn6PPGeSOkhmnGQNYjXDHidYes
Kbg2lOFF9MhIO/pjOH6qFznTtMFp8gUkwr3STO1F/nkD5Eg5TKl4MVHvQbCtcBmd
y0tMQOdlftAouDD3PO/Jy6YygiGkmrWTI1HgEiOzQfzjNSvsaMUIfZm77F3KXnhI
leMZ2PYNnF8b/eKPurNqUiEFsOf7kbssTMt1yHOK2cQ2jjru85Nk62oqVuDu6pjN
aaCGJfexj9PRJRkp/NdD5wiQuYPHuffC0NGpXtfcgoOQc7XLUnNdzktkXLDJjsJi
Kqripw10qbQ9/Lyu6SZZkuNXRL/dBf2tIrViKmW8fJL4/NBz8OJm9g3qcd9EHFz4
RvN5thfxXvlS6hHmYm5s6NPWMYt1d4FpJBJEicGjFmyAdMYH+B+ddiDsRBSwbNFx
cre5yNmeJbmzd2dzrRbujjuYHnppPOeTU4lBBGIxCHU0llG8i9bcKGq1Cg2HXOYq
i0x1nN4qi8xba7F/5uTTLcpNgtui0AslP1GzrkkrxXrkJQoKvqj2zi4eiLuz2JYs
C8AwM5Yi/1s3xDR8pjjJ/d421mTkFCMf+luFnVZNtyZLZepfKUtS3z6QPfEon7gp
0pvdGaPmGS8P4i/46NzXIiK2v/qA8tIP5PPJ+R6cgqvdMJ+Z0JFWvf+FvIQ3tC6y
8/gj7ZkNnxzxgMi+1Ri+vazEjlrXUquPBCrjOFuyw/qqj1KOdVDRTQLYdpcZxmEA
jhGMJUPe1FFmDEUggd1hEgt+MZvVg4U/ufcF3+hlI5a+kDFIXXP84vVYZuWIgtQQ
NKsBNZ+PEuWaStPdAyTGpjoorD5KauYEl9O2Xc8TzgJ3DttFPTs2uBHoBVcspV3P
6H8ANj9ZW1vnMmIJcZMR6Y0TyU7/8kZ849Qdl0NK+21oMXkjQPCWFmNkE0ljPR69
Jrmint5k4a0xr9v0V5EGrGNxjCFuMeLT2FpE6k/9jTvzDVLGM3CQJN7+XIJzC8rI
N3sPFCGklDewYw7/ZIGt01DsbP+cAe4RsBE5BJTQTvw+K5wkIvaT9m1+Ke3JHwLx
j3BvksXTW/d5+0VAx9ffKKm6gnLyQn3KTK7hKZqYRckshNeRk5l+YMd+XEVz062T
kU/UEfovIZMdKdt+V6zTSALuhukQTcGa6JcYG3SZwO/6whwz51YoxcI+79XVpm8b
D4pu0EeQKlPEGc1wHXbP8SFDZq/aNwfaNr8dbbVm/y0TdfNnt6l8TKMEBgStI0Ij
Xhk3fd73aIdM4kgRYVc4oojSO6jwUXTrwci5LVa4yjc44rh3asFNCU8o9UQQJ3Ih
ERqevdjC7ksEpdDf38P+TvMNp9M6RJa9U78v3kHTknNinEa7sHNdscRagBTZezEl
x9H0wxBIbF6Nf+iHmfqNAmyTiJbcV+As94D25fKVs3nE/lTUkZ1cOEFlS8s1cXpZ
Z/J9vp5qLflND+awxdZ0jUhI6Ymt7uQln5eczfQkKmG04ykcusHdK6RwJTZjwB2R
2ViSy+h8SPQyXYdRUa769mIHKyd81a30o+95YYxv5Yv8pF9b3yCGI+HIGxTL8762
WgeXKE5y7W898wjntgolj9sqNb7tdpp8gOGk1Gu0o4BxDXUBrA5KEI8+SXbhAJBq
9qrRVCqpTJIHyV99HoohaJ7TtjSYH5FvCO8mBXryEZuzdUr2wdV7w92JL2mFJq4M
7D4qPYE6ieLfNhcVW/WHzpAMXOn6TwO9we2vklqbTeOgLL17IU41T9uPHXqX+ApC
jr1POAFFOvDmG8FsorZxBhwNvhrSAfNOJ+2A4V9FE4fYunZs+MZEEiydsrGNeUHK
/iWvoxEp7Ow+Ld3PsOJmY/gllMRrIZKeWlCSh0n8RG8JMRgI6TFhf3D8j3yi41sK
b8yVMvK87fmRj0wJwBOFS3ZaoiGmHwZNWABm5EvZ8qPVTs03HCDIe7fQIOkBYQSp
5cQnUXLQlbJ6ofx5lSnTCAhaGqvCvZb1YYMsK1NHK4Yja2jxeXqZ65MRz4hybxCA
085K53WcQttdF4IDQXirSAj9YZiK83hz3g02jaUnO+KIjlJrWSiuteVzZB2gv85g
NKSAcvG8H7xcmzi9EnovYl49fvGVwpmD9T2lhr4kkLjQdN6HdbhLsO0bqaAWmrgx
LB9SZYY7AMEgKAclrAa0zSZ+FIYd3chtpSpIdE2y1mC4EP7H7RAXtZzyNHwA4otS
kVqxvXWjR4pNmixrTD1RtAEecXxoBLQYXykUfFl/Yqw9czUbc2n0TFlUSnJusBU1
Kq7UZG3GIJtA0c/UT6Cgf3G0ogTI4SrI9wsoYBZEt4L0HHZTIB4pZv1YAvUYV0gq
H3FsDEIHSsCFtzrSxWzEdj8FkpP3mX9L2BHPCPuGYQz64lTI6p9JLgQukhuSqzIO
ZzpaA44cap++Rr/dHhS97cYmTEdjKM6kRml3hZB3nv4aDH0EKpU/FS+GgfdxhTF6
ttgXOcQRA6ASVDPcWoe4pEiZDjJD3QVoGmLZnHPv9mfwpdC0k9GQRHIZdIemQ2Qy
x9do3D0Tw6tfm9iwhTyFEuygDpJIcueoGvvaDKa9DY8/cbVw9hKP/h1uzTPMwxle
ORkrDgb0QAtMHKJaEFjiXeq8QnUYTLmTcFi2QWPXac9JmecGGRVSeOjmg49+g98R
tQ8txdqbSyDP9uPxwmBZNM36Z81ltReZ/MquN+c5ztgJIiy3CbhEBABq9Vbin7zo
6GuqDhLBMms/m3mSKUPHqAnFp2WBD188GDT5odTNrhOLi9MvNFiNVne7ZSORzEjM
bh0lkLqUzu23jpbfimJq0LNsMrulT8g6Htkq09l85SiuvmXrb84NuVZdlirfdETA
D5JTe9vlm/XspcSqxCNMCjVO5cMI4F52f//PsHuW//1JybliNkrFuVi8g9FAHTrw
EsGr1nc8ox6DMVas/JCjbZRfHLMa3fTiNMbt87V5MNguy9XetcvCS8B/ifGEB6bT
SCypFTqvVntEspt5p1I2eJPCzunxIfpM12FBqcTtgQ0NYSTZuOeVQaMH8eqnslV7
qL7mu6GP05hsmOjoy+HRFa4srlrEhSt5RVkqxw5dcKWGpi3vhKYRmZYqT/8EYohR
C+BGzJMWuJBYED4MQByV3ai0QHjMZafD3uBQaq5cpWmahGhdV5WQd7RbMBYkeNfa
9sbaDmLWiiHbNmxSJ8H8CJWuLWHekV/5tQ5N6dYm6HV9okmxEQ8W0iMjMcKUvZcj
n8XG+vaBqxx22sXDUlZhj559KhTUo+bMC/HVpB9ZResMSC+zLvVZEYWJgLMqtCZy
ydbEJD2iosoPo6MdfVtmkTVg2GWuTBTvBXnQbOVJ5WyXADUPyVRBBOMRzvBEIAUh
NDQWhMTUzsbPxfigLh/Ikg/EPP3cOFW90r/iMqx+88eA6CYHN7AkQQ1CTz02Ay5a
iWi3HRw82Zpl53YrJfDdQ592Xb1Kt5An0uPprx1A7nS570FrDmsr2/RjF9kqITcB
XfuxlpsV4/vZFayHWe7WKiIBOCr4gA451bpiV53Qe11nO2AMjJoWco1FIV4pl9sZ
r+SCV/I2gAWuNNuBQ+sUkODti75L7Rl0/ChUqr4X1yRhw7nZAQiRVL8vRUfimak3
Ndbfp1RS/hJ6OhbxbVbi9dkwoQcTUpI5CjYZYNDgetdJqaedSQ76hI1uVt+xfB5G
a3mHURIB6MBiDpmOMTde2m5yYVrzp/fgMgWuQrszd5Zbybyhni1RmepqTOeSOMq3
4EEkbeAgB2rUyLsXFkCUQMFUG5p/gVmzKbjQ0dMHLHOz19ecbvZLym0+B2Rnk755
FnTE5yiSssyi3y33ILHvGPE9CW3m5BAu8stp0yuaqriXYmG6sLtavubYtCSGMLfD
DAgdDZye2paFsnj4HNrjDsiPxWPGPWYZBx40deTDhwVDWV9jOy5byX9u8u3XKxMQ
BdhGboV+7ney2ShcP4tQZ0EvduE+c5jzFEkcPi+EILMhi9Zi6V75OtlhXk6CKp6Y
kyLA8/jkV5d2rFlXoaK/wGrZIanRVbx6mwg5Y0JKlMuSttzrlY2HRbNK1aeIFLfk
ZRhb4hCgt8fbbmIL8RYuTmolvpfmoQPkmEQlZQ19jmxMTfastsK3bseiEZZfRJZs
u8KcQsZ10mGQkmY3XjNVq6hFVliYnAnz+HVXNkpHmcHWy75Oqdpl8rzWHUt+Cg8+
BAkee5dOnpimtzMN5ShPo7InCktUHoCuSgNlt9HXvLE1woEdrna4qa51cqhFyxFW
8IyRZOoac+6CNnNfzz+2Va1MrtXToajFfuWum1jeqTzN11AH5OECnvAAGCh8xdur
HvGsMBdJRINS85DpWqjc8fcY/Gwhe84dfJtmr4LZgaN2Qg3kcAAQVTmFz9qXXLAC
dS6zkVniWr7PMbr8S2W6ih8j6g6dzJ//ZMqUStFWHCbx2N0XLb2+vEZLjWl99tc0
8g9vEn/G89uHBCEJKJ5DNY4tZx0yUPPfVGsZ3uUhoWLklCihOywexiumh/HEnEMn
y6V3X9ufhZsu8bLDyNqGDttm6pS56qtR+kib+OCImbWKBea9Z+ErJeuOx9qMGjge
lkvSY8fagHYaIyk4t3U40BnetHIItPcmKHg0qZxTHmrf2v/W+SEX49LWwogwati+
KZLQFm8zRVgpHoB5PuAnU5hPxVAkWijNPNOPLmxKlL2Qe0U3WIUJWq9XmL+IPQe8
ipqWv5450Oh5IP+xud9yIyOp/tfidnxrvYbnLnCW4iiAmRvR/o2Wvt3uBRLbandU
DYSlHvik76ng9myZ1I5bGMRuMyQ3r+YwWCaRlyvrPx4IRWRZU3Z36ZrvAUjHS7nN
VU1jOhgrEOn0KcWVLx5jtipXjs492Sq1F84xUewtFpmgZxNI5rm+MNqkjDFTA8lx
+Oy3SpD3Pd7EdtT/ugSDYwXEqzXMSrhJnuBjhkzh5KUEA8y5SU3ONXUTVpy9SUTg
NUWac+EAcDpOT0690ziUbP0/LGeyHKZ+CgQsFLYMJKLkI17kQv2a+o9D2/x64Ck2
qjuO2me4JL7tV8iCK2/w3gETCrp6ARO5hX6O0RgRDq5ZicCOszOzbgxKpZ+OXTXb
I4OjX/WB68kGiX4SZRbNUKLsoStCnpaTg62MZfa3GzshTpfHX+TNacnzILMGjc8N
A9M5v8XhTvCfh4mNT3e0prMz3F4cKXix/T2QxwC0rlq6DdAw+FW27ULE05gWbQBT
kSUVsI/V8XDTXJh50kHTDkbZrZmNWJxEBnAepvqGPtW2HALAYYGu+R7UENVsqxKQ
iJcWa/VI1YpXPJSVU5WcRiJK3tIaVo2uani3tvpasTgfbobIidAcIlqCo7lR+NH+
0UrnFXbIMGaRrjPCSp7uGd2klNsufLhyDifEGCSq34XDdknzZsrep/pwZ07ag+O7
EIExveTV1iS+N5YyWebccN0oyM21MVCXHHiL/D/F23KqikT3LqoJ60m+U6jacLgh
3IQd/kntb1JCJ2R4c0NaIe0EF0+hKbiXghscF6yeaN12Ji5JntkeOB8gqsCcQdgT
+lyt1JaYOlD3U05g9Wvte3Xs3ol6GqOsdnAt5B3J8k6M0nYu9ADNiTtu80jqFaTA
KVoj66Jr0pfdpej1Lg5ctXji0JpcLDAoOmK09rJ5CIZpKvgV04KxpAdPozIpzMDP
jSMiDPMl8hxTrGDlQbtJM7zKLHDk/VyeyDkgg9QQHdcvR8O/NVx3DEbLM5ZA6BBm
oeTeO1qSEiHXP2UJbteveyCKsoMK4qIuckZZBI4tJlRzV89AXxgZgC48o5W+jiyi
nY2QU71nffQGn49iwxC5KY0RbYXXfdFq6yL88DEPAQpJbSOrZHzzCGVg1xV33D2J
fcpKNoTxRidDzGHYVvEl74Qwns8xNh1rSGehE1tDQ6X3usvRQNEJnhUECQ6dfGfR
gEKdXSDmtJPVuvBWaniZ5fNOc8u06XvvCg+5XRIUBTjOt72xC9TSU4bsK3OBhNz0
4z1R6LO1YG3Jifwmffat7wjXYRqXA47H44Ww271pReDTH4VFcVAyeQfG0l0GmyAn
zE8SBJJDsTqwKZ5rtCaxag/ZqLU5Zp6vSoZHSp1HlYBTSSPMhihLirkL4zhUZesR
UruUHjyhzv9E/oMS91CcPhxm8b3wueBNyngpGcjKl5PFP6c5HmRVT9gW9ikI15yF
jXM3oF71ogNlK3j6CqDr393qdXKu7XkMX/1vEF82MCsSzVZzMZxw784tafAqF9Mp
yobHoF77vMElJn+5gUBe3uMCmag/cn96EDjp6ey9fuw/QWxxtOMQyZvOKB5d0UIg
CbPPEZHBjZJYhBvbzeHyNTV3iOZXhF3lJNwTal8dsam/TZcLmMr/flMWKpPetAEe
VqDMuxS04BtfMcK7ptJV1xc9Ps2nFhtGEdtr1Iyu6ywhogX8M8iAtd52mWU0fLt7
is749LRH6WOj9mR9MchqDEBKnz5xs47XZs5WQ3vfuv1/Mmhoq+KuVd2VpQK62r2U
SWBWnW2yuqV2VJXtyySEm3O/efCqY3e7xcynB350Ci0z8YSS3at3OK0w1Gitc+GQ
pKFukh4uihyE/3VTLS+aRNArk4nCkRzTwvrDU2TYzZm4BBl+yZ7vGKJ14BnFkhC0
yoW9tHkZDr0mZ10KCbl7eXLDf/bNjAmWudIgiEvcFxl51sd+fXeGgZPLYkWUrxtC
+RpKR7iNG3V/3dxAODvJEl96mKfso2oD9pJud7NLXcpgN9QTVPiw5C7xosDz+Fb7
JVh+pBUQRBnFyy2DPiUfGwIj7U4gBGfv2REy5UbeATOyThKrP6I1DeA72mSwYbtU
cjFnU8hbsCxd4o+Fie+Yg5s+AEtwTtQaENKVyMLMwx6sqByR+LovnvqxKRwKM0Qy
P5vD3MO4lPkbq9gF3UxK5wESA2Ilg9Kas3PV4cqh0+XmsE3NXBnqL5zV3Hfe/PD0
D072Y8wQYHNRJk0j4nO7qCEv6faXnkS1rrzllohIgu8/odYtlgwjwUKuo+6IdUTr
AH866doA15ztQNI3O23FRE+6JqAceBQ/CRYCDnMc7x2zzkdLo49uETEUmL/cZJIC
uKIFNiEDq58jwG5oU4gZOJmIFDs28g/W8n3GPk8MwuX8iUafhp5ltPgKTvFrjlpH
Pj86/+HGrixr60vKQxr9QteP6Mi8NHeKmRAIk0TP5xhjZfHwb+CU4HvZC8RkYojt
rTfzBDyNxwZ7LZVJ5Nulxq2vhC5pOJVCtU9FGNOdMsb5lN0sYGryJH0NPBXJhX6r
RgdRQIxdUyN7OidTyXfzxRbqXSOJWXiDZP0OomPc66F03jjUieG1c7OKOU68ZqUH
N2JLdtNHa+vOi1vdN+NeSGgLc79qWq4BtHZHJb/XCiVd55b6ZAhBGA73V13+fuCg
6UHxVOX6QPPSEsvUX5pp8VeVESDL4Ex7JR/SFXI816bC37tdprskDB6j0Oi560kk
v007atLq8DuJbcdsfO0ohoXcRqQOWYET7lBcdMPcQTBdFkTYe541vmDacRYPG9HH
oA09dpvkp5kFNya/y+e7RBUA4yS6JOxzjEJRDOPSpmL3y3YMBVOeiKvC2SaAM0L2
sUq42jxyJ25JjTbuPJVwVBH1aMZXn2zoQ3GJGnn0d8biOic3tI5hHltC86kinNYz
+0CgP8Bwy9oWOyvDjmoTC0q5/QdYdl0uPG8tHxNWR/jM8OaQJM8mbY47yELZVslm
YuO0HxURG1CC3MAeeB5e9cbampAal+lbBmzhfxebe55a9fWK8a7HaQM9+lRb0ZlK
KGTisBYudXWpptr11sLJSp5flMlVEjZedc/zFnHUZjWe3k9ooevM/jfirN+MnmlI
kmZhZj9a3Ob5dKfQkY5R1rr/zeqo0P03wFyW8vWTX4w3q+FFEsbguL9h7K+h1VOH
H5irS8AFkXeywGC/Szo200yiBSSLufBN/jl6XrWk5+DLv/QuL153f25gX5S5K5M4
Hnp2qhxGhvK9DisoWlioB5My2jjVLVBzMbuZi3myptRCPhoa2o6q6CncW6mV4ZjF
jCadWa+JqIVuljQgkvitaKlg0HISXoRE/eyGydPWPy3ExVhGAhoeOvdEn+Mo/fyY
HqPK0hZSXYbEpK9OoJMuiXS73o/Thc1awj+bkucOq0JSl24QjbVioYCp1yKt2goM
1CXz88j9CWqNvvlUqgAsSGPCFB/2CIrJBaYR9j0NH918VbCRppDUW1qe3XVTJmCb
b80t5j4jj5DkH5Td3VpMcAUOfn+pmvN569NrM+QVYX3PYxlSwqVbfkY4ujHhYynV
UUKOy1RypqKbaVC542oevElFlTf049WhLi+9opQJP9mSgg52AJsDlSkvZcPSa5ei
1qvsUcJxZIHrPgM31NhX6DPi406FAdwWhM7uu2XqFluZXYes5bBH3YkU4JR0pG2h
/XRW5qGnBfa+JAk8rFo8jKkTxoQuvkye3WIjexHJwuLkZeqp4O1j5DLsnq+cmzlg
UED/FUNbJWvNKnaKUyDZihMlVzniWO6wChLEWoqse2bxE2paCjtrtstcvrg8s8qN
psj44Hyuid85LalZH8Yk5fzejlL8Sutx24JxwjP326unid7rOq2iZq1Bdscpmlna
vHE5fCzsLJ8ZVFtdh0NcwRvuT1mePnk3M5kA1nQ6yIodBBXbOwq2zOnxf/gksAto
aUda/615khMZDva6pX8QmVIkzDmfa+Fq2iY4ULlnj1peP23hWQYB90B4RGCcqgNq
k90QM/hGe8HznjbH/vgLEWd3ZL3DXDOcbQG29e0OgXoPlOiTBIQ9jQKQQ/1b8uzi
5qvopTOQKgOrL2WZ/419owNxnScW1LnEADPwTiQDiIIrQ4gCoKFW9J956Xpctp+Q
MtASQvhJ7StgtF3dV3CayyLzOWtIAa0YGlBQ5MeFQUTKfZcGasJ6b8VorJQdbJN+
0lsp+Uyn/FmpuCpZqh29eVaeAnbA2c6qJ6CfAkDD0vCrRjoC73ROBW7xrnFilseb
ZDsXZ76kg/YUZUsGqbamr7PIT96WOlvOtY+AAERovmlCpnifPJdAEtpS4zKirKd8
JBA4h1197WqE4J+pYF0qfGtxv4dHtBkCWQqyUW7MYutSnJP/9f02HrzYIEizNgOk
+NZrv277kD1tL4BRw6/4e+EatusehKpzEIlJTaZclCnaERgyFWSPGW0XvuLIaCGt
TikfQYmj6y54nZHcqFKhi1qabvkZzl0X3i/fH2jofyUZacEge+UlhNMPvGiK6ytK
D5tnNjbtz9xVxfByL6SxbmnxJ84WivMaH6d71gyoSwfVwWan0tjEb7qn3tQbPBsp
jAzhRVky0HmkYTVMWvJcVRp7/s2Dlx1AMYYQojGb/ef1e6tDkeFL+fcIYAbGhkpC
cWkE0iC+lpnTuyzfmTtAcO8XGcc46Jz2FMGUOeyc051iN2cjEbwmaOpZxRQdvMcv
hggHNVHUQ2iSDz0kOQebLAAPeD4KWuf/8m0idQoe8c6kLY9CX8bVaUxSH3KoVG0w
MGVjSYLG4NPn8WLAfBRQpq1uqSBqh55VX3VhJLSyH2SVgwgsdM3IP//sLxj9cLb7
ZHC+bErUEH0AX8p30Sk5i9c53T5CMOnEAY7tbtvVmS3qL4b4aWNmUc+BtPY101qS
NNrjGbF8mwMemlNYQPegG/Btv1hr3bxEKvEegiaZLWT7kCI90T0FnFAeMmr6dqm3
UW74JN5WFOlPXG9CTaZKAvHA4V6GmcWtBziyI/W3YyedwEvLjegi09KYDKLpHyms
+AvzVvyd29LK/F+lVy6RGifFhQYQRLwOHUxQ8BJm48gG6MCxPtdlBYth0LdVjJG2
v2bFUUEoToeUL2Hi9uVupB/L7BytZYK7nn3n6g8ZF8VzbbWe7PpV4BCLupReiC4t
k2r/QTCNIoWAGCGLi6Qs1wfRos4t8CsdFOca+7w3wK8cZlbFvCOWjk0zvW9k/jeq
TX8Dsd+OIn7y/mnTzsqo13VrKognIH2lf3Fy1HBq4QN5T1XDspBc0HLUo7N5O9HW
6SXAihQzTOVZRZz5RyZQrplcp1kylt2mkupm3Pta0fG2f2j8z3c1IpHZxsVuaQTv
6XRAZxAxw7wYf8/+IXi/lj3UZEVuUj/oFfsIyOC6gG+NRs4fCdOxOB8O5p8T6S+3
/NWX8QCEmknfd0x65Oe4oRH/xjXt3U2H5g2z8iIwscFjqIKiN6N1edNBHXck0XFu
Xg9T3gQ5hGCj9w7++kWZ2+RjLXQIW1Td9Gucrm4xE68LTIMuWowapHsKB1/B8fpD
IBn/f02HhLmdLYvuaMXGCiv7AatQN9fbOA4KbhmldYTurEEnRo8BeYPUiWEkUJnJ
Tt6F23RCYG65Ip1qLoVNkPSIPM5oOw3n/SWaY/wldSUm6XgpTvsmWeknHe1ZYaUS
IrUL4d4VWv2/UTrcS+ceLtoul65N91uDYkhpAoU/7A2WPhIBY4LwR0xS0EhX85gi
9kvm6sxJNnzkzrFhntCedTRTRa8EGsbJLfwEdPAoApA5tsXtUzc/B8K0b8wjSLVr
eMKOm/+gIUjWQ4KaHHlKZQGe+dT62NLq3g0rhBeI9KBhGwu+itzDkH6kf1WNU3sD
iZb4rB1mYqKrjWR2N+/a4RLbiTD7GIqFZXB2BbIzkuzR2k2UTH1Mhr4kvezgHhaz
ke1eIG6QJ36RM3ZdopT11Cmh6tiiWz1/SNyOxTsLqWFkYi9SC0azxMI5EaFcxgdW
uIbb+DO6TLFYNiHxGTHM0ErO4gx7r3jRb2stFyKITtae/0EvGgSwEspdGfhXnrgB
McnL5x0h4DuV0hEP1VjvvvmQ3QkN0u5r42px9ASCKVR25sn8iu6TOhzd5W03D5Or
O3jWStM2eVPVJme8Gi9Dsp/jqIgRBafXzz7ryMIVpL90AFxwDvxfoavD19dqIH8q
9HITaki5/yOOYcQTm6RbgQM64lqDuxqvGoNPOs6DBvD6f0/tRM+J4xIB0mE2Vr3Y
NjeiWoxRR0wAgL5Ad/C09UkNAaCTBC5PwdgCm5ST4KJNY1vWfKZI3RurBDpjBnKr
9qP1YAiv3d5VyqsDpo3XQnDtLasW6Hb7VXQBst3hm/DLzwHrlnQive3wrmZ4I18l
Ncc/aK/4e426iI6Xu9kH6UgeIJAulSF3+sN2srwWWSYBnJTq/Kytva5KODnfD4OS
u3Haf2TFys+HcKL8mF/VLUGYArPbh7hbwWMkH462LvGZDgjhJBwJvVT1VptetZVK
Ue5DqsmLyUgT72WiQicy6Cvn3GHFFhpC7vjvI/7JPVCPWoTjJNww3U2ZSrb3gHP0
ZLT1uskBAoIOBlb+B06+uwpby3EfUY6OPMJKyMnq8DM48enJXiIpc9wjN9a7OWNQ
HXhGY5X3zgY2zkQndbRTFGKEd0KE4iZ9KMeJb/wO6G/0UuK24jgqsE0VAojB9xpS
i2kZ9i16J74bfqoPFSInZG8VUxnp7QpcsaS1VDRXJPeEy/UcTjp+yaNv+WpqnFYx
kaHmZ6LRg03xej5EWTv1ZJqLGErYTV+YnBDeDSqt47549I8IPL4ZrjxBzbxnhgCq
TVwOF3R5cbmqAoGUhtrvC4cIYtW5xG7NtwAwAqvkabTw2VppJJu0FKKUL3Zh0oxH
dQhRhDXjOg4Nabg9Yy+eXL40s08c6h2oq/EAPVbBcqZ5p9UjXon0QABrZJi8JYgC
5XHJolfcChmB4gqavjmz5hGEz91x0iGSMEQ2T98GU5+yZK3BxgjMHe7yTyU6CY38
hKlHzoKTPywalr+nBu4D5jVtOymVk9zZTD0DqO6blz/6pHEKgVhLrw+4juOAntsr
MeXHGZ9D58shZKnQU7o99C5BipPKiaa27nu7oEnROn0Swwly/N+kg8zYjlsiVvM1
u9qyNhOJUb1oYbrlnhYmVlc4TubBTSo7BOnv3fTOQJjdfP/Ueob9cwzUDzjaURAi
r6haFED4ntNMVvnsgD+omOL9c7gTEJVmg5kplhyJfSQHFzAL5MGPWODggFIlj/DA
UviCHlpjzHto6eFCgsU9+HJycbgeRqD8axUomfxNYQ0/t4iOWxquN0uquDM00D3p
47RTXlStGFwLDzz+Czzrrx/wWSdpllRxK7VkvzljLgfclo+FY5R3dCEQ6cP+NYIs
r6830zfBj337JHsjfdi36NsV962+7nvCS6iYowW+CgJemleJNr4D4qOa5koQlWJS
JEf53IPmgnccXMW997/JxOXH8fw6cNNlbVhrVMZ5ddJ744+dyLuAIPwH9TBCv3Gi
fR+mLWZuA+dTIDpaEAvbSLMQWbLUT4vgNUASXZx1b7HrRdtM+WTqmIa5ZmL1BZiZ
2JeenJppJd3ZQjzcuIIuKlsDMJCnbo2tVmoLaSDJler7ajRfLtWjyxjQIjcvY8uL
SloGpRLfoUdOdB7sf1gzYFZixv7WpVroRd2qxAPp8kpcdfwxtmNJJcsQCJ0zGv8+
HqSJZXAV+9bSx2TZt+1+f1+E4CxVOMHUz44pXWwnurkhDAbPOyLlbRFmABbV4saK
2yzRs9Zyehj2BHJkUpcEJhYHUc+GQnWmo4tHBQiqzfrBPPBsuUOWhzcmDJfZQkQt
GxKxHCc0cLlBq846B61VggHMvJWPHMtG8St0F7wv9ZQaw4lAkqF8b0nYy8rwh1Ty
HVagFIYqIfnD2QTujaeYU7kAvuR0ox7U1hZsMi3w5fPoHTOscrQMawrsNw9/XOWR
LH7o2Mulbtpfg4IKLRzLzR26EVIzGSJRXQEfwO6t/nl137y/AD+EqVvMjzGX4YSL
by0+9wom5gWoetV84gGqErTEXnBkLh9NAwniWJo2fUFenV8OClqjvV37dCEweLDS
m/BEeUt5Rr/wa2MHGuYdQaUKWdCzkgtP/ekW9EycNH+B5hDs4GieYP3wO+QSHk89
Awgu4lFMHwYozcFaTHCNZFVqE8XJ473FnF2zu8ZEQQYeXVJJm3RCmHs/xjX6Thfl
mMACe+PjtVeR3grE0qDOPl/cTxUfjfXVFVcZSgsoYoN+p5/we68T8FMcU6HuRY4x
1LibqJs2ij6Zz8T0RENMBZijsLMCwkyrS7CoaVp9OVFSTlrzKTS5reh2exu2ZhbW
hRYw+gRat6Fsw9zgLno+sUaR/NT5Lf2OBEnCzQUZcrXbmzI+t+nh4J55zmclkXvr
TQLIv0AmUax8R7eB15fOwlvdE3dUdnvQruAIF/x+XJgzuVa8U7HuBtQfdns5OJv/
4kROTDghan7HwGifbsKW+XyD4/EnQSUZwmGMMNsftdOQQomHtKSXErF7CpbLYTGx
XKeQ9hINAra20zwViEcoDB9aJJSDoJ5DuKxTdTlsDUITjSKzl51X2wP+kvyGGJQg
9+3x1vbAnc8/FEm6UzyqwWNf+ev8noSo/hstCqb74pJORXd2Iwi+T1F5Iw2GWBGw
I+4/KjxDx9XWymocLadWI4W6lkFHapcayFjC9zrCz+adMAtcm895YLKw2f3dSiQq
V0isGQzQBJ26DJoIn3pX4HXct5XpvzW2Q0NgmluuwquEDC+MFeZ2n0GAyI9DUskC
5tU5FjE+LHmGCQErcaKgwiUbdHvh+Pta03lset+mTW0dnoW8whriQaxT+svg0hnh
1Wwkhj7ELJ12Ct5LAfOYxigSIXQmiAA7IVNYSqy9tUpEb61bIBjD5YgSRZ/8RbXh
xi0fqbla5Gnr1iDhQXO/2+Re4ysP6IV6Ym0yc+8RH8Gtuo7hc+q7WcOhYWsNSuWQ
jD1sJsStGVruAwDNTUKL+FScqpjp8ETONUO95O5Y/g3o4AU8GCM/i214tv31FF4q
mHJVzTxXCnNcI4w2DdoJbNguhqJAKxBh17piozDOfawtfuuByvA91gsgUfR518Is
MFMa7drLNkmkn7Tb/NG5B7SPb2cAiBK5vAgDnHbDGpE7EzsS+IIqI0Tu+xrzDaME
DWfTADaW1rAq82UIFZNfjEObWSumRTPYlXeljiYudfXdc22l7oJSQFsPnz/wuk+E
xu9xTJiErh9NwDylLUAtGjH5+00IEqrHqElAXCHCP/ZOsa+E48bPVO2NZ38etPcu
V0Cvmm6YgvQLD1qjuYZQAOYBgjAWQ8bj6ZC18FODPsKN+wr2PUfipM3hwkA1VQr2
SvFKRiMeXbKKyOZo7CS/tfTIyjEIMgMLZ2UYUIKGqX9zthUHMGLalRIE0quG8R89
YzLO0W4gGdYKtuf79qBwnQqY4yuma2FaDUJHB8uR7ZdhVoPNn6TFuuQZ8av6VfvH
ECoBewzKXOMYUlcPNNTsEvHRKTdHABQ1AZLtjiJZnEmfP02WSOtYV/AhjzOhnRyX
LAUJkZpc4Ov8rryV43GaJeDhhH0mESSUwI/9HzSMaXaZVnVooy6+9BuVZU8+TG2F
E12s3MIckC+nFzxWviHBD2UPvU09kVifRuZjWKsQ6Och3zsJwUPtWeokv6U/T0Um
Xo1wQmJxhFEPd25sUdwvhIS67FlYdPpBzOVUDO2hdplZB4NnEII6ElbRHYyMlMmi
dZ+hQvTc7C/6BmOG1tbEM3vi1awF9LLuG9enXHkOiinS0MmzODC0lcaNP5JTH49J
aIS0OcrLNcHBfVA/j1DqGlBldjJM47JAKeSA05wtmEb4Keb0p5lpwaR7Pf9EHRjm
HZV2Cgn6zif4Upz1sK+3wOJ4nP+slHwoo8RgguSTu1n6jTWTqA7/hcUJxNG+50Ec
a4OzA3pgfuMcklFTK5qM54dgcfZhSnUCZjDaAX12/5L6cZPiJWIMnpnrIr58ogb0
VXDpHXhapQ+USEbRpSeoq1I1kV8LrqOfwBsRILg7bOyYXB4tQRoCYWoTXtg62j+M
TsSIm4C98dNoeJ2avER7NKUKG3jptyKfEyyFFje2eQ1OuxiYbYV3PtUPFk0kvTHx
NgHdgtcDOF+Pd13ZS6exPFIP65WDD9yv0368kVJ+pNlGJ2mS04g2daneVAif7X/D
O0Hq0KttLTiVsni01Z+WSx7icvlYEscTBvAGK3nqBwlvvO7Gcs2FbXsaaakkJVP1
Zjq9JHiQizRIsWAq0pjqqEc6nLLekOTxm2z5MHRQnP+WLbU9vKThrpL2Em/x2ltG
GOnUjI22HdwDXGQmJFjznOmG+QQIphOUvcjAjRSmnbWGgBdgw93ogX4wKGjau26m
Jt45Y3q1/UCIMeu+0yvDIPzII/W1p8CrLQuSjcmS/7mLqNJ7AQJ8IMF43xcZR8vV
2TuOFHZfK6JsNfIgKJodICR8Jv0mdb5pb0V3thFpHiPHq+ZqcMzRZ0KJUnGG1OE5
EjdPP/jBsvhLSrrGKp1krIXqxdR10Y4V0UbernqKJpBSuCTNeGae5tt2EehxuzvG
HVLQc3WwifpH9VKTOmq+gmuZVFp/2EOKkhQk5SExhQNXYaZLa1qk60O9NbdMyzBb
sZ8B9AwtC9meSVSsjuSAiExR0qKrhE1DgQnQzVtagGk3F2MPxVO46LKYD9Jljm/K
1og68HAmrZpNN7JTNR/u+VqQjGfY+0HPQF6tQ/XWZJhk7wzo2FM5s2/8eDIEOM9x
XHu6IWi7ECjDAYOg8glAoA10dbYmZ5lk5CrEUinbS2aGK5tEXMylQm4fsefkAiDE
7LIdP0Lvp1I4D4BQiWh+Kpuf8W2RJoTCvVR4dfRXM/A7Q/CKBerAQyocSHBgLCU7
RxDosK5d2Rt2TyRseru8zRufyYUBoRCy7v2r2BSGxh/9DpZDySHGlYITxzBzXEwt
NtJfKulXsCYqErP7e1C9uT5PGhYPnsRswp4Do+ie8KsI32K/b7ZnqX2IfPtjzDSw
GRZoTRD+QjvkyvJib9q2m/jNhOEvxS4VzqblIPMGbO7Jf15zju9UBJQgRpZ64zN+
ou7qzSe3N2ZVLq5KPBsM+pyDv/rSATp6DCePWK4qdew4n/PsEIza6xK/LEuZe2kV
BhZST8xAE2CaamDXqux0/LdXkbcHBSsJWkW+xsH5Up3XQhppCMq0P8cR8Fcpp9fh
aprokCjIpqSvVQBdpJySRwfZ5890wMgEv8dZmHBbbIjmatz7AIwyaNAwUuM2BwoX
BwaQTgojhibtepPIF2HZPJx6I0UQSa5GhqaYN3qqnRy94Qr1sVu63g33JCIc9zXM
J2SXGWJQw55kMWUXLDDhkFP1NSlVg4QqWIraAYGvdqboWK+A07BqNJmDICqhkIov
I6MmC0ANUnm9wybU9T+QsCOLPLLdNu4uF0DDLSfFpTvaD1bDKd3WL3pLNFwOPGzT
i8wbFsBT+JFHXZY7EFs8OoJugzJ6TptLYrmCENF9ZjMTsyv4+/fiNDQ9P2XFdCe/
RxcP3XKnLplqlqCoCWgt3s6KnmzK45QBGfVzTeu45rVRtYZf2tVtQXwkyplrFI9B
KS8hc2mL2z2BRi2ioOBn/05xp/TwtTWW+7DeQnydnehNx9nYWG+IDujLh5bL4mQ9
bAuwlA7UVUsevKML3pN1+MPxlinZS23kYPkwj9gOAVR54geS8JOoNj2fu4nCmvPy
5rDXloYxr7+4bml7Bcfue8Js39uDFkQcM0oZvn+1R6bTHvW9aOc/tFjGINvfXxYr
3Eit48SEqcUdV+AC84QUzF5514dtuG1jjqt6DRoqfkI1IJGi1HHhC/gtRaYSiDAG
NFy7v3E+fBDGcs2RRnKAwbjFb26zCtKAby5EDOLtqkdttj4Ef0VmbCxB5XkNUpME
duhLH2VoYrcwnJXU9/iT8Wdi3JE5MRU6EJrkO2uSf4bTQMTwOfzuyPSwgOmdCoSe
b1Mi3FSPCLDo9jymD/D8HAv/A+riMDInLotudVQIvv/NWGH65MvwdjhFp67v3MaF
Uny1xrs+glZa/39sw6MbGq8QOw655bf9iavi3iJN7XAVBJ2vhOT1fbyABW93Z0xH
VMiPIVIdRYZVqc1DvCHF8tvXiAIiMEUis8YG/Z1GO7NjGPwnDj3fpB5T9bgtAwlB
xWliyQlDNDha+gAIYl38VQssErQeKLnSyH/tsi8Qu6GQoInTT5Gwx/O5pfbyX/zG
1mEwoSGHc4icO9ltEU2bCXu0mJEtoiv9DIGAHhnpOQ5xo4oLZ1PllRkh4/uwAYuI
fYCgT3p2h5J71WcLRa51vfAIqyOtACwCO36DPZZy8l5rKIAu6zKlJoOPDFiyhdx9
XiTBvyM2beJNo27QmHDLwx4/e/NPGOO2ZjgKOCfArfbDv7P1ZogyvptkBa2N9Pu6
mr8YH1X+G+9qrB4CnAmfSFTs+8HYbgAZz68XtCm6sVZJ3lwWNZJSu75N9viJij+K
DzRrTH9f/t1NATZI7bAGIEqexD9KwcRoToyr1++4hg6/VMJfW9pMZXDaM2VdQayp
bSohTQ1VNEqMpSB3i0NJJlu08F6WgKWjNPT/ILGu9Vid5AJ33oXH1M/xfM0iNEfF
HccHv+4SOTRSY1Bx2yO4Pjrrmluv3c869UnjQ+Szdcn2nEECOmhIcHK6shkcmWvT
UXZ7da/qmqfRQU4WZIQDGs41GwuuPUiT44I1iGBd+b8WBygDzZoJPB9XT+i5KBbb
WyMvwpyCBbbgD2GykkcO17hmWTkr2KLRJ/1wPFmowgxuVfoQ/sUCl9HNJ9mof4ku
BpiIHjB9CuNfVV+oZvo3xy9Cqpndj9pkvvCPX8SrVJfomG9ZTWGFAFXrvS5Rusl5
oEkzfwv95vRlRehEJm4yjj+5Sve+TNn2Qibp2kSJVdf20cfDu51BriYeOtcvc/09
OejKmzFZKjaKEgxRqE3ZMCCdqQxbyaBRc+9CCF1U/o3vc0i4qiHWhW3K3yl5RpG7
2ODSG8jtf4+MGQdAgllp+JJfCFtWb3xt5ZS8p3XllHfu05mx8XLbTGrMfIM22g+j
3qxyQZ6ghMmJs2ToF4mE/+TnJ15gPxBXXjDCh9SVucNkAfD7eqc9z2vlgPqcw5pR
+LkWk/rOmt5TXtlwkymmfxHwTGr+EIU4TnRMrMIvUTyQSGoNUm63rr2g6DmQyX26
1BNmATFzUSl301CmJQwMRVA6Re0+auBh9GgUGj7CCI/A2BGnseTsKzjjtmGMz3As
YRkfdcgGIvJFkVxOZB6Z7YyI22LeQRieVF9r0oqRMiWsZqPieclr2QVLQIYwNxE+
+zeNuhm2DPL7ohl0YWRfgqCeLbqxJ8J2PobkgiixhAgLOUDsERe3YDhDNQl9W5if
BNGqLY7/b1R6Guwog+LxcJIeuSIv9mQ92jSQG7LcQruUQSLy+fXFTVCJCrzGz/nF
zkaKjG2fVbE9SL6mXsMVLgW5Nqz6qvtKKcwj7ZYnWIC4p/5844CSJEJthQl0D0dI
fD1c5qAbJv9Lmbeuw71FFKgba4WP4jSlp1d/OOm9VhuwklAK4hgX4K8Hov95Mckr
SbBZutPI6OWhXjR2llTbx6MbKQdWQHm5uARpTFhhjYoji8GNI2P4srCVoNCx+aZU
AMCKIMZBHlczZ1Vn4x1dkAsA21ecswOsz5/jusIj4qctrxQHcBsSOnacctA3AQoc
9LVtPb9idQhHhMAVtvoj74ghLZQFa7P5TLmgsDR6F0ViqgcWK466aIbkVYh06G8W
5seWGBCailSi2ZXSJoIULI31rLwzRddBgOTyR/UYzLf8BfwzR9/eH4LnalYhY7Lh
CC8b5u3JORq65qMdSTqd/Dk9m4OndEwI6kE3juUCFJtncQjQ1ME2UVQ2oJ1SIfFQ
ml2XZqS30j4fnoNfY1vKINSsx4QVbBLDxga0PdLROprJ+7nOrPEpkjo/vuOJT4/c
tO/FuNUH8MFrIljkWeeV0plUvfkXLmRYCNdyBcFCjvZOtAZA4KbFrtyg4fY3/lvy
TfUpA0mkqjNJWO2G949Jyz2hr+hPO8/k9obYxMcmAuqkOGChEOagfelSqYWOvTif
fqHg+lRyYFg7X3MIaJZngX3FbY3ulxGBBJNLT5KAB/BEzfNejqF/UjC8OxnFNOtZ
X07p/DWHxafFmHoq4wIAXbHySgEltXn6pdcxTGJfupiaGaIqgpYo7hyFB/zhy6KJ
mX5/XMBiGjO2i2XhKeaaItE6pre7UuKkoDHtLEDeQVhpD6DSmjl/C9jR9hVNaUeM
5ASrpP/F+2g++PWP9cl2Mhv/4xDGYBEasgMP0MWIj+UXJdZ+SUJ0fMkT/mwLgXOn
JSq7ubJohFt3/5dbOIda/sPCKG3Jv7kRbZ1Ii3VOBMgKMCiWN+8tdB6vCItWItEL
ztueNb9sfReBc2LO04Awjs1HPHpkeQ4GMBcNsgtMzYhC445PzlMNMhGCQNSWIIY2
QRJm2UMx0lWeZTC5TfCO1rXHM7oVtuVKJN0N+fKDsdOvjcpKrg60g6+3dEcozjKU
yRWkl+sxdGPyOQyuaJ6C5H7d9RkExdgLtOYqXB8TzFWbjHozYhqnMJYcprHN/jey
p7Jzz0mK1JqT6XfpAzxXNKnGmko5HXi9dDAeC59k2QCDC7zDJUg2cXXYBhaFgiGE
EG4ysNGIL2DDhG79VIHhkoZCUS8Rf6hCwcLm4G6/WjaHeineQS1fQtxrXNcODNzP
7oWF1iDJfAJSpsuwxAajOhuuB1xhUID3qhxVGbwDEBv85EEuZLrYhx1StSD2BytK
9XAyi67Kx77xXkcBEnl7MjB7G0rAYY70HJy+gzZi/G6ejFH7rPZwy6hvvUU52diI
t8V53i64jibExYiUUdav2UOvlUKWcav0YaiBSpFEUfDZiu7gNSRHG8DMqmn7iI72
l3zgBy3VNtFvYM34h7l8gKK/P0fDW+STpQwIEnME9at8ypRaV/RYG5Yuxi4Ml80J
R0r3+b0JP+M38LZteWcMPgUc+II3uIZdQsKO8vmRpYyIn/oBHn88s4GucFMdQi+Y
BNlbzrn4juGvJ3rsoNLTnhJjsZwbR3yiYyMfmPsdTNweCSdemRfXaAFy8mzopfAQ
NQgk8n1GI4dyIEvKDPlffx38JGAy6bJtezZwcdPryhMf7b3qFcWcIIg3eE7dBk4k
D/OOXBewWtKjBpyjHEYarUu5lVd8JU7T1b5zQ2H2YmBZaiOUZoGd//lhkK8n78WK
meYX9Z/L+t2z3Wuqv3eJOzJK/7Xo9nFfpoJq4NDkfTbeSZW8JoOlezUjqsS7Yqu2
d5b3/yZmpfPT69V0GEK2xpw6+A1wGuNy3e4jiY9g9N4X8iqoRoV6iPkbClHazu6W
U4Ak84Kl2prc3DWi2/K0JptaDOaYZMKwyM1QdSgK1ESlwRIGZlkHXsC6+54kwkRy
6lCJVcp5LfR9Gx8eyhxc3/4QZKQaVOoaHV/S95cZAed/YQFhilzrLcPNasN3SASf
+VBrrWH0b/6hQGCxAM6tsHmx/QN6ne+5sq8pnLiRvWD6A50Gkm2tIyrB6bX+mnjM
/3ZfeGbnmqlUj1+ZAGGaorfIEO2yCkFPmHqU+AwFklxFloSCxs0pxcqtWmDeW4hR
w8yibmIT9JCkmGHheDyh2YmB0gf80Tpx23rjC/KObatIg+nJ6ux0v3yC2zudlfBu
j1zgZv4RfzZEkj6iLcxONnNDJo3QfjjfUmDxxrht7UZG6P84+GnXp9lrRMv3SCKb
uq1pEQBB1yIm3yR2pfYUEl/uA5d7Nryk9j+NTcVZu+tySV+BZexYNEkDx2jH7zv4
GGKDYwm2ZojMYMusKhgHp3xp/phAgH0IGh0zApKlgSWFY4UpeXlBglpHLAZgJhav
x7vc+NXZlptKqPJ5p+U5yyhykfBoFTJlgGvIgFc6YKbx3NnCC7bzJE4LLpQ6/Exk
hgFsbkeoSnSUW9A29w4TMl1Y/cVBDU0yNngRm6MTY1r40uCQU2m7nxmUD/xRTlxN
ZhHFxDJ1KKYUs4Wvp8QhgRrCv4DvOgvQ9ZHX1I9NBmFRSkgyLxQ52WrNoS54glcH
ShdNwWrp0MQDDBxEcA7CChrgggWyt6vvlRq4AUVfYPRbAczauw2Y72jjPjO/EG4w
3qjY9w6aiKRC+jgQkoKR/+XgzzmxtrYDj8DNjuZ8glzhgHqKiZcGJMxM+gX+Ds13
Oe6pH/H3gXk7sUI1PLowUuQs8gszOO0pALjI2VOF4w7ZSTMhssOUhU7pmIWDKJfm
tmhrEkpxLeN6zgqv1wq4dXnnTMs+EckwRH5mlc0rpwnUOHsGRlIqVgNj5Q6c8Uz3
ettA7QJ2sahWPSqx/Wlq/KJGm4crKWzhzsL2ww6k8iGF+n4mAkY0jM3oN2nBoPOW
9vz0z+3k1Ki5tsJoVbzYfDQjIBCSkjO/aCzDhROXfmZ0TiGMVfssMLTGDDe2VusA
vsnNFNcYp6tDbwMxfgJTHvmqWfwjWtlocvfYPo2Y5xz9lB8SRhYpBb96pfZugJAS
WjF6d6MUMRCJ67KKSASwk2qFWRDyYQPCQMM9GnuWeX9+eruAZSjMLNj5v8Xh3H0W
l5CUSh0BiE1M9MuLZhNHOXPHHbZ2VlJrW7tY+jqCtzE1i/IiHJISvNBdYV1w0E/J
HZ4+M661GXXjisbIRnpf/9pm6DLqtkQ5w50/XqBQfe/QmytAS5aK96bejveeCvl7
EBjgcDsjX5XIZ8ZgOW1MeWgZC449ZgxZ19OBQN/GVWvBpT+1KOChBz4ZRa2jcm3X
qoO2TZ8NxG03jAjHEK2YMXOqaZ93svW1lIBSvho4BqP3LmeMwqQ489jjzTfc39xG
BQf71TBrx6nrNswnLvE5bX7h3q6ZDBR48sx4Y3mPn5lUVpxHHMPktx/AuPUiBwc9
p6NkGb7SO8udg5aCWqAwzApJLBRKAJh9T0b16DKQzJ1OiYCJDIGPzhxmzXY3BExo
EiPDuc01No/QNwT3s4jO+MF70vfvFocaTFXYzw0epAP38p7BAP1pX8IVG0SNm2Ss
5p3NHkaLF979hm1zvrljjF7TvQ8bUWeCGYvpvw9KUEty1AnBVRMubffqDJgRXPQ3
WJ/hEq7cokEFcMuchERE3WXxFWzZaPyitlHiFiSutwuBkzfPvhSWbX8X3+4V0dhj
aY4gh/7VNnGXMnpPdsy0P0qwMea791KGHVOxbkNpbmIYXE9xK9RAFmuzQMzgAWGQ
z2eyCcfJ0B6UywdCNzNw1VgKVSgR+0Ykd2z3gPnYHdDR+G3mGfhDmweSQsRGRLja
NEDM7RHBv3rEVTQHkYGG9f3jOQMZs7dqTG3/1gWRd/G+p8lMAjThO8oQnGYAa51j
HgpIf+32NSqgnXaZ8OjgIDkdHk418STyB5226k+XZr9t7JHRJg4vkYbKHptssa+2
oRRR+UfR2aGQuf2DrbXrIVlpjkAhlk0uQiu/UKhtKNxo34bRFnf7jiu5lyFrP6Uf
QvINUECzkynmZGrwRwZW3/RS+VEyqMXrbg1OQ9y3UsxlaKn/M5MVHDxA5drO84b8
GRdE3ymWmEnzcUNkgNEVVjFCjxzjw+4KRxVADnEybKwscbRQUZAsQ5sMCUmkb0ry
FFMhM0TiVJyd9awCkVSDa3BuZJRzJgERpqLyP9XpyfY2vTGQJyf6r1SUFQpIL10E
hZzs+PUUXeTU8ZqdfqvKbfIJBrRdnD6nVEDFJm70/JdkTIhO89RMqu/eRv+9ipFz
p7xkzgqDdUDcP7gyIY05tBYG+RfCsQ9wRIg6lYnFYNIFk0RHcmioFoRL1QENAEbt
cP4JfCxRRgtZwiJFH2tZqSx2vAV1R1IWckeTKRRWVS4jxCKSQl7Bu9XfZy2nuGHy
fXeUwSknDIk+bag6RzEI6Kcdrp0JiRw3FEY4SsVzl5dWg3cZ0PkuUpU5G78+gfzM
NXAxDTidjtSTv4loD5i7nnCgEFO7pn43yUXvk+ipP+aqUO8eQO+p9SDT4Hrb1am6
uRO460nUl5Stn3/uH9XXbVAscEHo/NzGZ5s2aNCfyh/D8+cOnka6ZdOHBBiOaVvA
uSgRfnd0AJshyGlp174JNgD69dJivewudKr40FnteDevsgZD5awKs1qlg4sXLVFs
ep2Jd1/U0VFGh0B47kkggXNbGtbEQU23aKdY1I2t6Wi/mOaaOxX5fgLU2ea3rk22
XOEyGZocKWa/uK02N3LHnVgCbTg15XdfqUlr989V5y9eId+H5QeSxB0MauLYrjMx
b08V01wD/MQK0Q9Bo+OHqM6TpwJmrIbYo29Q4IS6c7+p4+xYlnj53oqrNdOOqouH
AJor7V5FyXFKbgm6cwPs4XmyCNeC2b9MzAReiKBGRjdzTdo5P4DpAnlSS20t9bPP
pAz3aBTCUCuMXS2CmYYhS8sgdPWxqUhydE9wA/Zuh5LnlGp6PYhD5asHgmyMRAtG
4R1UhZK3ph1HhUT8dUx7eemd1guuHDk0KflOHlBr1qH7GJqKcxmuz4t8ybBM0zuL
rT5T6K78+zBzVDQ9TfIEM8daXIYlPai8HJa4vIzEOEijQHCZhq/2WjjPJneaJVXb
bYeUK/WQz4BC+006fBjjEsbk5gmoryrWmi+n2ynlQdXKLPewHgOwqdbkTbjnylog
9hVr03JLUBL1CfRJ5GWrNDnhyOHUWIXMaOrPDK8RQTYtMnlHXxjxdwLl331abSbV
lTD/M2wJposmm8IyNNhmwVN26TtMrT5VPs1sR2bu6UyR3NhPKOLwdeMiKOR683mo
O15UocxiH7vnRBzcOPQNL+NiYeVFEICT5lEJqP5c/CfS7Ell3e5zXCaorADereQm
/RxHmbufBwL+JIbMkglsRHIEvJp6XeohIlH7+1uF1OfLWdK7lsDtrLgaRyq+K00u
u7DzyEF1Cxqt/ltaKXVlD9XPvp/WnepZeGxkUfBxPvlKDoDeqh6WzWEJrmGAI5R8
fvwfaeMx9MoGsBbo+i5ZmAJ07op4NV301jy0t8No60V11w0B83xxHv9byHKvYJa+
Rm7OB81M1by83VvgKlaYjvV2MwK0AQtJSWIU0NG1agz54XZwlw3DC0MPViPWq3WR
CaNB+2mrkp8eoAnJGfSla/t0Jrjcww9gpYZYUlwbKbjdtdW230axlH7cv13EOvM6
PfE/e31L137m5vWHnjQvoZqcJ5mvvuTZkKhzbIiuURkPbeQVISa/ZmEzVlrmq1cD
hSVoIj2kGYsh9DeY/Z0318tMllqH7um5QuZqDxifGNczi6adUsvwRzRuxXQvoE2D
RQavKuaF/wXijUK9YO9ls+OENr8QjcAufFbUCLGxYrqxDJOr4QVa/hvwgCQwmcRh
wJIZQtLiJ8Of0kEeDrlawG+PsAAcp2o2Yiqije3JVB96lymKZ+QOXUio75QOQ8CY
lWYE6HJUah7ov154yImymNO0oWiwVg6BFIGHCgWinkIeCYxEYnjEEn5xs9fw3Nf3
qpQJ7w3Yk2X8KfOtFjOteKq7wy23HHLFbB525ytyrC932+/GzUrtVo4reo+QU/2y
TomEEDfOLCAvTr+YDCb0RWU0YAY+b9O/N9f1nsBBuQsPLIjEQrU9cxIjMWRUu0rn
QNhDX6lWxVDI3OZHBLNL3XR1YHPnnNEJdXEMzDifb59Ujjda3GIwxsANfzuGyjfp
isKOuPnYy2eXHrJzwpyFLM3I5WN0i1V+XYvE4+Vnsn57nyksDOOkmaECSkjULoHP
4xSyx2CGwxJJZv9IiTO1J9/S97tMJSJ3e8pEGkIw/aXBoBroOu3zNwz9h8Xmii1S
TrMZG32Sh412HgG4PWjm/zoOErwjkXKBW0JkUvuJWWKUpbUYYtdxpirXctmGwtYf
pXejP313HeMOyX6qEgKA7Rca42p7UdY11UrEeJdyF4PEOk8jhwnJ+uFjcYNrKswR
aF5X2vRhiOE/8K1yl2Fa1heSHz1C8QOn5w26pS6bYTxtH88Hhpznm2lRaOjKVq/h
gyqS8osRg8utndKxJBk3jYuD+565DJWT8JmUda9mZN0wjtLMIM/SZ+AewsmqgIa0
3EHfkiIs6qaBVmr3bdMxFaosoDx4zWTSTR7KBKW1gLwm/kRmkDwv1035hoy5Bai2
/F7TiSZUTPeqIdnx6FIHsLJ1gcrhxoJR43ksTcDW9N7GZhzWGfFTgOtX8vAy5M0L
Wn087agGlDxbj2I8tpXBIAuVM/shu+usIf5FSUUjaIBOgX7S1GI3JHsmBKZd6H3e
IK+tlBkOA8Sae0Zk2lkXgjesCZbSx+VqVUSgq5q1t9LpE4ipaEMeKOggJDmJqnLB
sIVqALbfY4RrT6lNXy+mErvENbBuXmQ928pVyxM1onzh1EvnKz0FjKqTGzg/ug9u
efH+mvCL68bA9mpIwHjxAQHc2jDpnGTUJUmUu1whpmw3T0MSRrUUMbIADtxA3qRQ
WnTMgoGPFSUrIgyFn4ElKeao+6kt+cppcRMwzaJnR0l3XVdBkL7VjJVYmhdjVNef
uFzD55JvVe9H0aSu56wUBohhyvt2YC8ED6i+z1t4oZz6Tec9kaK4aF/nSssg4+BG
smTzGme0zA/h6tUF/vhIHWQiZmyFzTYY/SB1zHDHYnat6WA2etJXYe89eXvf4Y/A
08YzB3O9T6Pk4JH96O7Bs/wWS5c1Qr3+6sJZX7zqD1TeXteUomtusS0sve6QlfSg
dYRbvvBptNaOP3nirKNTbw6QKo3saOCLkkPJWkVE5yRIEFJOG4836n93qYKLFh2B
9YSqCUsP3NgxhclsEroe5pbNsl91ZZYKcdjhHl7qJsa/+kBZO+NKyVEcCDOdrkQr
Y9lXOISsTa0gl/77zrN17G6+CYty0eliABWReBkGBtiXgWgMzNMvrj2hI0J+j9n5
ujedQrZlDZQKpbt9XUYkIn7OyDqJD/UYM0XPKRjdXhz7F4phuHm224YJyHIGKTfm
81pnbGYvqeXxpx2jQA74Xw9DnCAqPYoqkEKBKZku8+haDyRonGW14EdPoRpKL7di
ikioL8mJDdRVc0WWad4pdL8cE70SAPip/n3gxH/jUspA/F4HAbq+ezJ6Hcjm5I07
OdPCNzS5RLA8xi3IgjdVi4t+VzZxlMNHrlcHQT4UpofVj/xiCMSDzSYYuEky1NvZ
nxluuJF5tpFB2QXRCD3Nym4HDT3eJO1Lyhsj9vKgkQ1dXiLasWGcHq2d/ThY4ThS
PJQT1xROtSmULfb0pLsizhr1kvL700cQ2fVbh4zaeCQZBclZM/pcZtxjm0cGgSkB
SjXcSZ1pXDKlg3L4wGkBr1GQ7LF8RvR1aSWPFxTVfFZmz7CY8zK1cKG44ZJ4AER+
Y9RBaWPDsI+33avYBEYF1zRLM7J/u6AtyI/L69RSaMyjL6vzj0NJhKdPrNIY19rO
xrtiQdmlNG7b2p9BBAB8vkkfCkC1x1YyLtHvolmbmLpnLPdMzutg/iSRs150EnZm
hDCpVx9bKrTUadgHKoFgq/JNKLHix0FPGKe7lweE+2ca1z+MxJSLQT2L5CQjFljT
iP+Lo6V6uhUPA6KZxhpIk6nbbgpToSvnfWzQ1Yr+Lo65YI2njwB0zNhDbTih5Fvp
s2bgt0Z5v9yjJzPDQbpwPrYdqcumROjAnhOF+pmygaWghDnNp+dK6xvWIhwVR1FR
uo2rW+ZnpBmfMH4juBbj+SPQWFMiTo0fvP9goxKnRvFqOopa2fWpikDV6XGf1bRI
jidGVZgarvlTNXb1RNNacXB/N4QCSQrtU/ktXI45h0KOuwn5Li/WJlJMlMxNhktr
6+XL7r2J/XkJ2TrC2Xvcb5JdLeeXd0NW32lNZHRtzcFpMV50hA9gT8HYyOqdfyWk
HESqfN2yw8+/ZOwfVLTWAbVTLtgE3ktgf7CUi+m7sIzjsuOucMNuyYgLzRMro10o
aRamYEEEiAP877Gwh+wC0o31TxLAQgcPQGrhuZqN7P/bPJmH+n2GPsTdwTydjmgD
rBkl6xbTjIozeLNJ829AZY9sqDwxisPg//A954M+hTXmc+/6uSrbcB/tD+0xBAPM
tVowtBIHM0jD7+Lb5IaEDkv4Kfagvk1jvYEyvrEDpxwz6X+jYJfaeF+yZRQ/MLnY
WWTJ39RYOf2556tmClRBkrpjoV/UysXg3BZMk4meTc7Albiw4/AmCtXKwTW7ntCZ
g8k8DgRD9zc6B4CBZ6ohSlv01AoFGbVxKFf77d+5bg+9GrSbmc+m5xeFHDrgOGsh
4vPlu9dzDu9wlGRcJJXSh09HQfWo6n5uCKV3b83nkAKudWnBbhDdzWVpAVQn4gZw
Zfld4zRB6xKu5o4WSc4U1cS/s86/6HsjfiSAdY/DwWeNrGFsPn5tGuMzKCpQA0t3
O1k6OzEhYdLjY+pzn9YPUrdkF/LTVBoWL0NNRRyAvli5kUyav5VUshwev/GfG+z/
0Bjiu/G63TpQ6nY4Ou5PodLxv9VHYk6FvpuDcML5kuh9ZPAm8f5Fj4taDwe79kMm
GZ9XIL0KagYcKJg7ry1HMXe/sodARGafXVjih6nKkPrCvh0CazN5Rg+duCo76Av8
ujjcpi2yCP7e7ujIEY65IflDMCb8S0QGExypg098QvGJ6S2/wwnsLNos/Wl2Ct10
H1SxNRNVE7L3XXUN8VRO8PzNoblsGHrHT/L6f9wYAqepe3FjnS+yPaW7Y2q0VaNs
2DgwgpVNg/D4ThPh0Roy+NluRbPqfUzPqpRwnJdqw/wnzlYrQ0GoYwvSaonU6Roo
V4LxrOx2TBp5RUgjqGlh1Z7WuIsI74MCu3kSRi867n9pKJwG5PB7jQjt8bBdNDkP
dcYVkQ1boL/JIciVx+UyD/FcryJg20/o1RUupJQRO2+Q5jqthl9vL5Xnf9nv62iq
rPpwRJevoajZKOVMLigcodVl1iUeyKES2K+XkGltQaO7IaeYRKktjowa6aBJvKGh
dmYB3Dq0eQruQvlvbCrmeaCJOUhdHoapR08ElqhvpiViTlwmyGYFJvTJ0IU0UBIB
E5cMe4g3mWCHAHqg7YX4+m6eeQzy6FDAkzP+hWm0Rar2ALUx3gCu9JjhNzaQr+9S
9fLSXi6zk8NZzxqxr3h9WfuAQAxwKqewH1piA48oBwluxx1pmaGljOCRunfFOlM+
v8aFgHHjLTHHORaAAElkDg/XTq9HAaJ4ajubMcnuavhiNEjBDdEEbHPj5Yq1bjND
C6m2Y+n2SqY2gyKcuXJFTPFI4uhtKrKl0vyWnzANzNGr/oEvVaPZtdDis/x1tiVt
OJAamLoCCVjy5vjKI+nOWm3IvrwxIYXRZeiB4A9S/zFLzPO2TUAwqVkY290c/7H7
Cqdp1te53dX8wQHXt1HtZLqIKe4MPVF3tldMUXHtk8b3erS02lrb0JjeKANY56Kr
pMWbM/Bjh7pVj+eE3UWFmh2T7V51b+Qa53dnPZks/UXOgizIm/LVcr2i8eGD8LcM
qOwX1quuWB82akJ7P3PoRdm7CUK2OWoDFYl6jPNFI1w6WRDvsTafwN6/bdYPMKFK
6mDB28wdBf+vx4TDcijBgFjbjyIwl8E4Ib0SFEIhlm3OPljYptgCT4TEUC8TGwha
c6QBTNS/771QIj7sNSozxovALivi/Rz5U5x/jghgisP6HU4u+qvkJC/bXdTOTGZV
yvHe7zWj5QmYTytx3N/XoEunCfcweGmrJI8KEK9CHkCo5TGyqmX1ZAfL7DxPkp/h
zsEfLHkEkvI8UDoytggNUq0AeVYfTtwHevrCp6qZnYiVQe0J9EaqfQvaqZEbzTy9
KslIM4J/OSmR1fizW6y718+djZzvRosz/js+hnIt7mJhjqVu/xzra9sJxcmZxJS/
jxWrXFjLz5iSbNeT+XWpGRl10Q6fLADMUFqO44xDCTsvXogGBbJ5KQfw+ooBxlgS
BH0jEhYXLJAQrUcckD9HedhtHA2R00eUz2p8j2QnK3rVjt6Bw+GBb6Zlandvr9Um
b6akHH9dA9ZRDj0cnSJutW4m5pVgtzX3QiEZ0x/mRxhp7xolTZ6D1vlAroMeds4O
rgDR/P2PNwRECyFxAVo/Ni0IGUBWWdFk/6ZPxrGb9b/uUur5KN5m2t+0cutzkoiC
HnoAoG47ZQOGbzrICZnwa9ZqnoTj6mHTKC7wYh1EMexDzLraBYnmHOoqx4GazM4K
b0xh4MXg8h2lXcfRW7soS8KnMAiDHPlaom5s/oE8mRgCF26bw33apRyXm/nPkeQh
327egmYXJtvc61fKYOLGJy5R/5J98BAiJg70EcmqXT2SfOJVdg4goaVAUCrQTJTx
LOKPleBHANhA+3mFslmkvhEHImoPtFroL1zTvgTPxFcAU2uqx+lIlTBgwm2hBQQM
eaEhMbQ4Z+bkj0VRDrWpMe81TKGk/GGR8I6+DCZD2uMZ70+v4Jgm447wkXC5Weio
8wBUF3/MowoCRQlf10luDL3HC68AobxzvcXTVN2gR9k7sWpK4WZHO5sIpjg+5lK5
UNWdma2BmNU12SO1GhEbO+vevD916HfB/kYmbqfDLH44JnRBk4FaG38vMBBktm50
OP6LDqH6iVFi7w7GeFhXfAT91maQsLjZz6JuwgmHcYVTOefc4BXS9HB3cRZglmx/
w1+270I6wtx9yfm39DZN3vCLab41GsYhO0sxwm7SHFneSgjyb3O/0ymfUl0Tg4L2
T7kAWbe68uILeUvMLdmgNitjzH2hYB6MkIgZRVVyCLFhtDR1X2ILFKI36Kbhrp3N
gsE9FRqkhQg05SFkq14Q8Gnisv3/+uNhFirChQ56tN8C4B6GB24rksGpNATbMiKp
wxjhfrT9Ae/g4WbErdDJH162ltmvTbt3b+42se9d22FJ+u4G8NcCFm8FDdkX77GV
0oRypSVTPUwezlJgYs/aj0/IeGsN2lW2GXTWevKGMujsOnnJKNjFjfcdsLus6glq
suA++Yh3R9fjnXOiUW/WRmGnOLxPXLi9aBpdSAagSRgyRcgbKQbi+ZoDhfALMhV6
6MSvgXuXWoah3KbIQw+TNhpxBVAKZa28R3h4n9BXqxYeAWpmnEeSun72v52qU+l6
hrxSWsGSb3fCjK9H5I48KifSikgOQ9JUYKQfWOwRwHoA4YT/UuBuQXe8RU6azbEo
8+ZMhvqJkSkNgY8dCUxsgWhpCLes05RGuEk1FlzGFsGbgzIQpZW1Dd3CCpB8Deav
JdaP6zQaBKl96uH+EQkfenW+GrWQV/EFyx8t0p2oGI+mxaKqgdOxCXxbxYhS+SZ4
m1hdpiOGiSspGa9DWVxEJc3tJA7qgBGGmHhwQjDpEd28jEX1WCX0w8QyySMP0llh
EHea6ZxDQ1mRS6EZGx9+WmsoK1v/1H/7cEsQZKGDVjuRdsWE6KmpWMX5A6L/+tMl
yXm7mVjtlj6lj9dTu9t1iXdubt4RcPmne2LdbiIKUPqadiV84g55NPfBFFYYlWce
R8TIeRoFVXIqVu5ZV2ZPn1damY2kIMYPWGDtD7HcpdZPtQqGPBddqIScrzksn67s
mE4uP3rNQnGqWPxMK6R4fBcrSWc0ePI9Hdqmq5D5NYHkBI0SQ0INUaV7q+/K2dnf
PrHele3d+U+6ZmuVbW8ugXdNzo43dMVddznw1ZP4IQVxQ0FSK/geJmsWA9hDGueG
VPFqfzbq1EqBmQ9pFPJjz1eDDG+TCjg1+VGL0561XpkWZ/iWcThU/4mbMnIvXO5Q
e5Xau1VjLrSUcsNvTMBE31lcsOf2mj5gkiA7+f/VkT8WvZsHoSciqajRhH7dUf0p
oGoO+/NAGjFHdDeGtS3oqcJRQiwLihkOr1YNEIAVxcvvwpBJVFbQkBFTF1zhclKF
ZCDTHUWkWdE8BV6IVwGk8UTr177RQuFfHHjTz0nY31UCPgBrmSZpUPo7D5RKGE65
8EMPR3GRdIRMcx0VB9zi5sG+lzA8AuzlPf84+KyE9rOXvT1UyafD3buLsN1YTSM+
qB5vjF9KPXDMpWK1Eq9a2GNa5GEtBTiLdprSereHcglFtkz4wMQnXk3r79rOFDsO
L0I7cVEEYbOk2u7K0E831/c+zrTWYnzzguAZpHLkBjTxlpD4UUZo7HS04LBLb5Nb
7QjPAiPT+73+di/KlHIQOGzd5GORG/sO5JBJLgk1iYlB3gmHsjbNQgvIqijD2bZG
W6QUY4Hco8b+t6dEj2Wrb+NlGumo1PBuu6EzFFdBvGufyN0GAN7hvGyJWMh9LcCw
uEn9IZRqwe787X33W+rlGeJCxMdLQmnyAYaiUa0gJb5L65NXagnjaTIktT/n2anX
qYrBtCT4ZlavpnpaEltGlvU2DDJmkP0ZbMheQLq+XdSF8oruUDZqnFUxZDSWJsGv
ds/kd9KStMVaVjZqa/raI+VA/mAwfFDtBpsx3r1/FyscBHfypVhE9mssx+KEJb+W
y4JUmANIViTVK+So65SwZYNLmUxXr+cZUupsKW2GJ6EMx5KLMRaG4gS5wSEcuSeH
XtwlaVsNHk3/4B+vi6jfT5UFE8lfcpfQm1itbVtJYA9H+CYjq/rBMwKAKoN94JL/
THCcPOXXcGPI33fM/hu1XscES5V37y/4DRzDXb5xWz/x1Y232dBbjZAi6O/z/Slt
Gp0t2W/27VTIVLULVLP2inEIt/Zihc/ZAG8GWWhU1QvNxUS2/sksBSNV+SQ8PO37
dER/w6FpfyFNXlINhWjoMDytUyDsLrISg0CaGFk/zd+q4DPdHh7spsUYc09sa+cC
sCLGJ9sMyRNagYp4hn5GAOE2C0q27SjsXrEqdA7MLqIh2RwDlA8di3DJ7Vr8igv5
nAkiPNHXhYxNhJHj0p8GhgKrEEo+Qvwu3piqIPbbpSk29r2kCSWEIxzSgAO5oJA1
HqPAPLKtbfUCRdYJDbhNwYzfo/mg4goLPr4/rVgzk795NChjA+4gBgb+veATyW5/
UYJJhMzeizSpQUlF6LZYLvpxtb8Y481cD5iP49drCbN6+Y7tAOfugcqGbJF5pd4B
I7YyJ7JuhFCL08LvKkt2UkEthxy5Lv6ghOO8vHEdzp3IMYKItp1Z6Mb1X3+SvuFF
QYBq2pw0NfynFqrw+ok/cU/KCYWd/RjKzw8oOGIPYtx+M38hnigvBBUW6AFpznZ9
rHmkdZHKQmg2K4f18BxC7q4Z7ntWqwyMaCze+VHSMooFMSQ8xlajf34LhkAMX3M0
q6RXwHQ5BizxJpbu46BCp/lBpuoSIugO+azCrM9tItpMH7AUIkeEQase29ZO6BKA
VChzx1IkzSSb54ALQF6GuU0CtZztEzbquHVHNyfjm3qzEuNJEqeDxa7kXqGOACui
zQFRrKqOwW5GfCU3xtugKtlP+BU+4GVYe/vr3uDA2dd9jeC9sWOqK5pWQxUsOEH/
e1GTfOvcTNlY2ZgoLCfuRBberksZKZPcifReRjzJSWyQyZChj6cLK8xaGaRK4+mJ
JfED2kNydsC9maUz6IuGt6GsJoXhArFTDC4t4i8roajlYgqhdTzG0Gquw67MZwUq
XRUfv+ZV+dmPNBL3Q3IAy1kkLppyaO6ZnVLo/YPNEzncNmhTvSonuS1VlZRk93tf
4pEjYPPJWIbWLJq1PTwnzfylwCByhEBYbVdKZ4t4yvq7DLJnKJybCuXLYTCGTRdn
jogNkapk9duz2jSrQVE1puWdBxSXtBT58Ob7nUFzxsa7w7pA8nnQU1uKrRMSq5tR
BCtbArHEncASaTG0cBL9mDfIIIMeD9j8kiP+k2MXooZvkktftshkCeFpd0nIcwjZ
ZsxKeOgKFCyQONSBvznRO1VoiXYxdEPzkCH2XLTRuFHewJW2odmjBki9dohvx6FE
BPb1DKUdjCP9l+RsOg8CNtMtbCkpqF5/8VarLkjH53akFByjmLQOZhLcUTEuUYbX
+1ctPS6mxnDsV3087hp3xiAoaAk90zNYIp78cMIa4gUfLRikL18/4GMnxsLHO1hu
xxDBvkZuVTJ+N+v5aSOIH7B6R4W/uRyZ2UQ+UGKjNLU6QjQokuDz4W91gKyOoVMV
sG+mhDLMUHYL+Cbzu8c/fpSVqYgxljOP6pAIxdrYoqLgzSHt1oz10oSaR1IkS3oI
tuT/80zC0rAZyNszd7EVuR8KYruKFWc2WHw8uD95O1Y8BM35Pcsc2nfUdMY+tmLv
Ff131i3tbhdoAwaNU3yB+a6qbcVmrVzAfPa6dQ4TmpFzGhGSJ8C4AOgBhq8AtUye
JZMTRCMzRrzlgytxYObQyryu1E0LUmtI0uWVni9lttGlKd5B8CJa9ycBF6vUgPwH
GQYnqN+yMHWpEuGn08Qi5I2OmP1Zd2M4hJt9nsDZMeF4kTTgZa63SaMkL/jmNRx7
Z0f2fkyTlfwptaOq6lvGi90ql7JcnCsPKiq7xk5HsZGeqX4bvTtXL12jKpTdhJ0A
fuqa2Dit45peSHyuibrG737EifoBC2yFawstMBYDBmQe6/qqJHVTVrwtl+a7+889
S0SIO7O4uthkffiVoeo8VcOWL4yegxC2tupjTFu2MdSEih0ADLPg1ItEs66rDDze
EK+VLp6FRsRGTkkbEyiGuFXfcwqavB5ap3dd8jnkW8iD6G6fPPyB2xvW8/4G1hAD
idrHwFf+4XHjogMW8l+BJL9c9RBJqoJyAbk5lASJbp3AaqSqvsnnxy28EsyW4LRR
99883of4k2sQNtvY4TR+8OYSd1hSaF87Efm3Nr1dmjhpCSesjPwd6isTav9+PviK
uY2fJ1Gt0krX7yWB/jYSDvFduLhVdOaNLsSruwdV19UacvC8FHJhAbC3NZ6Xtdu7
Hp1qW/X7JGf/tJPCmOZc2SYC7+EDBEgzj8S++rLFe8QOUUvhxF7Zja+zV8HBij54
1wBunlDwMwSG3JJqdsli0YiphSwSJuYudUv7wwEIdsnvZ9eZevQtmozjb+nsv8K2
L9tzrbBq7tVLl7IRKwcPm9svi5LQyhnm38LS93NInh3Ojy4RtExXpuNx2mI+FHZp
KtLO97wsmcBVN+26s24NfYogFqGGYFZWAtBu3gGxXtSJuUDzLNRY/JE0YpyZNpVY
pq5UwfNNSKxRf282GVcQxqx7n8e4s1wyTT5rtLq1xKJyhjp6PQ27zxA3j/EM880J
MLx+eh3LQeKLQQP00owCZF/8pXmy9AE8cGO26p0Hos+XMQHPwfwCA3MX3fMYIcGG
TLk/3NyrH2pXm44lw/z+ADVImnZZvgU7M/FDCX11/7plPElXimq+3VYSOMCEOG2o
TfkYquVltnOtCZaWVLwnbfjGFRKme99Wx0FYNHJO8NeEAlOivx4BPrNiofAJ1TOZ
SFyPFLcKEyE1XcdWZvayK30Tbrz0gQcKn5Hvbesgce7V2iORqSXsXneoX+rLH3UZ
ifF22OSTPQCuF52gSCktZ/ULT3D0vwIl4niMnrPBgitH/iKQZjF7LeS+bEhpQcTu
Aj1/cyrWT7JqGg2EisWy8DKOJjWEyi/0IE3I7UpI/TTmMT50CBEuBUs8EGUgIC/x
/tiYy9h3jm57tH0tyVUVfSZOo9g6UiIWhRttsWpDDYhdj5nFrO+SaI2zsnVrQRfe
txnOJDfWOZu5HB0mH+U+ZbDhL18TyeUXCMr0ITveueNa73XpXEsSmNLn6fPgA9am
wC0wV4dHXDWzStLO0H4rAX+yOa0yEYpOPj7rO3YgSbRmo+wqS1kzcB+Opi5Yo/8z
FoAE4jKL+KOXyc8u1fWiYL5IuoP0souZW9OqnznCY+Gzu8OdEP1dh/ahmqwYro9T
fEgOAX7s1mNkV3wgwOaZVD1vi+F7dItCOzrShYNCGvHn6QDc2sWnvDfK8obvLXWF
q0bvemZd3O9Rb3EfbIN+zqCMX/BcwDoCLfWTlZKqLsUfntXKV7nl+XcXfE0VorNK
fwG1P5cCH1WF2Z0orrTSDnfnt2kMu13aMNjJGMf0hasQzJHfGmcyr3bI//S2BrIg
HwCxLt+HCfJsWrMYiR+4gnYzaVqMK/1cD93NVUB8rEOVohSGr13kBc40grd/kPQI
D8OIyR4OcyBBVzI0hTTRjSw09ryJtIfqtnP5uRgZLpQ2aMDF+zHJzt5ZzlBgEJYA
gf6jO2kzcD4yXGd133HQN53uwxh70tdb5MmW3DuFBWGbrVWi7EK5P12DB2ehIhY4
gSwejezRfVUmy1eDmWEc2m0ciEmIPjim8vPMAfGfnsfgl6oMG8uPpSv/wb2LTe4S
fr1xZ6O5UCOY1MIZYPjZGu/a67o7uVRF34Jl7/sD41yd+URgCoydjalwaRId+xIu
BB0IIK/cAjmxP/UqpCxlhfGRhq/VDTlnehJevxnh0WB5W24g7j1ZE3/Hkdw30Awd
LvsL8jIwO6P4ihAcKLQ64j7vgx2Cjogif1lMjqvb2BHpgKRXxid0QKKR3Z++Zy3w
NkiyKf3bj4g6bE/vS1+ypSTLR3SBu8NrRHHt8SM8kKkwkIIDzvFLXqXH5QFNyDH5
MOUCk0YSajdwDLjIwgujiftiOnobXh56DY5bQlnmRFZpY+NSkil3lDAzQjw8gCkX
FssLj48DcOq10NYLK6yXCYwUao+tyfkKlmbN77d8DnWCWxpbTmdNQaA5qFxxirYt
jl2m7WHPjIpm3R5ubljaI3D6VBHUG/VNkPA7ZOC6uGTFILzjqW+F2yX9qGXD9V21
E7a7ibVAeFhuIiczTWrlZnqP5qOteHY8OAmXX2ruhVlpx5ueukR/C2hGbVMhkJ8Y
Gd0sBc005TweojwEHMKzyeA8Nua1p8AzYjeQBmYxMvuW4p3YCdhjudOMbsRaC2vb
v2LWe/2lwPnj9pVABCC6USNTgarhwi19x3MnHD0jWt3ZZNvDekOMDrOaekbQUHx8
ncrR+m0Nhw0CdR2tHXfzkltBXcaNU7pbjxaSOQEJcjnvz0+YFd86sHvtyw5wJBOI
HbGdbtybvbVeJeX1epVbj3AwND+lRvz0xTGj9JA/M8nLlCiGZkx2/EYkaMdYwq5M
AEa/4UIb5vGXqxHm2kaY2npYvVnBl3P0ImqrK6cg52APMV1PfyzIvnaQ/O3l/3Ji
ll+Uhm1eoQTu/Be//NgcV5+F2KACG0F7tJFVpXoU/wRxWi5/I/vqD6SiM/v/DgZ5
W+oGBf0PcCy5tuY3I4opS9HM9nAFDA4YFr4E0W0WNXSEUMkMSXdd65MvejSwk204
bnJDO1kMtXw6CdSYPx3hb1OSkvX+/8s4+gyX8K9ae9/3caGMbudxyGNTVwCa45ai
rG0Ki86O/8QBV7VvaEEnMkEy/fNBzD7G6QdSt13Q5rUJXdW4ByZyJkKI4N+gLc3h
oPULpZLr9SKl/x9pUJJ3SOoBGFaPSyr1LSj0KOUOBSE8b2CynHLXH0pm9Kf8vX8V
6/7VbEtmkpcaSLQYGgoi0Hpypu4uqQ1RCSIohgYdRQdEpltOpdG+PCr8/BQ1iZ4B
TADfMILG8tIbVd8Q66ort1bVsL9pU69093GyZy+zBFgsYRpImbEPeA8WGSEHsZ/B
RbY+Aoat52EHAjgXcL8ZBSPgUfUA7FipuahJlDJMqvIWH0Gc/9BJYuNsnrE6wNil
GnXaBjiNjZsUi4HiAZ5A+lVP0JNfdWb+IGj+OSj1awE2TFpnffsh32WN+4Pu90W5
BE4r4MV8Wy2lUg7M06RpaHMittTDl5VgvT02ymi3HqJXzd8Z4Yys+lY1/TYKwO0C
BRpDsbPlbISX7AMZXGqVjh327WING5naZ1DJ1uYqnNRCQ8eYt3JOsdxWyHrYKctU
SOEFe+HcXDvSCBVoL7tDBAqPIcl/kUDfydPrHXiPFnNjVN23QLVZ4iJPMOQYPkJF
mvHvUZ4iHkx9/9t5KinLv//dIgcBYWnALzQRI2/4gO0TN/TebraKcTCpxGJ+waI5
kGSElxRBYPifKAsXjeFMLXwlH6RzcxKcbPzL2Ik3cdqW8QpMqzWprVbw+yRd50/u
1fNNWIL/ObrgOetek/aMykK6KQYzNkZ0balg4lYrfLBlBUH1LutCwGvSvT75qqIV
W1UcIvcffWJbkUmd/U4lktpFur3uHMZedEUFhW6evQQPjc/uzcfk3+c8/90mSb6k
EdqNpwiVhAWx2VeY51hUdzysAwqa//6MzE1h4hrdRCRmxVkjMDwo77eL1FNPSYvN
IlzcrN9LlK8Sh4okqz3eAhZ2d3sL3xvoprw2gO8lNmo4cZJpzlNLMxdbalfCJqg6
hkK/3RppMVyhhxPl/oj/qIdoxaSx0AmSOxKpZ6sXCPg0dcotu6ZNwHF6P3GluCCJ
aZX4nqxVLt+k5mE58jH+qPldZH5sostrRIQ9wWEIqU2IvSrolZwNK3cgmoZQhL+K
o4iS8aLpBOGaWX/Z0zrisi2MNwZ4jaZMxnBUWZvTs86lEFd851Xb+fhyFM93Tlvn
tFACpWMV0NFTS3k8EUuY5FcfbEb9Rj4lvXlka8Oj/24+fFc4IUdk2ZJ9EnJ2bl2a
ArabESG5i7bXd18JOXNUGLCBs0nbgiWVd32fMW+94khF6l4rxjeoAP2LB+AG3Exi
hfSzp+WqMRRzlUgXgv2XyaFwO4tw9YAZN4NoJfwjOfHCF51P0eKQ/4eu8bHfyrm0
fUAFgdtAmV7dhNDE7kk6ernnvcdBoJOjDYZeg7R8omoevFrS3tk0lU9nubxKTsyP
vBm/1VC1jAtUHaIVj1CV9AhFMiETZFOxMEyBDVSS+DQQx4VeczBOluPAZCNfYbnj
xUq9JtFsDNfOsuGiDJ5B3isy4CSLff97pZxJPdQE2644AkroeY0SAOX6FGlHJdtO
ZkRfNPX6p4Pirc6l1uRZHxr+leWrWiFZwJXTEax2y/T/RjpCP/qkvYK01psNzKQn
vNUcB/ctdzsJjRJwcp8MLWjLcF/9yMAuLoFiFOXTryRdZigybdL03HzsKwmQFMf8
IFsjQUjm9cqI1wCtcByOBqZbO9zEw4Z7ExvxKCMJ4ElJo6SGxgBrwob9cZsuGwBm
7hr0UX3YQDt0Dkg0KNXpxNq8ezVsUUtNe9DB9IeNqnm9PtpHvD59qU0BVjn/Gw8A
LeTYAikKl1NzPwdhGG21LuJrRus/bTztDPioUYww2D1D5FrPpyb7ZWYgw/nBUyUH
/bhnOjq7FHplPVSAw9GGvVHTsGgiUiFFOTLNYLE1gdNHKeM6tJt5iFpnqZ09/cVg
QmykHuzR+itUQqmbW+K9uj4CLg4S/2u7SwBGiUSOUaHnnyQc2uXRVJzkCLf79MxP
lBwKelGA2fp2bVzoNobU01HWYk1mWUwgHn/NJzU7aR2CAnW4yw1Ar+fkyLIYvWFy
lQuHcNzjV3APIgult1bijePXOD0fnkyuqcFdeBLYasLrDhC2/Uw52ISYrBx8avZ1
wuZj8KV0h9fDdvIAu9GsRV7sUzYvZdexXFQt3QCsyRyJSOOi+4+3xCrH7WjX6ucm
P2Cb9VjjNL81bNIwwn+OMIFstM1fV7s1s/vzneU9F9OJko5QITFJTeEsTnGZTYVm
LGDdjf6RzfhJo0aGHsfNKoVAmnsR1/MuDY3xR8SoUS3Cr2XHuqLMziytPYsDVSLc
CPIYkSkDrRv4fCkGvMPWfdohY2yBXEXU9Rx/VNjdEPTY6lqK8KWS6v1CAFqwqXPQ
Rag78Y3sJ/0EfEiKTgBXhaPka5wH2TebUNCUjLAKWZTcoepFd41TACvrtLBC+MlR
ki9h6aDq+9JNkuk1CLjg0zo/k/8lAxXKOpL1sJ2FaBQN04amUfK3Pxath5Eg3w3v
qdfqik7bftB97c+5qLw9/nl94jry1kBc0rD84gDGTXzir3Y0QJK7xvGxED9vDOZw
wHsYN4Kg9cMRKG+BacrRppkdMKwwMcRIHRgOx0eztjLccfqQF0KhSPJ4XWDyU7hC
LWf1Dxj2yTYT8kkf00VbJKfzrekCi0D77fO5EVVfM8qOKL2+bBzF9wLHCgvq3kfY
AGy0Ncu2GyOt3/XJmUNoQ5GXX/LAZQv1yxoBCefr5/DWAK5fgafIXz16lYiN8lPs
Tjo3Lzl/gI9zCZLnztp7t/9X/DYig0Kqh1gi/qVnAOTUn1mHhBTIb3kxmzK32ML6
uLRxW64V6H3TUXbnakKNGo2wywzvpaQTKAV8xw2JsaO5ZatFFtkZXMNQUT925qRU
I7DNnTI4mWJbbyca2kYPIAbVl0ZTQD7pKoClFUhX1+eL6Gf5Ct6CGXYeUf9Hfymq
ucGeDzOHWWqQ9xfEWkjpAeKpmTn9UChYeeJ/v/R8dzhvalX/3vYSq1EczMpOKv03
MFqflUzibTDQU7hLpBi7z2zsV+qkLaehc9bnVOs1D6AuQAytF0Z0ftRLaSKERj5H
LFLXRTjSoLBSJVpI9/wDfF9dNpkV8yNohEpTXwmVQi0R5Yd8/xtffLtFhp8/3V/x
aMXpmxSS9PnY42gRGG1ZeHusmrgfIX8kjJnaHWUi2DpVo8bAoyY1v3/Ai+bHh8Nk
DuuNwZoV5ynBEv70kfjwNyO1WZGszpVnbqkMzXqW7IgQp3a3NZ0kLKS2f0HcYqoA
HWv3hyi0lLD6ovPsHW4Sk3uuyH1/1WtpcVTIRIetTqSRKhBS7J6u2J/mmkSn7hNu
zQgaiE+mJMl+Rw3XBPU9crjsES2SjqayS1lSbTNnxkyBsZ9IIro8zqzRnzq6wLy/
yK1uO1ZC1QYeDx7bax6gFqdR6+cvPpdOYuxflwBLm87Bb0+SB0nHLu/e/stJNZap
ZV3jM8uh0hIrjop6afroyWoEGX7odFUTUOZZd8m59TtEgSNV1PiBKGs23g1/Pj4B
WdhmgAT0lPHzCLMsbnJBB3Un5pdFw5fSSEDg+tRcXVR32SarOBw0hkLKW5Sf0826
RZ7H1qcqs3CMHiHebm9scpkJajXJZrh36/LGmiOcTEDdV7BjJMl2+lrpIEV72JFF
ruBpPtXwr19yxp2F1hs2+TVDXECBXi1OZ6asI1MkAgcOx4yetlTaWVHdZgKzKQcJ
m51GyBtbx7O1lFLlddphPkHF8fGav5NcMwPiVpoGKUOw7e6JSHqeVNYBoi+a38PO
/W98dCKMarvKes9KXmgxyaFZqkkkqpwH82qsxhhG53TLws1nYR2Y/pGOg5m/JgyB
nfSHeo4phP5od8tRrovePbbt+O0Br6LomHymsbBUaWd7xLGLMr/aszubhKAVyazt
pzpRe4QdbAtlAkKNdyXLKncCkFmSEBNGNKVnpoFO8O4D5tfTTu8p7shoKx77dXQr
pKyIe44f95lC5wIU3civmagZvIbAZGugt5bwLyhGsfA1zurfZtRvU1h09Mp74mn5
CZ3/l1kxFsPsmwgEk1u6k63a3c0Zes+EU++nmP3PI7kTI0qyCad1LC93ZmT/lKhP
VC0BIArruLNJ+TR/r7qO5mBD/F9xImiP8+MEuVAjkKtEG2lnQsqaDbnf7yubtWyp
L8T3rJ7hyKPRbUnQhgEDKFM7T5dzbJBO0A3VrQhEcnGXydeVJCkH6xC8giqWFxmK
mnr5zok9flBNjLqaKfSMaktis8VJHeh/L0eT7C4VvkcwRoklFZOeWso2x5reCaVk
a9Liu4PVTbrXVEqe6UwBafqVCgSJ5/YLHyQEvXftS5dwCZ+wC2BdCGVsqmoT6Uu+
vjpcXDNN2kjLvAXYZSgWwTn4G+S5KOfNaRFKzkNRCsXH/B8qumKkkvf2uaXkgl77
uEZqdyb7b87jbv0jb3uw6KB0XAXXMZKw+FhlDRXO3KSQ/9GfBu5w9dJvuj1Jc2vc
F203CKdRqh9HekczjKWjHxUcMY5wqozvRRLd0InvrRYOrInyq4rA4ERsAIduNIyj
MHOdn1NexgaE1saEx3ydqrSgqax7KRdrxfFxEBouuVH+dDHXdzEtYfyuL9AAF8fC
FzHLnRxB9NK0K/Fkixp681JrIkERsnHz+S6fFYVcKPI31mhzOezxFfZ9d9Y2WjdW
Q6uJErTRanWnJF4RRovJp0wGKacKk7GHF88Qk+xgBh6hgwjwRHeaGi0Tran4C1eK
eZGvDP5r7BBQIyU9aeLGWIibLWS/o5Ai/xn+HEbduJGjtSGLMYWZZNJXzwTAqk29
GrSHXrQfj9zDzfyuiPxsdsnCICA3Xn8HlAMQz8o/oAeus5hO3fHF9k0SMjRIQdv5
FVEsVv99tBfnzxYhjVJT4P9mokGs9swCb80wowen8s9uPIYqYgAuDti9KjNQ86GN
+esroKIBpqI27UbyzIGNhNnuLP0q16SsUxDyDhZNhPNiOMZ5423BOr8FVktOgHEw
dnDX8fjTdYJo480drBj+Z9OPnWcq+PBio2dtuwvUsgxgZFiP8+PDPFU1jkVH37kG
AUOQfwu0oa/g0xMN868dw0mBrrLDnU61kXcDFg7cmdmsE1NLckLRJa0wVcKj+rfF
ZRjCXRVczPXyZa86GenbPcc4Jads90mwWmPcxYQgxjrnOHr6HG5qsVqIqzf6u6Rs
o9ePj5evtGSj5E0Ao7L2ne8d5bNsFAVPK/N70scjELsMA5zaw5WYboMNtg7yTkZO
/OQW86GNs3eKVmunrZbm805X8gIgzOVb21i6eHIZ4d8UcT88EEVM+dJT7GIHDkTa
vwMn9aBXpkWkbDVVczUw5iWA54eBv/nDXyVrzOz/caXACeriL5CZs9ruyu/fkZeo
2FT3aSO1rngiYOrPT9CPrYUU+MEnPb0tj7x2dyb2oshaNniCKHpJFPWjCjuGIbDF
Q8TmYRO6KKzunSq1zo3yL+gZVMRdD0frVM2wrk/ZYdwXeQHWqo8McrkezGbQB4rE
iR7fYsaatth02RFXzDEeixBTEM5Fp+/gwU8+b6MUeCeXKzBKKpZKY87zLPgIERMO
CSkjGIDk3QeaQYZNvyH9hJG8CRWiOmhMG59NwpLv0tlZ1VnIJ0UjtlG/aRv4OczK
opZGOi0QhsFZs2FNaCOMMw9pxS+RkgCt4V4UTP6WJJrpNwBb3O/S6TW+92wnKdFb
+mpEPXcDq+VUDllpDLt3CJ5YQjGvMgJTHjt36Q9veiP8NDsZj2GrvJzENB+qQcSK
5GcbgmixMrj0OGFWu8a/ZzcTzvSnU8k56QnCduuAhDGNKUimeCgZxGWMhrb+YWdK
LKK1q4p78U0ERZbgvUOTm4JWuReIpfmKZRrjC/0qDMB1+9cgbbqfdU/JtOIMmzZJ
V8KcuQ065JDCpQM3eZxUYhpfPF6cNZiKXDy1af5/ihGqjFyVkayWRJAlugDqOxBc
UnoGN1QY2xf9k9Lofdhrfww5yiyrb5dfZRGTftXkftWG4RKx+2FUl+MgAZ5QAsuI
s1is0uUay976EwGCpXfYma6/BidAnlXqXqxT2LUXj5EkfohWBgP/fGqbtJwVwYMP
PuIjyglB3EUTe7TGkMo6JegDtLdQG80Hcu2qY3Y1RFtfyxSR+lhsPY4PQ3kyiYr8
jRnikQTAGSw/CQCkR4azTyZ+igsvYHFi7fwbqcLqqUQYZowgdi2SNVJ9TTrj0GpT
tXqbPEsLRLBYqKx1BlVlJzlk5p2Gq/sjBbqmtDZqDFxadPq6dWEqrIFo9T/FvKrD
3ETbkn5CfXpXea9DvK1eVjBX8EyEkrJNZYVFsJY1r+Uej//IgigdvYWdHoaqaM9p
sjUGZSXcS4jIvu09VsYP3gWVsulfuoJ/7YL2aa23DFHKNhTjkrl2fLDU2W+S9SKF
Psrzq+2l8a4fyEAWtdmwn/xoc6vaquSoRO5hztk2MbTrcKeLhiF0dzwYhp2smsuT
YMzqJXPsc7Pzl34xeiIszrlbuvo/giYdzc5htXNZi4B7P6eTjYu8fAsuLeb8suVb
oXElwTh+xcU294jWy71nxnTnu9ATGs8okyimaM0yM5UWhZPS4U4gfSWKjJCTFQNq
wss9KuPItaPLZS8lvwy8MnN9cgyEtMaU76nUvz99UYwAoP+eTKwOZSLIlWpjeWNa
o9jCqgLRgjBTQP0UrmXua3QthTfoJNh88hIjpqdbtKUoyRk5+pzs1P/criXXwpd3
/+d0pvkkHi62SAGG1izRRn03VeBd4efO4fd9w44q2phD/OnWQ28h5Ck6hYJXebex
eEqgFcLOOncdhc92h5nJzWUSsiElSYgEQz9sDjoi4/+v0DG2O8BvOAI9gWgbMfAw
1Do22NkGwOkjUQJTQpAxfNsGCjoDthxAdVGYj7PSDjwiWCnogcj9BJswZqeCNIVb
FtINyI57cdlEPcmjhsJOXEmEWFXrmIlWT/GS7djsQo/SyvyAssbG9D+a7u42P5El
3AIhs0RBOj+VNpBTR2a+aNniOO9RDsWH54L6SFfKBN7RQqg9B6SBOXJzOxqGsf/u
CSbKoKQeTeWJZAJbqZqeeLmsl7VaZC2szXlyXI8JUJ8LfetSRp5Sp3A9A9PPFlLf
NKufEKkb79aaWo73xWWK54Av51Oa455dUsWbWhBn0G0S7sIumXiDT/m8hVL0gxaE
TvUeXaVrSCMa1Y56g1JnqWIJxzsOxQhTPFK7Sh4ati/6kwMms1EyfWMS/gzNKV+2
4rsd0mt++L49zbVoed1CrkQkRz6F9y3oWtaIG3e9v7omjQLhYwxNXKCAp4j9I0Kc
5v4rWEb8KAt+MkQYjt9WVKRUMoTbVJcyr+dM+tIheLkoSuobD0eefYT3Uibv79b3
72CoIwhnszCqVaJo2KUDiPPCNz/ltIkUHTwgAvVDdsQ0UydSMpb+Cl8u06tfEojG
ApjlJbuKO1djKjYMp/v2YdnimlyWasp+Z90n0+kT3bBGorJo7eZ8ErLl2/xaqHZx
47piBVoZWRupOt8XFjjtI/62wwNWZIJsW5AlpDeXCBCEt9bvtiNS941JxI/Wx8Jt
MEl7aKu+SihMPDvkLkVOTlJ96pLLyjUhdUPysG9wxs1JFpxWESXXfNDU3kSMFz0C
GY8QrRsgRCLLRIOI4/6Ewya4C4WjHSGx1ZL8lvMs4YFR8g6qcea6XY4MCDxX0gUf
tnJ2fveQATh/Yauu04In0QzC/ZIx+vaXD4zqflEPAXqLZHTDQ2i1ZYEqVR83Q1In
6sGjYxy806Gp8kp01JP8GepytlJM13VUqJBKZI3/3qWYQizTHE2OMuTQm0KRZV8V
tZziYKtGUXkXbtNmTlqDdg6uRPH1qHcASQy6cXJ2NFeStVh2fbiHS7HxBACymNnX
/mPV/H+Y2WONmm1uIfdtHpOkM+Vy7J5njEAVh6R1+XTXYfLgJOJNNRu74FEoStMm
2pILSaEOcdfWhI5FcTca0HQOfqqmbyaPATivPoYx+Jjo8jUjnMKoj/ZiyVMQ+azp
63ffpdbmFj0qdVd76cBXTnUs4ybKI/Ew9pcqy9bJXNjkpciSu1nfrDiH7f5USdI+
7rXAv+ptvN0FBx7yGvSC8jQoo9LpIuNiHVSQ5sTQzEtZFxdoOuLHTDEyvbfNBvJ9
b7K0gAO89yLGJIfxu8xhpQ3GqxZwXQUxVm31NWxuCA0rliJweDBeS4tNU1KXGjo/
LflHbKgfWzEb+BkLOC0ZUhd4P+uVo7o+oyS9ffUSxzl9LjtKvZ+j66lR2VLkeBEd
jJilzaYHdAV1mfpxfHYjn9DDLPMlqfDVkABFvHHf5oYlp2bghyx7XYZLQ/qbaLWf
SquqGPFtnx/p+BB969ku6+VjBmmHOB3izymESee/cfBTx6HUU4B2c2HYzSuVsw8q
DTbcS/RkFyKkVdcvGabdV4xIQXdsfQrwaQnv9N0+Y/WSiMNICDCxLuXaqP0dBkBv
vtgBuWusGpUhyaJ8qRqmlzjPoZIyJ/KbTQncy8toDVjtnHlFR1Ru/h57P5DwUVrM
/O/eww5PQNzLAlq9CpF6YjdM0U9+yetVUq+fw/SHZ64S+cyDmYIycXdC/w0D6gF2
iJqeFwJFEoLSdDJ+h0rTmO5PSJ+FxeTjAP27IJkjJRtUrXZQo900kSRqgeW7A76u
v7z9toAIbfq7oIyF531ZB8TPKc6Nk4UPO0T0CMMmvCA2Xdc9yBLRsLRNDbbbzAqD
rgHD78N/sngFxPsLQPDanuvBW1wq0dJzJBTq6eMp3oXSfUeXdFm2GHTsf68wRyiO
eLrbSzZMkLljR6QisyEgdwY4/6IQuGFSbwwYwB8/3akvLKYTJYNlMA8xtLEw8Fwv
YoLxytjPEMB9a+X61qlJh8fwzb1O6JacnLxt+LjU2yowp2FKb0E8NSL8Y0VNlH5L
942wTXf10WesiiTODNWS76XwTUF05lh/OncwEa+KOPJ5quPCv8lPid+t+Ji7BUN7
cJ2RyQO0Eu3ITkOrMwtpc+DuezjW1+BAYxTvRJYxTaufqXOG73R4EmaJG87PZTxy
3mPMmKrJ1Zik4stLkFlxtSXi463YNU70s25OxeMDz8fIQGebC7Jzsn2Qq4Y78R3R
c5kUXN/lX14vpmvuZDSP8MWG7t/4uz1WO+Lc8rlkvjTBKvFJEbJaTfiGKlRU8Iir
nlQQy6WbX1srZIHjbuDSE8OsyozwzxZP0+t8ZMLEOLWoEnAINX0yj4l+1v+J4799
m7ymw6g7VfvpLcYF9PsHos9v5CXyxLNWgsuV/Rr8o559seBiy1zNe1Y9bx6OY9SY
P0+tyb5stMScpuKfsacPhK6mcc8/utD1PwFzrcFTcIz5+n5cAkiWSNAiw7zmKQCj
zncKBDwUa44p06kxQufhYhMO6ewncNlvhABuH+ZSxRSsUBBiieCvAcnuCUWSAk3T
trDFvni0//jkqEWuNzMYj0/d+cwmGH5MAUfAJMc1dtBh3wPDUNzrWn+fdNuh87Jv
gQLYp/Fe7MTqoYJUqNtmjQyntgRoP2YSfd3YK0yH+5NCuVRhgujh+AydFCfFdQfM
caefmTyRsKBrEpIaT4x7YoXgRDSvuIZHIy0TwJQ9KMKcN38Ofg4z8V5lJ4KxV/+J
zHKRpFEMkgfeuxfhRrsAS5KHCqaKfspLTCGFW2zmFqFKVXjnEEN6myU9TyXwQHVG
JUR4ytr6v4vKSL1FPItAbnMVCTjkT1sGoLk8xcbwjVzIltWlNa5xcSa2u6hvzjxv
pKJWUCFZW9Y7O1AO14/unwGFd32Oqr2nHJ56fHS/MwWgJA2i53RaZRpV7wIic9ML
rZlVqhyPDHv38xoqY6E5OmoYhzrCKv0w9nKVPcrrkmPmlukZHdB9eq6szX6hvOh8
DhmdQoxBLj+uD5E5bPm9oGA3DRIqvmwPhnEaaQyyOPZatLn2v2xN5xbGpgNj/I/A
HhGlp7pUVTdJPz9PMxv5gFMZhrtMcFXToAhHKniCaoo+nJEMzgB9n5FXNzMcY9ZS
bynUotejBC9Ai+yUG1DccdxhXzRrVjY9jpe/FNOL97ZQ4/gU99QLGu4RebRCAW0m
S1CB+siv7qMINW0FF3m3t2CvVpVxjXfQfJqRAApJ588T5DobVV1yCjWPXqrsYXAV
W8/2e1SaCF0Dbi32n7ehrti83xCvDu7NmjhGl27IMBCWH2Bo3roJEDTU/m5MQSGf
sRlOO6qC5Ugm2vyCPpC87kSvfOXpaRYUHi+cMcGxe5AeAnP95lbaCyO5nmYaQ8dY
dSVbtz08zdGWmsW+0wUsQIA8dVK1tho7dEWXgqmJXlHBjH0XNtmiFdkw9aLba85w
MmYy50EhsR337kFFxkq598ZhDK5ifmqlbYRrUnsv5dpAAKc5Vgp1NPuFxMpNFxTE
O+v0D1WJ5RPLjb1PvnkePv/qB9RaRZ53FTS35/NrdvrvKBqxdbia0q65N05UxoKU
DyVQ4KbFdZp6RX9knthO97ZQS5+RBpsPvtwEEyzIPRJN1f5GF7zcLmqLNK8qgbSH
i4pk9nlTLZ0MmrRho82uOzoohjwIDX7GcVQoiufZrj+eE8qYt+cZ9WqGHtnC08xx
mCHtUvN/96kl4cUC4jXGWgqhLvR5WZ9lB1pF+ShQRT34TZPOdLjg4rQA2XajdC1Y
0BUnG21NzSHO0a38KIcK7wEzWLhNs+LzJ5wyNWHsrZA7Jh58TbRG0u/dNu9PsxmZ
RlAKBwnaiHzczZwIjEMqYLB63NvAl+fHG42TxzKhFq1Nv7/eutOqo7U2mFyGpSDu
OQUMIjEXztIYE2lIK/jG+KD1VRnsfWrb+MvUlWAFuQSRxpeRUKGjPrb8mIQXUKXt
aTt9TrWq0NnMWw/SWtYVfJBOWGLrPNT40FLSTv3i/7VFRjxCuMj8/7fvVxjvSmtp
aWJrfee0dyIFDZ83dWGhLCe/fF20SuU1TYjg0axLf0y5RMQqXUZajfoedJc/2doL
xRoF+/ZjxP28zZejhSbMI2eKwMWBfL2E1WyTltW7QbghYaFgmRrQupNsQV1sXnoM
y086yH2wq0PjhDbka7IDpoTZPLBV79wGEq8RtYwGLnXAGymfercgm/NGhP8JsekT
zNxDFHcZ84yozgTFvJFvwZsFVczko4XgpVqv9vIT6Uy61hFQHLinmYYO/F1uD0RI
uUOdJPGeUZUQgdCDROWzAfv2GxGx4hdaGZmd4nKRYTPe0fS0YTCtc9/x/325t5Lm
+H3b3g+QCjQViOqjxAEvb5pBdH2t4Chbd9ZnlHsTEKRiDne5Z6ypwruaxnXfV9GW
2uvQ35qrlRE3+nnWOMCdrPvGbFSwg6go5+PZ7iGd00axlV2kvVTDfc0BUMI8nmZj
kmKD34dBw1jsn2fHMlwFerV+Z/PC6MMKeZ9+dwSULw5P+ZweqDNLs5FQGwoaIfnL
o7mbX/MkN7f7gZR+ik4c6CQSiFRvaEMjp63+hNpNdoGk2LukYWOduSJIRbYEoSwH
TPmTZhtXKkTyZpugflDIbtyoFcC+EvTMuHchsVSmHO0m+xe4AVO6I+Wbb89/AHxV
39PDyoBn+lPpv+bjZ5zKmuROirc/2ll9zuCwpnA2nl/PAto4P5HCfFIYlr1HJjoN
Qjq0KtsvtS3IiSSLLPsFx+jY+sW+gdb8xVrGMAwYonPtzYuTnAiZyZwYiyZthN9G
OHwZmwt69fT21bLoIRyhMUbjUCAGscbK5Vl6+33UCcETcTQbEtqyB+eX96tT7OZZ
YsdLbseVMbBvUbpxBHswGMDwU0XUuCLpslnDZajuw+t4P/Ovc5vIQNo4d9bp2Mpm
rVRmg48c8FRcGftKnJ1fMkkj37tcYgxejOQ0qajSfFMyL1FFyeFsDCgvq9OIDxmU
XL8lwwWo9sRgAIwW8ckL5xkpRZBPXbTj/fWenXREbmxuKMvAj1igxfJ0ZAooBXMu
5A3JrCJov4zVDGaR2nXdgm4hNYlpQcaJuarSIR26r+oeYaVjtfqZwzvrYak/jAm3
rCw6k4QQiFJoYZmi52GmCnh3EQioZb2/u/YBz/yIkvwRR1AY15IiXRg3dV9/C9UV
P+DHhMscjCnBoSn4/9FqWQ4IG11E8yFPi6nq7CC6QsGZ+V45zkDPp8TgpXYopd9k
byHmN6Kd8u81IMs2VhRNei0AKWxkt4HJSxS7IWxI07pn9Oq1g3zICuEhm/OJgC/v
2s8guYSDqgBM6hn7RRKRGWhAlb124m1n3NWtWIKydkpr8qORIlkcNPGgqyI0bpUT
VfKPZBQSefDkduMoAkle4XgyNiEZARtxG2xOHAMII7+LSwwBswJ9hP0tK/ySyHbc
SFCJWsLBWC6RNyNspuOYL9IBLXTAoiJMhl7c999hHf0jaaJH2zPuUDNyxwSHX+sn
QK6aZHsZUMF8PfteA7HhaSm9ZsHN8D3ln8yGgftL0TJR+gGnik8f7gzVZABBh96H
+QxH25PY3mSzk8so9w/JpUPm1H6YIrGBuwl3Yui82TGbn0DeqiQh28lrbGKPEalN
+uQfKdrlzpbgzpGv3mZtepJp4WyIsjJvkIx4fbaZxEbhMT3yBK0juJXCJlxs7qJd
dsQYRcxT5RiztIVHN02rDA40gsm6zez0XZ1ZMzn93LI3uYGiqdX61cAjbZRODWSP
R/L+hi9p/telA7PHuTAhSeIdDdwPUAcKCSb/zX+rfcrlY4rWiB4al5sCzaXlsgNK
ZpXuQednvOfxY8n2VDFQbvUo8a9Q/HSFF/B6EJEVX6AyZcnVOFqhK4aocEC3XJUj
WLeS1EVRG0lEypZmyTk9N2UPcboB0YPWOREZkiSIQRniADba4ftoGXdXYj+iRmOG
M/dQokOeGesHzTb71IoDVB/7BtgGOiw/UykQwgxcqf3d/MBOnEQJY1BZff5zV4S6
eXT2nicvBxmSahgu/HuBueL5ZN/EgXvtFpC8mX8iSlnk1mquorYBKALzvXjeZILY
FTtWj97y/CXosbLtBm/H6Y2mYvONKQTOmMD+4ssTZe2ZJ1F4EoufzbrR9AwwyrWi
L5u/sK+RPAVlPzs41XXUl2c0tgRShVkWZad+7PhYt91/1UsdFeuA96rBrWClSq5s
63qdrPkp37SCqRKq5Bf7QDRMSN2hSYDttOiH9OrdkTcdlxQLkDpwsNcBX8bek5Ln
EK3vwSXVBxkIjWNm+ANIDsdvls+JzI+mX6BqXpHDfW0mhZKzOtk0qZD35eMZZHzq
p0+sVr02ZAGGqTFrTg4tAaX1hkB3+V+/T4pWzTPcEpPmYzvlx3NFam+j2dpGWu4X
ROtgJ4IFE99C2/sMSUy4G8mSgPw+xjJjVPIpVdkpXBpiW0DMgMCiVQz4l4812dfM
3rI9x+q7YCZjGMkXGsaNp/55nQxvRuA3zr6rSyg0U/KBa181GrfveTxxHXtQAT2c
B/VARpFlB6nwpsiIPXggEr/O+q8EGV8pEZMrP3pHw/uD5JoqwZzyQfM51yFAPP3z
SyMVl8E6ZD8fb8EhKcIjbcJy45uYmruJZAtcrjEAak4DhVJJUIzt6+XM+Wkkum6t
7U33YzojSviid+FW5zjWT+WpK/k5izRdI1hhpXFFWXp2FGCu2Dctu3bhbBnellrP
upVfmYiNeUs4DqHnWCpHznbPEU0ifSH1KmuDuDt7tqJx1v7eBfcyIjsHoIGtYyCz
NmRWsepkG2/g6zRFVV224mtQRXL0yp9CgYSRieaYjHmqxqpKpPxkHF54zdvPxlUG
UWzmnoyKKBUkrOjGR/mcdRRStmnKyMOvksL0YQ2ldGPdt+hz2jAnpxH8yw9Ic4ph
h8Fhz4E5KGJoKb5sVtMzZMkBd7KZHzwwVhxgmwZMDFKe+NCaoCe6UhZhfLhz7NDr
F8BmQQXkm1V1uaRKWGtHQcSJF8A8rp7U8HnFTXi6G2LKSg/TGC358uajKK517JWS
aeB/cCxNNI51pExZz9yGrQZTmw4CxncY626ZmVpIVyi6QQLe5aD5tvMs2BiEoaII
o2OJ0S1v0o2CSBe++6EpDy+n+fg8yXz/Vlq/V1coU5eIyWNvU/iZb6sCkWmoNZ/N
IsOIBzBIxpinJlt5K7twNZKCTXkZle0lmDCoIq6GTg2OBRB4THWVe+gB4CgCmA1B
VQgN2ordPazxa/JzZxBdjQM9fUipbuA0E7RpwpU/2l+eiVN+L3t9XDjW7tVS+su0
xx84R+g8epL++MzofR6LwTv17Ip2Om5AI4T/nBDBmIt74cW1AVUf5p8dC5zxj0r2
6r+5V/DVZ4xyuU54xyifyGWUIgDN/E4LzF/uwZLLlTh5yxfp1J6YpMa7NyBs//bF
eeva13O0s0NRzfwGci+5eq8IH6s8Qc95EO8Bs3JibSbJ+Siv2cFkBdqVR2IK8Ix3
xV1uKtcBDWKIgNFeTn826jbihD31jSdnScyDvYE3v+w9/UEcj4aoevu6bp2/Lnvi
mw0+NdSaj2GaG6dTdW6mDevk8Qm1Wf0FNUzae+hoJQ6NtVG+Go6C1atfhzlSIKNl
K7t5WO2fgTLlG9ifz0Nsf59B+XFs6+4d44aB78tlM6cfwkEtM60GR6bja3K/BOGS
YY0tkVLucdjJKk/TKnsSkHYzFJRIDsSAgABYUhaL+gWSYfxcuLlhV947t68vJ5Ah
P3QiUXIPA7m6+1++dZjYPwi4vPQJBQ14AXcHAstEuOXCNSGgvYjJAZMn+amRWmFS
XaNTKI3Pe0Hgtooqg5AlpUKEH/gd6UKfmUpMm+CPKEeHpytoP89wNIMaf9io50Yn
FNwCV6H+rLxZO4Y4nAQHrighct10xb0gPLTUDKOrEw7b0ccoZZqB2LWqML3vAJ6Q
lWGok5K60rVqvocPyu2fLOOA0Q84KhslgKL/+0dMqBLjR82HGd8CPh0XsoWFqivV
DcsUXx23fh6toszcZG70j9zKbqPwbNH/tYLdBZYvuNh+toR9vh/UK3mjhv0ORCz8
ka/gX2xHei+HJ0WUeeygE56FP+gTFK9+PzcCtXUWXab5wj03Vh+gB1l0YxEMwopB
ic1K4+5Y2iN/37LDe39SFCDaswOPw1uL2GljmiZevLqZjSGHWOzHqEQl6gYRTDf1
JBPlH9ZVao34PDSPvZlBMK2LehLhjdnWNFoOVZlbuLxECD2azB0MTQTbwjmK6iNO
wNngMLZEp9k0HG5zwVGxfzuKF7VMpj8dGrhl3ILdmQf4kxG1krOzPn36gWBPqAMp
zUf2USKtUJhfB6QcqMRCEcgOK5QE2eXHGvdGQy9sb5FtOokLT/fL4krD2pdEZ07X
pyD57jFAwRYc03PUW5UOsmHRcIcTnROFsgjOoJjcvKGKyCpmnzIhoECC1jXbfcNF
ZstUsM0cK1V4tvb/X1iSrUVEGfI9PLgmjEWwVyAMi+dPNbWVpFLi/0EJKn9ZKiJ2
VtoJnVE+kDRaQF7dP7Wg3b1hqNlWKtn+EGsQugeragxY8EfAn3OF72kK1o5SKLLj
xVbxdn+V6xQ6cpOEHbjwigHCIbiQ4rQg4ffRmFNXdGtUDcwhjZurWhGIG07jbzS4
8qqhMjIbrl7wvB7UvG75Nz2mr+rYbppRM2bjA6iE643+Ydt9j2sCgE8iGl0eKVk5
VYt67bidcSsckgly8Fx1wRBFYOJFo95RXUZ1iIzc1e0T2Jt+yI7ETnKKC1LqxhQ3
rSfMVGPV+xDdnupNxfToSm3uxK/oTM0cVWseEx2meScBjvrH5nXZFVH9yNsMjxSA
wu7nYAzld1UjW9yD+tk/c2YQYnB0XkcF1gfdRvm4ffa98vMtte7QKv1xm4h99J7u
ClPzbsM/G2Y7jXxw+csQo9wjI7D3Kerg/W4wRebs3Fme/uVxzlDTpx77RExJLixM
fdmQlCNvm234RJqUbJFT/RSY5OsCZZAMqfzbrlQITL+2gzMcxIsryx7W5I8yJY0H
APfBrhFWGcJZzhSxufTvvTfp6jHeTbP79MKhW84+/DLRqP+vdezWfYYCATfEn7ki
zWnBEPVf0AtBaIbSKu+5bygkrs8z3uFh9GWEsvCSWAJPkds7dxWKlUYWJ/TToE7r
ruf5e6K+QLkN6oacyE8e4LNx2j8EcAJm6wm8xz1e29rtOOUqqiJDsDlHUbeByKDC
jytCpC2K1pMPDMtE2iB9d9KNJTkrXAkUUyQhOjG/Oo9cLtf6on20SAI4HUdw31dO
RQxJEpnd0jcY/KD43K6TyJYV2OZRPWZt1qo0ZyRuh53RNu/ya1PQ9JyEosuUwHM5
DuqaHlBOjfTx2H/1PDbgYVM7zWCKg9O9h9hr0MhjNq4xEV4QwCGG5JxyDYwwO+6U
66Hqi7p7WSDGuqhn6ScSBByY5Og0nViAxz8x/dpVFfQ9Q1gUkuK7jOj13O7eu0Om
iv+D4GR2bHjhqVG7Hq4OQzqRV2ZnUdC+xtK3EYeX71lNKblBGee9qNXoJZ1VgszS
L8x75AOWOdcbW2+O6JK58pPNnoDireuN8XDLHbFy6nNOkYYEkxlnMUoalcT/6ACS
MJ8FnioirYcBSvBrqcW9iXgEaAfUF9uNCSPeHOnM7y23g/amRfe8/Bj7uqP7gi/I
mygJNSTepRbKWv5j9W1pIqiB1t7l2f2SoEUrZfDHr6+VYVzuMHzXUZhO3HPDIxec
qAT7Dp0VFbncr4dBD7RG0f91R0boxHC6VCJDFPB1ezgBAzCZK4kts0FDY4dfnwAV
slDtKZu3LT056i5b+OCaBL8zFSXENsG7bn1Bqx3sodR+Pv1EGYvtVca5s4vVF2lz
6GDT1iIn54uYlwDG4XorJEtUooUMM4QC5uc7Gsb1CqdjBzUgCtr99c4mrXW5Sqd5
byhmOymJd6BDmgDiuCBRaH8GgYJN/OM85BF3PuEe4L4Yr087G0I6jI6Fq1ln6GWn
rExET0FziHe+XrHgsEnrkrXBywkRh4C+ydZGzNYpRvdQecdufkbi20Uq4XxQD+bL
rNEI2HOcXVeuu0TSaGF7V80+UfeDpRiNnj5KJW9d898GmofCnrA9m8EhQC6aebyX
m78gBoiVXDk86Omb2HsdCx/rQVITWnqkFSAaSM6nahEKn/6LiYU1yYfP5AWYSHPT
Gbs49jNP0tx4lJkw6Em7o1xVcta2dfSrd7OkE27EhOTeex7ptRBQ9mq2vNi0NCL0
tVsnQGpON/xSEuFkibICnTZh8/AYLgwutoVJrRLWeuEYaLX5kMupVzGlvjKO3+sq
jQitFpqRpSqy56tYauMHzsw68eXsCvZvUBadyHNrPXeF2cLQZeA8hVEHh4j4nPZZ
WNtsf9fbeXh9TLdPCYwIgrbJ78lCa/QvI+flE0Cmk+ZqIV6B5BZraGeSD5QS7lf9
IFCICSW2ZuyCErmGE69psSPXkF+eSUbyOtA6DPNixgsP33c5JDHZqAe2gbpNd0wE
wATKv43W6hovsWMZALsZ06cqHCcEx0KaxYOyk6Q2cBQDapzgj13XJbd4dhfMel+v
mbHLctUHIX7+6IBuWJQiDuecV3YsJfGJuHYraV1DrwgNhDhOUqfBI7gbIDuLzemj
Nbqo8xBEzbQsssFPC5c89zXR9KljE6BSfCwnoxk2CQ9vQuAY3U/u8G0w1QUDXN4I
exRPaAnQlkPJEJxWPfbygjefO3TRzMwbyn8eS81LHg8ogFAPjkEvzNIpxJPrA2Vs
/8FZ/7RfR6t0y2fmKD7PZ5lzNDr16RfOHPL8BT6aM3QXaUE9JKf/RXcANQYr0Y01
OfEAslGy2Br50s5canECd/7WoreyPcaLfU7+VeN/Ug+3gVyvNZMlPSELF7ZldiGs
Zy/vLwpVqRQXhIxquHHNWNBtJX7bW9OZ09gdjeM2f68WzlIBnzcm8B7+3OKvX6bQ
8FUj2X0E3mJXQa/PMmL/cQcb5nfLRO5XFMPUyN6Iy1o/i0EUIguEEW4KFHBCbyYE
avsM83U4+36Nq23ySMk3XK58/Jmu0eWmvDFiLS+pf0e3DOje/1zYQHzBHLgfIwx0
03VS/SnsJNUS+letAWgE5PUkS9X8qabsmJCcjnRpnVnuOvsgXNcuD7d45X1oOPoo
18bTSoB9L5lUIrDlWvhgxO3gHLxHfaZsXzkaFZ9WF6ue4g/kLVMaLr/lLCS3k/eB
qH1d6IzoD8tbSMKb9YGU6efhdvGH2M5IS48WNEfeGIYKbMpjlprgz6nR/r5OL5Ew
EOaNe4Gx68bwq+14CPleYfRF+OgXfKlzrwG6ihmauBhrFkBnfd0H+ezraU2gGdx8
LhKTgioa2i9BrPtE73+8km9JgyOhXcZHfvsHqmKwVHCCulkAsSQXiB/PtP54SOfL
AaEZgtvE7ra+VJJUit0m4BUwz7ynQvSxhtsWI/QiWPPUiy5I42Me9G5fxDp0yMLy
Gu7WYhsB2KCP4WygI9AuTZwYOn2zbCx6la3oVNLkRiXc6ROTYE/7szwo0VrRLPtV
ZpV8bxCEHE1++vRQXXM1txVnEQPnH3Xrf5Is1v9TFIXKMG8TRHkC6qgOjTMJKrA5
nXbKy/6JDEM82kYLiND8nwXgWMLqSLVTcdYp46Ts00JdYnVbjUrydtPwHYkYhpro
6ws/F1ZyNFSBSKyXJ6ajSPr9LBg2SbXUAa/Int03x+aJbEToB2fV0+rGATVwLMU1
sz+Cdwsr64rFH111svGjZ2zCF1NPp8NbrK+Z+Mz0uLitK6eD9mYgX7656vbh6xTh
taIWmYBcRlvc654jeAtJyvhnhkHCBDo2eMgozCeWAiiKw+DQ9jeC+7wEmxZkV/hn
LC3Y49VXByCyM2A031BuEcz7SDvImYvN+TsDXvrrqvj2jJzMD72FJUqlQbn25fig
4ai1TALJRNVA+Q2SEnlvLH3p1+4edyDYB05Be9xG2JzFxBTuUdooZTKSHFJozwoR
8KWgnoKZ/AnKsXnD/g9aUyUsFYVS/rU2wa6dnEuv+jw0K3j1fkTi5YQnxfh48V+b
D7ufsT6q0cHWmcrATUkn9fiM1hRepkpiRx280aMtCoUJ+DDpFEvVzRCS/uvGXPOx
mryUp4qA8xaURG48PYDw9e8MJhBi4QP5JQ/ivu8HoOdMDo1xWe4vV4J1SF8I59II
iFEs4qr6cpY0wsxMDcdyFPFtjuFg75gFUPO4PXTb3crwOhP3yLI+sWEAYDL12FVO
GFzrcfFP2v8L0jJt499OsqSWSS72Hoe2MD3msqTPGzNnsxFNdDfFh9GpBjDDK+0g
LueelvlnHXaG8KP8Hnv6BV7mBg3fiZLEyxW/G+AS6WC0Nlw1WaV/M1NiQ0S3FTt+
X1mwbueFRUr+uyldqvpeM2GXNTWrDqpzlfWXKNjfnXoBKtPfmBige7eKjV79Bsoo
INiq+pmO7lz65pNnTo5BHDtvHJEiXuvMoYAxTwOhStuH/ZW64RoS0ABL7HERkolm
IulkK0pUt7HWJ5P6RcrTs3EW/GCdDOzgW1ibWLlWmDuBOcIG07dDNXkAemFttHgb
vFcVaNlUxxZ9pZ2ljzAP25ABIOY4dwFle7u1x5pHrsT3KRt9Mqa5CdRuj6SFT2Ki
jiREN4RHrzs4Gt9stpWiKVx2F8k6DXKZOzzm9/2Vx9gZVmJbeS8Y2gsf07TJSzGU
o0jSJj0zuuTwR4DvzWQi4vsCmG1JzVB9yqtFp7TsHx6JIKSc+LE3Ac2dHlpBv3bi
l7hQIyf3tIIUL09IpqEjIc8to0ROMsWgzImDfptn4zz+1GEIgkdbPsnkVtBafalR
k1+7yurI7KVaI9MK+/7ogypYbBw5kXp/3Q76EnRLa0Eh4bP3HDVqUNFR+qMKP6EH
0Li7/mLoIfzDM7IHXydry/5IcFYtUC/FiEqbup1WQtcv/HUEMBaDjtXt81j27LrB
n6tlH/okN2lMc7/CtIv7YK+fMmeExGjyHEMJ0MuCLAY9qccV2R2Riwrxz2FLjIF5
zJyPKpZslcNoocxn986TwfnN8zddHCGoFqjuIyvhhpJVeC+npc1VA/RL4RgIJHbg
Evdv5MBhfsM+qDEdswoskBVR5woQOIlc81uxvlj37yMTY8aj5DTyncme9y6UoHmR
gJX1R+lr0aAqt+EVEOnwO0wALajoXX9njtu41d7rAdz2yyn8LJ9jRKKWODcVOluk
z17jNyC1MO1jISLZBWjU8fMGSzqXjOmlwVVYrcspmiPIR68G0JU0TJusmgcDweU0
ZkXY/7uYIDMTtMXxYUAkaCJhf5Boz34Z2XI2FwiiuRpkzYRCc5yEdY4UiPbqGoRu
mr2gAJUeFOu3bvOMMn3+cpIX2Brix/Rq998EsWielfTBEWcLjq4Pq9Da8sd6716q
+IRzrTvLRZTB0LruSKpBQhLRjz5plVus4P0cqPGZAqJoxPv9noYzOh+Kxu0ornFv
R0+qCAtwGHZZNFe0mJ1Xqgn5VT4ZRwglyKukVdKefu8h4V2WAn4DrLNpYPN1Q4dz
YSof/VWxOayQzd6GspO+Tmr8oXcnU05z+07KoinRDdG2jeTejvxj3FHKnjjvhMU3
UR2tAlCeYUcF+bN4tAE88w4HlhZWIHkFMEJE2mn5QVwqxW0c5aOPUne+BChCH17r
EGzHX0UfRwloDaWaCSSiVoQzgBDcq4yfbZqanbMMDjmdGcSJEEVSO+9aKvp+buXZ
SgyYr0BnFlJV/+c2Xfi4ZpbfDgbaDQOnJaBmudp8jp0gKK7TxDyEbH/X77cVsrJw
somqVy8zirbmwRwFAyuqHx4Od3r4oIuGk/gkC80Tf64+YM/BlaRpNqjzbXm+3VTU
Xy4tkU52o6POCX6HSkdBW/PGypLm0cnEbifFPqzks+DH/PLO3aB40dlwUTrTnKhZ
5WfYCUTMW89MvD+4THAMubF31xH0pt1pSvzVxJhgjGcf4cagBNcRIyEQ04a137kc
wStTVMvvFkgJ67Cg9uWAmIX7T1UY8a6aM5r/6LAIkIiILzGL2Xpeaq7ofoiww0sI
35w0oNSzjM0b5mwA6AX61rS1Vs+cv4C0g293RY3xaH0oKZ7M9C3vTuSH7aFhzwIy
wskfJ489hp2qTa5yBwv+pZeUsGD09mSFA4zYPVZOPTyL0dQPLJ+lr2BJSUbaAoyx
R2Y/xCVms+TBcD7ZVzRSLvr+QcSAUcdv93wwSClGiiHf46bEqpWVWDdf6hbPolUT
oU3+5hU2mwlt/7FPoynYqtMc0MPtvhuvOQFhEv/Aqii4+NmWIzRYVuSWUSGC3EcN
O3It92ZKFAmjXd7Ysr7Ruwkv+UVFETS4CJBAoLSe1AAqlo074liac2cfH91Sulwd
6n3nxrAnMkvP+m3rF8IAJa7LxWgDUyBF/4227p4NFknNOuJaEQF2PVeksugrfBPL
e6Z0bYkL3oVIkN7GYngJ7veuWI7PygXR7fStwcIEXphFQswZFxarlUbSMtzj+PDU
mxXOhEba0dICdamcvcOlQR1LI15Rtf2v/HdqdvvAhaDQyk6lGa+aG09HxmzzSF9b
Ru4ag2leqPs1GxAlF2UgqYe+fhWjLOuakXCeyQr0eTQ3OFcfZ3X7qlFZeQcrK6WP
eEIHrJP2hyzpJTsNvABd8yBQEnVPYTOmEEufOyBCdAc+qbzGmpj3i1IgJGuwqKAj
SrbDc72HcSFwFZGTNbU6hJfHD2bB9fPwuobiNMlKIfWnDzNHKM92tPG9CztXInlz
aAmgmDZCfumjuN2hRHWA9416wOH63eT0mTuLfcwnLX/jsEJsD8XEEYAldz/UjUpK
T9GB5OybJbjziS1jLIzx6+VW8dgD+5o35BjSkeLdmUmGGe529ID54KOYmswEwyDg
qwr1OJEqvcM+Y+b1iudxGtJI+YxyPfs6JpO8B7fVPvySZVw5ARl2B6JiYUn5kTDI
Jl1ncxR5b3Is6wfnOpUc8WaLodkA/D2gCXGvrRwllDRcfyJF7wHqA1K+WS/KIUvX
eHeSVDP6nq/w0fjfvkzHMw==
`pragma protect end_protected
