// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LWMCBzFBFKR+G34RiRNaPLGp/8PEazhNTROG/tgH9fTcu/j74ly6mY3UNkZggCro
Kfj6BxJgQbnUfj0qatTRhjZepn3rd+mNaisAMmB+il8wf/8ORDZF99DzW5W1xQGM
3V6BYNmvLeSlpbiwyJf3VZQGCgwqKRecfwfeQYpdkXE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16704)
O2kdyYGTNgO2RVG2I2kQn/lhXBY7hHsfd3sOx8A79xHvZ3tzy8XMHtg/3xRg4qKX
U9E47vb6tMD9PzH3lP4CMFg1JLQ5L7s8fdUCGvFwoHueKhio9IDTyo6W0AVfgMf3
AtGztIbKf1XJyGU5NG6QXVbusl9DihpklDc6LieJlt1ELAD/0rKB9eRkK8n9QfuM
g7q7GiObzjfxh/OqCH1XCghxrWbvkZen3po4nghxgflLv/6n2j54htL8sTIjQq+T
PlWfnRYzp2a8yUETpvImBbon0gXkq9zQvrL3qA4PdF9jIA8W6CO39qm0PvbKYv9c
1syS1YjrxDvM0E9IxsT6K+Dx5cMBm53+1Wxz2oQoG+a3pGIwFA0le0oEWmdxWj9P
CvcETXKMh7/cH7xBf13VWRjJVB1FiQL1s/X/OckdhOXhsGJp+G39O534cMTRhOxy
ekB6OxMzywDyowhYOD7xB4Nd8VB7kxlPqt3z/lTqm3TwEv2KXtGmjxVFOIK7eN2K
4h/6SAaFcbrKrF4j5VX4vQ1mykBKnR1KAKPpKbFQftTZHohBTHjUYHZzuBJTFHDz
gYjgSpcseVu32S1PlFmCFGzfWzFj9HYgLphOWP5CI2J9GUDTL+EGq6onsx2u0lm8
plrx2WcOOHkUHJ8edGgKjR1YmmENEfYwLESoecSSgPI/Hi0hMrI6AVXaDcCyPLB4
+/8dYiv/8+FDCZqlrO9KJgsg5JUUO8AOO/TsS8w36YOiIQDwCP9QYViR/uf+hEDt
8DX0Mg46azFr6RAk2UAX/nlqQzDTzMWqquNYKBULyDV+5zBIv/fBghOel90fEVw7
QkV2d80r67SaRZooXjRoo5/4iCQXJUZO3XWifkMvPgGSY1BmtxUZi/r/S7j7Filq
MPij5urYThEQL7OQykCmZcoEY6BTADrgiMB/u80Ivj86Gna0ofFa+V/rqiefXlO7
jEK8jFCr+4H2lg66KCWHCXPPi9WBq7BoWaY/PeXXTL5M5fiqUDZlw+Fyx4MPLbnS
CXs4TDQkGECQrD917TsOX4H//oUKVTsek6wRf7Q9umyZ98f/dzF2O9rb7cYrADJq
PYbLDcJMRzlVVKsWNja7IMhw6+8JBp6tp2kSRVvat6MExgshAFtB/u9tuchydL5k
PveAzWnzVvqRqBBxcOSws8ppT4Y/3/WM2Mjxu4UZQgdKzFQjhwdatRLS/NjJZRXr
OzL+O5i12NL2rZKRXdmJiWTF/4HDmLZC8pJ91fENCLR0Wg0QjXL9ldy6EWUBmc18
S1WCHPY/jbc+3AyA5ejaB5swkQpSyHixfBuckROm+5U+m0EDT1TMNCVj6Q/1aJVQ
R+4R0hzqHxFd4/kAX90La4XdKuy7KZCClWA8S9VR0JZCtARc0NzRKPQfVUhZlPgi
nlX5RQnTI4kg6Ap6CCQVEuTDHhwwMsdbPLM7bTclRRWKz6wrYhvplW3DwQei4Hu4
rfOC+0FNVIVXVKH054d3sZ0Lv72FHpjvPmmKEOmFtbP9KJn8KQOw1LfB2toPu5pc
HazyK8dFR+EY5M8PcLR19wImot869bWUblVLCm6o1QYX0ltELOnUUVJ1AiTh6gSL
W2ZrGRrJtYhn5I5BYaDCyX7gJchI6h1CmgQDmsCsfq7FwOcNQeorwUXqqizeTYLw
ZnmDu1gZRxBTbIB/BposEH4S6Oui1U14hdEwFfwnnq8dKzmX+5RDHTNPtJzWlgFU
tXvHkj8lDJIZdctHXTk5r+J0RqojF5rupx7ZgjWvn6Mue2uQeb4aXzxft3dG1dJT
z29DtTVCFjjMPK8lHAwqjGaD94IVjK7IU3xoHvUK+gaSyJss6pd2M4PuSCpL6LMD
FC0b2wG4lucBn9njSMfMH8oWHatJTRp48SBd/t5MTcjj2nQchgZRniMLuSpKX0xc
/JaJfQASkS1uK8fhRcTCEns1m65bi5LRA7tSyaycfzz74pvoy3BnFEedsOIVWSPl
swP2J3ZZOWYkzBhzfYyQ5DNE/AtSC2JG38BqeHq9kzupRTMAA7I4gtidoxwZ0kQn
wHaZWHeTFq4FDcPqZM51Uf8LC2BbTYcEr5fZSHIXZSGa+QuBjozZWsSQOPhgrJlP
znNqSKZh00yibUrORmlP17SXQPnKhYGVR/qveKzzOcrXR2tddVvlkt1+OLuWgKNG
PTN87yhZoPrEPVR1cdNJqJN9vFXIOdfHrXsNg8OEjEu9vJG7dxejCaN8xaoPMdOs
3ouCrGhFu4fDYvz32CkxNrI3OvOHSd+wbwA2uuqR5K9H8JPpYU/HhhUGmLWe9wtF
+cdtvB8tTfOOBbv9859LX39bG4nRGj3/vv5P5Mx/ctmWuwsHRrSnBYGPBg0GY/Ni
rGH/rOl8JVEd+bJ8uY/uWtT3fo7fhdqr++GNgm/3E18A10Uv9HJKUM++pZSYsWbi
Ezg/hDuDj79e9/UwIA3I78n9n2KvmzBYRwa55t9/CcF8IIAF7VpwEEXA5zh3cD1w
+h5YplqhyTiMG6XVL/C8jfNjjHQgxmFSrk+z3fK/XkecRLoI5aXj+G/YpwELye2l
T0p8giFU6jj247Yl8qDq+ttaeqj68i8+nP2t8pRJPtGUua4yOmPcaqfjz8lO1+0o
djHcIe8jyRdZqHtCCG3LLWeR77KALFdgdycz2URC+WP53rC5gNXt8DZ7jdgZ0zPk
3PPnZ/cg0FeGKeo+rR7LDp0ROo+JbWjd1gsaOID8Mq06T/4YApxjTvSfPvlopuhL
gCN2rEiVARQHODgJ3gmITDvOGRbZ1pQL0oKDRQBIocF0ShqXW8whCqTr2m/QfL+N
mlZabT7M7a3qUGT8WIiqrM1E/i4NygMkq8z0rfj7C/aje+JTtyRhw8VgAflDp9HJ
CcahaMpipJGktKlqWC3cRm2NWlEwNXfz3wozp4wQc313tXbpFSNav+500tJq4cXx
h89Fb6RSt0Mvf8tk2BDChW3YrrqCvmwRE2U9MJ9kGrHKDDyWyybbzJdFTeV0vDGp
lWX0m8eUvOG3fPApECMaR0HglRJ6wV05r8UvQ3/3WwMxRUGz2PM8bnBPqXHuovWn
MzDC/pqRSq1w41L5ZioRjG7/vsUbizdLwlfTC1/seQPy2QOk9VgYvuO8hdbkQNVH
LBNnyMb068qbG8ka85RzVFUZ7RY9fn7Hxm1Whc37xgMroOE38EEVf9p5Zgf96Eo/
y47JhoAwp/qMjZbLPsIYeB4PAG514KQC3gtsoazcdWW/oumG7ifZcscNHkmDimn+
G5rjrTcPQxcoqZfzIsDjDFo3U4X6ScxvW9WZ//L801knLfbR0HZteXSdwh1x04tm
g8BUAYACj/rK2H6P1PwVWiBmj35XXKJnfIVjl0IhjbbZ41J1RJ0FISblKShD3hMo
BhZ3doOlgg6xY9OzKtEMODF7cZv9BN/pthp4c8sPrfJE82yVCgTkJv5ZZRUYbJ1/
gwYZsfja+wUaHA1hIFjrjdhs6wx/Ltgkcmmz+cjK0h2j3KzFedyVLXk5ebDujeol
aoy8Lpw8iRXlOXkNfyhFSyXiIHCCjLJQjFh6J6zgmRKu8o97j4GP1HCdICc/BNQl
Xt5J+iKxEXYbNM45PztH8azMvttd6v5vf9aiVNmgTsAzR1x0LPjH0LO4MKvc4TLk
zIveXYFqpm8pWjBbfOevjBi/EeYugabqvBMdmqq3mqKRUHhLJSKKrrpPacvPP1CU
mHiViwc/fah8o0RyZbWthG31GyN/uQMbyDlF9DGE5/ETl0uVJtWMScgX2mmGZVB3
4x8if2q9HubR6dW8Uy0trLwm9nhmI7fI+SPunNmRDJnl4U1PrP4oiog8W+4ET61K
0nL/kgi19AXADA3ElX225iI8SSBgalyUgkBbYrnRQHrAu0jRTQwQ8DZzxOWeXLdn
d8qdiHQKdmX5aJZqIWobte4DpIwCUXaBHNP16z9sJw7zWfygRbhFqCN2RNFxHszC
dP53SpPALRzbdWfcNWzCjR80aHS4ubRZhpeIhUhlTsvcCkTKwhEw5laZDUgBGTuZ
S883NKffp9bEDO3K5LMptQbZ5TnAgc06qYenUIb8vL2SguLkF3ApaiJgXnl3ECZt
psgwfMqb+PAsTgYE/coabcCik4ozg+J0CO8pWfW67Pdb0funjD/T5k4KpovaccJv
Z60EsQnrjFmkDdiP3YvVkFuZyyX6g+y20YOkND+xdyw60jeAxRLcP9gwAc+tvDAo
c0lAG/Fuofu+KJPVYYnwlYua2hkCJBf39I+WdCx2kvoOd4a77yGxGYazvp6M2ZwF
bjnBpKk+HD08dw2aXdr69k9kIGlZNUw1YsAx5ni7x80goW/IPtGrcjWPWcDp2Sbg
pwnJwjcJcJ7M7WSrdMaZrmfhaUdq1+cc6fGbDDmpDFvouCJklav8R4z5y/HvR31G
sZxx6d3E6tWoPb2RUXlR8EuHjmtpZp6vn+RG7L8v9APu35cE6798GAS39ZvpPzmZ
hitdES/voojmHtkEEi6myCmj87yuxb1xLdM+5S6qFWlB6rkZtBv/IdpbT0mGR6Q7
XKIO3itFP46lCF3q9i7pW3hF6/+DNuVFn8EhPCv2EUTU+XRpjRAymm4DWCr/Voxc
YG2W4MrhzB3Y99YDX8HVSACHAYwVXRFTKFFc/Q1u59D3DY5bN1g65vHLuM/M1F7a
bQ9MbmgA0fQuqpM/AwmklENdHh0n8+Qk/6/N6Sfy2ff1mmuNknGpi/DE1JaAsLVj
jcWIaJugIGJeLXiunsjY40H+l1Nqh9oL0xPh8tcoSDdtLZDXnL6khsPa2tCUPiol
JsFLW78pvkeM90jIxT+r/7bSyoMqAl9q4A0gceRhQa6lkAmF+WuRiPk7NmxDbTIk
LKiQF5YTKebqd68jUDz20o1SSOA/jKJlXprqI+DhGTNIeAHyHNYTbHqnmSLYSFrf
WsXC2iDOnLWQ732ZNxeoYTtNwMtci1pqsdVxgypOfjQeHRXIaLLC9po9hukw4gbk
mEo2qDxbcAglB9UMxCWl9mAnKG7FsVser8ht7ZkqStYrQnCD0tf8GrBKHynRF8Tq
h5Xe/edl2dy0l5dEYjRiupVZOPYRKdcaSTp1nNNF09wNmOp3vjCom7kpgw/X6Vec
jmErV/l29xO3yH6arfyaI5kzlm6seENNCGFJn8UXYK/NpVT7HnatyMDaMWQkK6U4
DQGg8IQzEUlM3fEPGMQvokZArAxXAiai4kOxmzW2X4fCHoevHrBqDKV8LUcEHPY6
E9Wo8QFr0zQcWiA+KnIk7Tr2CrRkGUfvQg3j92YFVWWn4pjpZYWE7WecjuIL7kyZ
p3MiBo6gGUaNNCXpH34W91to98wa9NOuPMEFGDVl6/fxzqWVDF3kY23xCzIXCz13
dFpaq8a1w0YzNafEF0R+VzFLyKWo+83LDiwm/eZvyyg+/LOdr53VU/msybfdGa0B
06Y30rk3752E5Q1z5TFC38sreNSw5x+cA4QbrtRQXbkTZTcpfiDSnUbUEF+9OWXW
Q/NNo8nhpgkFgyLsz0GJZrnvbi0pGcI7DDST/mnloAo5trYgjSsWDO6BDb5f7htD
lECpCfpBDmSQCan6hucrIWoMEnlcRZ/MmQi4rGMMKaoX52Fq6U4Lv37aFOeCmHrP
JovRpvxlzwIGF4QA0T1MIJ1gNP3enpE/Crqq1gajgRcP1SdtEoHWEwkqEoOsoy2v
l9G5Gfph2jOz7OkSSGMhyZUC08QaJuhdFes9UDuKvI5/SQhpMF8WmNr92XONllP6
pBz4rrlYus4VTGtDbbD/1sgJArDdfdreTdrwjFq3yqX0dewGGxWdA6CjsNtz1Icq
GLpTsYIXmO3NzURdW7VcPjTDIwM3tIIi0RJE+ZmCy6MHUazRabcOh5zbHam0uhbM
PnNGxl4R8VrXjUvwhQOmtkQ05/mYeh7eJoRbxVzwhCHDbv/KhFdxBM0/lWVoYJ4E
dZa3D5WL0YjYpkdDgOK/es1p+o+D1fhyol2CdmmQw3m9cgDgz7906MOizVcR6QG5
oLesWOnHO46q+6Cs/lECKvDiZAGqw8LKT6eRqAfNP3jnPQmAQroOM2hNjh50CdD0
a2zG7FbD+3+EfnI8aYut0fFh5OhLKsQxRclzLP4bBHHCNxPbzXKpZwttiQE9585i
dLy4Zq6UFFE2NMbsllgwYR9P4Yq2XDLnFaLl2fZgEYoZFfHejjWDl1rpIXz57Y1L
J5H4NydDTO+GEAfNOBfYIhJQgz30Nu46xn++ZnILBVFOBHnU99TYxibNXTUunQ+T
hOkmsSoXWh9S8ea5vpZY4Q3g8nQ5XXNB0YiPPVP3mf57X5rto6kmexdVVq+BN4H2
/WwthLCK6v2B6P8+G2L7T1d0cwLANhZDs+iQn1akHi5DG9BJd1DiL1iG0ULwWczl
gPR5YXse9kOtdYKJVwRFJKsUb7U+Ir3oaeKT580JYwsBIHpejlm4ZD/7NWZiSgzi
nwfisEtwJdu4OEHunUJDiK3Bz/8ybFyAMhTtS9SMqtH4ur/M3sssQoXZN7uH+PZE
zsvotZpZBz6fWyzI8Zuw7Rihvw4PFqutGisJJXMRb5s/apcJGJWKxYK9heGVClIa
QQNvyyUiF9zIW/iFzhZUWHu4JAxuBUEfXW3mYoTBxz+GKqAdt7PGa4v6BoaqiXUW
IqqRBDFL2rI3WoH3T++KFHTSYtu2BrcDUk8dJFsApDpSU7dWWMMNtJS8+VExvH6b
CKsnIml4I+rq3c2eyfO9mx9ejz561Oo0aFwOGn/6cAySptoF3RmBjKFBtCVk7+bT
iOVan3BkJO47FBdxT5iaVT1P2PwpwzWIF1CpBkvCdvlelI1M7fRYjXQMPTFege+b
rbWYeGggzN0664xJGTNrTWapKHBxdhSq+tMvVgIav2ai68uH87XsR5AtCDa1ZTOG
AtKOKx7Ku4uaq7v/s5bX4saGzb8BjXPiElwS491olPT5oTt5zh22b/oI3j0fFXJU
O/vue5XPv6Exo/5uvYxZFU7hqJ75G0XtXrHD8pmTEKlwl1weEkoh6b8/pccEaaVT
7k9uXj5OIAYSWNFVdfqRtHmsbUKtV3ZxcxWK7erDQgRRJHFCeX7wKo88jNHeKR52
BmxTVJoZwmxm8kRyBf7lUb6nURtQBEjmc13OuOaq0HTstJDpLgH3j2cYHM7vBq66
2qiK+yb/eqHz4gnu7D3HIwbg8ksqFa73ijLl9cGkYOfXETaErE0bJsJaGlCUP2eu
UlQx2kFcCcxKtoOh1GfAJNvd7dEueGZzZngjJ8Qbzz8DP5bFxvY9/Vn6At9eF+yC
pcYBezb9LJmMTdTajnBrpCBRTY4obv4xKxK3r/JTcJ6LchrWDLuwpcf+5iYH3hS5
WDG8hfVnUlVGP5HK5/7iFAod4Bna+IybO75RnMpNsY1G58df0jP434PSXcM3GebE
pNCK6sN81gv/On7+Uqh35gzQmVU0Qrcou/JhmYPOQX80CS32y+Ep3ZJtPZKvAlzY
7E/JnEvqP3lOTsD8ERxxBEtCdzZvmjS/sDK20CVe4JxvGlnwQp/xzdOxzdsmGYjB
UXXZXs5ykFBsy9o1KkiDLsWvBxQMcUPlE8II770hGsy6u/TfmmShZnh7GdDF0M1j
Vqdm/uN/Wj8kV/+b3g5qIw/NDV7pkANxJu3XAEaP+lGe9TBlmQjtO9L8viSn54zr
e/y8bnJ+l37d2X1JuZHp5xbEpzhqW/Ra0fHuFj3+ahnQ4Bc9ZmAw5yqBUn9bw1LR
aXnGizcjbrGUKsq6OQIYkDjUWMnJq0YymR5AvLVSZDVCQvSQ+AbF4zim/UuxXx70
o/zT6+r2BC/ryTKszhaNGi1TjHQX/5/9AFQaY3Ax3dekNFDp3b34TUNvK9o7aZ7z
L45qale5IuRV2aK3pPO0nXchDa9iNeke6aE5rWYPed3ATpltHDVJ+nu2IOWYP1Mt
UKK1nU1YSkxTpsnVexsBlHjaaCmxok1cf/KUTPYUyp5luWPRZFsJjMde2ElaQ9Fk
B3htP0wrKXZzDxgn9FaeVngmOvD9IRpm1ijRK5JMXiKI8CpJxZ1el6GJqRYER1b3
bVKSI4EIOjaYkKz73vZ3IY3ajJzJ0sWs8YuXgDiipbppwUFWeB9FtgQhAKIE255E
WSCXNsQpP8tXHfFlQKa3J63PVSWjdHsLeZXALQgKmcFvi3fOZdHMN3khhog3J2k6
deWzohzrkCBBOgKtoZVyH4p7q81N0g4ZzkmP+/CPjowkUrDVVO1FQbd9LYeiUVyt
xG7ofdb3T65NHXmXofT5U3I0uwRX7Lsj3Px4K5zcsJUrLKJRCfPWWFTNU9aRLgLM
2VGlY5Sv0imqBn4zWXBjXS9Q3J0DQOGTtDGtGXAvko20ofMs1Vzb+binXMeBByM6
rOtIL6aiBkqWKMLkfTt/H/hCEM8+J7EnM35/TR4Rk40wBf0nwa2RE7zm3fdGd+X7
mSS7sGjDuxzpKZen9coE7KpddseXG0WLeauif5OYJx/vVCosyucOvIUHSPXUHe05
Cfm7nIqjibTI0d0ns0G3AIig4qawfZUPA/h65SOygQSqZdOSA+E46iQ7hJd+so5D
CV/VXRLxaxdovGY27whRyrwyn5WkvXP6kglasm/yJv6sKSduotBnrGmcA3f6nljK
MPITf4Cy8uL1J6r+p7bh28avmm+ZEUPggtkZThdi0rnUlbgK/BSiQAt1zLcTn/x6
kS2eCADd+aRAUMmKlrkLy0W1kfGQnqntNA/oBoWmp/O8tlMwnV4zLecInBRts/e+
2QlSXiOcQ/3Z3CzbR0hNzL371LWa6GPeu4NwIHV54D44aUzw7TUR+AGRo0e8noKl
m0SEAuFUdR0d7cDBAZ0LQtqkbE3TkTGSvxHA6KGXCW2PuggDGjNBuZvVl03KYECX
cYSa6SMm7wbGXfis6OomxFnqD3PkdLiLGrewse99IQgMWLVEGKIlUe8AUcrzdcdg
RV/PelARhzla9U0+/DBJGmRywJuKdZ40L6UoqsSBC/Ew0tba95MjJc0MztExDBw2
psAft19W1iEk24eRlZ9aJbM+pUWVsknNuJRBPqgOLgAVrCojgd8oCwSINn+5JZUv
aiAHTNvwNtScxzGEpCl0ez3vPVA+zy3BDhx5OM6PPQBIWzVZS+gV77OgspBzCldi
QGDhoikyYqnlXDNc03vJA12ty6wLqjXIEG1s1hO9Hqt3YWBchFfU3ErJCKxl7hDO
AnbHKRKD5Ux90JdJ8d05eIv4H4iLq2l5kgs94ca98cqb1jG1vSey0sgel/ipNdgy
oZ2hXvxtkVfCraigwaW7KgmgOSv2L3GpCGHfuJEDeQxFHR4pODEypnFSpBgTq/9n
+5IiTOAwJg3pA0mIb1DC55qmwtOFEJythGZY3SSctZxvoDcJY+fY8+6aCOGTN0R7
TFC+r6wlH3G8e+0Lmt/PM5kh7D5AJYK1Ce1OgZtMtcauqPca9rHtrP1rqcodHb9U
Og+IffbbQNXZg9/lSWlREtEVEaXbGN//9olsqPpW7oxR0nYoGHtP2XpvvyLrhBez
8NCy6rTbFHscjFJUtk9pvgWMkVORL/PgQXcj68/gzXQmMT3uZlZppqrxaCufjFeN
q0J5gXd7LTfBfpFc0y++DI9Y/BU7+SyBY5iI0Vtmd23QBzbIXbezJqpLQ5M7e3ac
JZzAAQsTBeuY3tDvCJDAWhf3n22gQmarxplCGROHWKMbZsZMSC7WX/4CpWEkq3oN
QiwTPZd7yMhc0IWLvNFxiVPBRVFMw4wARZvFO3Dyye/hsbPlPFRuu8zUhih4yr//
oCqTDkNkeTXWCTK+tVdLvbpnHqz9nOWWmihh6jKAQU6Luoons2K0Jv1HfZcGWH/a
k6HaZohSzZO1sSm8fUnzxjIPD7P5j4wh/6/nlEQgT6G5j5RmZ3cIcWhN9LHacqLd
XLaZ/S2scEtjsizX/PWE8vv1txCb6Nvf9RtPCAGcQMcQtV04m+ZbUpFd/gIoNUiW
Z60PI4agWfqjoqGT71SXlNfBOpBXUB2S0giF/T/l/00dfcDfjNHBUN6cqErVs4wO
MGc3PG12l0AgeqM0+JNatuc8dORzM3t4Bq0JwBRjOJjYodgYfZ1qfcoQxG3xN/8P
2Ovpa0NuzJu9/PGa7HMI0SsZyBlioqHzWwuFZYdL0GMiZWxK5zH2f2ZO+Sf/Chbt
DIhuq+0M6ki119pzbh0xHyPyC+dVis0WpM/tM49BsJ8eNU/8U1fSMqQlfIMgyW33
xcCr1VxMMzVUdjdlCaYye/b3euFxjk7pLOSaxFoOWOyl8FgvVvvm0AFxNXsiUkEr
qLcfxBqmSMdRsPf6Yye86HslvFiiwllRR+y3dvJxNNPiEwg7G8u/ksGu148EFcd6
+FtkIzb7oyPubi3GjXcCxRUS8mSuwk/CKqP+YnZuyWaC+PgM0pdQfMMC5yw9Hu2d
vqH5d0si9rAwVNIn60CCAufAm9DXfiJV7rJNUOEyl31zAm3Y3Ze9hN0x/3PgaEib
RwDBIgZFTCBvUgB5LL+HiLXnvpUfRjmtAKjfqSFjmgPLEp7BqNGidYCnBCNUpnG8
f1j/mIGR40nTzlASUz+J8AslFoJUbwySLClTWMxJoNI/gryeezejSyOIVG1khSAD
85i5zQ1NZI4ZeNdEL3bF4ui/Xq+kaulejsP7TMI/i6iifCpdinPiUU3/sM6iZqaA
nNM43CQR3BGtKGu4do0ZLPUDEnX3eNHT1uI4iMGPvKlahY7238Us4sSr2LJVEqe6
kddAsDAjHpfSFzHLBL0WF6fXbRAKcEffee+h2d8gCOpnxixITD6xDnReBYPMZ9d8
LaucWJGzTmePIESsseHT00LCBAzu8ztfnc2jDknW7GyG1f0S7T7TYtCO/s1dx6RH
Sw3oW4m9suR6cO7ytnn/uAXwiYEiYSH2ouipjxy7tvC+zFv2qRqeuJ3S9m3N6cj3
4GinBVP+dm1MDxz53TsquBIv9nOtwBp2lFe54Szmjk+3LsmPl2YKQ19QNDcLk2ho
Bpc5N6/gJXRfDNkBoJtZsgxhIlEHyPsdpoc29WdEKyStLpDfTJ9jky1fZNhPaN7u
pJiJDONYOl9bDG6Lh74m8d40rVK1RaWILCP95ez/NQitkP3AE8vhZoqJ75TcLRR6
dsss54Y0tsNCJASFYLJ1+KR7AyYetvKwFJgBYTMI3D/+wXfOxOwLHUPwpMcOT/K5
DVnCTbR+0juW2xuXv5igZRsVRSXddLS+fG0Ozb3nxy+qlj6HoYtl4rqoxJUzZhMv
cj7NBrjjYx6PHrONrdM0yd5tTmvH7AiSdguWh7LJ4mRWrqGChPZjYAZKf7PGHHSy
aDCyTL/NNzabqY0SIQMUOrm41bv+Gpt3/ad3jm6paiO8yOXhrqg8hqh40862WjM/
/q8PYUr40lN8fjFoL3XIYOW7myfaRnaevv6N3sDN69enR32byMhg6dIEvSYInqIc
UK3DV+dvOAWKjolUBXpkTTfOgWr4FscfQ6GHIt8i4W0Ch5kOCh0f2JEUq1rp1hnb
6dBoEHNWKBxENxezMoAzI1HSoIwQtoFDZ5b3r+UF2s6jv2gtV1faTXpK2KNay5Jq
rHsCBgIuZv9tg6pHeh0T3cHeQM2roj/2FK+81MpPm12vuJz0I2bcUiKM8gYdjfhl
IZzyuXAy3U5dwc5wx6bN9v/qHiuP8zOmp5xxfu4HagfkzR5Hyap1aIg4l3lM6HPa
9QZYQeryJ0aVuWrvPXXKNIQ378aQ5NXK33I+k4+o5qE6ycp78is2f4S8O6lzRtnS
mxES1Ig7DX4HrdPPsEdzeylcIFTt0T3IPDMd0AAzTNAdMazpOvHQQbH6KLRJNC/z
tibhG4+aBfldIF8ZcB0oz/nGDtNMO2JBIWPVG4EWDxxHzxAVaewDyXYvWKsDrZwf
kKGdAUAASMAJK77XGWJuYGEl3FwU1qk4uNZ8xC/tSl+cpXaC2//x6yMKvr36/MTE
flhgDGM1aIhOrPsPg3cJsdMbENNGWaqXvH5KW3GPexI8FbP6qeP2sjj4VuAg2zM7
MWBZatgR4dN8cPKutQR+XZqHHN+ZLlnETSg+YGVNvZRe1PhCoJFi4zAJvtmBgBzM
ncnxZMX+iDkA2DiFh04rUZ6iRPw4/6U/97KDISQmIWaWG0s1vZhKgZCMX9+Gq6fI
kzLPsNvS0hK+XxPFpW5qYCjVwLyBGDwfRxEENVFQNupbNe+FKemA0s5Hy+cojVvN
wQy3rI46Z5M+1R9atty8BVAwaw5Mfml+XDVhPZPeGluHi7Lx8NKwzwVZD7QcRK8C
qxkYw/LPylAQsenkB5dtyKGG8UJkEcT4u8hcTcDxJy3qgdyJaWm7Y25eDxPux/fq
SW+7Jxg5jkHjsGQaycH4rPY+YQc2PkHv0A46QPvRGs6oON9FOMVu+7xiDHy67pHe
R8nTTZRKy59Oq2fXD+ieutRoGxLayf0PUL1GI6YVe5xLwt3gEmdhVHsb2fNv80Tp
wiiJsXlUR3ovA4Un7dOkhJsbXMkSgYVtg5+rean0iXXq8WMn9eA5+eR0PFBUCfLB
FhvtBbHMtRYK9NS9tk9RwgrHTFOHTCxf1/cb08Pl0+R8cQeU5Yl9WPRCDCFTW4Zo
OoHj1HbFm9aYJffDRggH7GMjZMNWvKI20LfFCR5FtDJsDWzfAv67fbjFF0Pxdx/d
PkcEN5uyR2FC5Ue6kpx67KAW663pWoJb+/NyNWDAfi1mcQ7jW8vCQKNjzbTm7sf3
F1/FukYvWoCGAEuql4w7itr3L6vc0trSDo87RNFVA0xk8qh6+GmUyKnexHwgWLsb
dqwtseplTCKEZhVo0smu8e3Q1BU8/I7zMxa7v38mEHwoYuKpLGu+UCWrn1gDPXl9
hlY2TAPadMZ0zDDZweadXPOu6c+QnJWlvwfhMvm+TjmILFVJhMoxGaWXRSgkbscd
ElipPJ5SEjgdVwsSHbzEt9WLpmbKyfdGcLpVpN3FXUxjJ5IZymGPw7EzalZ6Ri5g
s7+mvlBGJG1GJ+iPyk5SfRM9/8Vub/TS8CH+GtbbHhtVp/arhDWWN3zV5RaA59U4
A1/e0zEi+i5AQQ7hKOV87mLYouvy2MfAqK/YG8OxVuIrdFpNMolpA85Z6iagaCWA
YmWxma8f7wR+7teke66whap0h3mYXD8cX+ImHjKURZQQcNJHbCUi8/fnGYZ8DX0i
JcfD97LwoJxDKO9rogdsbSf+2cbndiNJQWWskXptq70VpARHuoarBK7Bcn7NG7Bt
wZpRjHieRZUtSUmASl2N3U9PKO/at4h66OwoJmZWjfH3FX7vdqXrkxopkYJBtZNP
33JzTGdveUf5WV1F+iS5TILkk2VETOki8enJR3hY1dJRl/zVTwwPoiWFJ6VyqqzC
0D7HEueMWXqhVW/lGsfZO+Zjj5rgDN0OnSsiKwfGRPUOnzJwr6V2/zkXYbgCWeXE
EbzDxizh/6RZH88CY6hyYigdM1Mmx/FR4sDotU89L6Da97EGszHY3SCgOe8p1pe1
XdokqsGH7CMB8zRlXbWuQLfo+QL2isIuBgRHaXlLPuurdsQmoMziWdOwVkoX1wKu
X1uisDIdCycksFK4VJ9m4t/54xOgLpA0NBzFY0wzOWEhdpAvaR/suiY7RNEhJvG6
jKivy3w8BD40swPkyTz0HI+WERtJ2ICFlnDNW/BbvajDVxbkbzQ9hoa/VO7TmMfI
39nIBZMDXM7LEKhfflzkjPLMA9E2pZHEseWyoCYMPu5eQNpl1L1ms1Joza4+iMH4
d1FT3b3Rx+iVQ04LbAECfU5Z9mB+EB8B1a2xp+0HhZvzhJPFG1ki8mtG76wdQT/1
sDRLsfoElsVTcZTPiOQFhg2uFsQ85WAezen5KLG6J7r+0SQp8rrLCSm2YkzKeczM
uUgQsmQJKieCymqyE+FEm0qGSbddKdAUcF4GKbJ14QCxNH9eLlyhrBe/MVP8An0F
+B6XQCSrOPFmVJo4vV8xN1ft05iozX8PcIhcFobyEqBYUDAz2lybZX2ItUVIdMcp
NKgiUoe/xAmKnCbcZmpg7j2+ruRUFcKnUsTtKJtIMrRB8k69oqeUuWwf0LmKQTBW
YYYjp/wgkh3fVtn74Acf9uyTw4DnSd9jjiv500sCCsXoxe0rplMAKDFego2S7Dyj
yub8NOTaV1cizmDjLOUPL8WtRF1tja4ZKMNbI3q5oKWGQadbUpQcl6vIYB31JNmS
Fdr7hL8PbHyBtKXQt4c3wWUzy+foEWLuftBXJ5Dtsxb7OFbwH89XC/cFtQMUChGP
VdyGQJ5f+UtaQtyTUmg+gENb585fDVyXU58LSGSf7ubbbpFbwFlPUyS/OYFtVW0j
htkD5SyYxlT0wFVLY/lhqY75JtrOtSDMh0jnfvAk6MD8DhHmKHgh7QeTpZiRsfTx
R5t7qtSvzbx2u9xi916ouuvC/WHu8RfIookVkN4CFL2OBQR1wNSYc++yRDS7anHe
kmIjKqJPGrsRv1nBODHmTbO7n3OCZLPGFP+xu5wDKpUOKBijA71gfqlv0yMpOnF8
0u1OqBbVwJNA9GoTS7PzKEC2WoyF0BsJjdRezos7vFl5eh+ME2slORm4YDozx1Gb
wgx8qENMYZMrbauWI/1oB/0TIuLGeBKC04Ht8QeDTDq8xw/+nXbuCMPe6YAxUVlf
PrJOB6d3yOfN1nIT09KcBqznDnzpKb9Gxigy9jX3uAYoW9yggltvc++ZP9QPArJb
ByMp/h6E1IwUXfqXLHNZ6lKGfHVRPuuqGkhSh7kf0o7dhiW3TrEK7u8jjmWv86wv
HF+59rk/gdGg3VxYzTCl58t43EsSkMPMkUDAk9pQ/cjtHUSTGg4i6zV4XJN1HF1k
RNI8/8PSBzta2BVjlCMyF9oIxcCL45fAfLd3NAZWCBzQ/xoNM2x3C+vHLwwUYU7H
KXFSMt2Z6dfrSDddSItGbauQwvqhJIvBTz9m3dYtISz5Ngn+YihKeDXBpJSjbHbi
1F1BNJonWc2gP6ZkuZ58KoSWGgoVk+eFZGsSWRcxq+ReEpgCwtYey4UjqHDHbJw4
RdRlf44S2X124t1AkOZErESMGF4jiFMB8OIeNBu4bj1vgl+hb13pwOnVAh4OSU2R
yUHSFva7n+E1XitaFt/D8RqbHOBw6i7JBVoJrrnLO9JaCMhH/G9R8GqS+Ed8gCYL
V2Y+L4M4pAxMNRqSzAU24k181b2CjGObYtPdowG2Hg7aDzN7l7n9KQWulM+FZdew
RG842FRLdG1RN1jQMZlkkpBBRVSAzH1JG62eoNEDDkzNVRfFiuS1YvWOXb+nKswP
NY/hFmYAoSmNa4wCuRKAKsHB7HoC1cvSBneFgBfX19/9+823yqfMq/Sm0fBLuuN5
H9F8PAEuCoID3GLxAoU9mwcGal+VbZEHdcne48BRFh5EnElJeP5u+mVGWBoTuehA
F4IvBd2W15uY+7hu7IZL/k/MlenVzwaWhOweuRJTGzhBfoRGdMtCBsh9Q4ExOGSl
cGJO+7a22w9A1qkyEbndV3vnu65hqXp+Bg01IfGpTuqox1g/jhXg5MW9xoW7WxUL
9LhY6FbA3PzKOB0uAd3HO+rPkuZkzANBKN2nL7Yfo5bVC3bIKSSXEIKJzHlRBiCi
9mhMFbJbHyaKLzUqU1X84jKR3dRFrh0dpPW5aFRp5jvRFMBLGsggN0TnG/4oWZF6
Gaep346gU2YGqJVfAHgEaGliEK6799SF1LEFeJMRfTh8kfNsPNKcrMm5ILfmrMrL
4FqRceXJo8vq46XRQDURaismmjK0cpGBtI2SXKy8tWn11s+CjRV7MC0hehHIhi7w
ksN7gv5GmhZcBVg0OM/cgrEdqOLKCailLIt1iFepL8jZPG+y6djet49CxK6UCOJI
KFJwuTcbgV6ToR0NiP0DqEhCxzGc9MseRGLV6WYYXpPJfKSsSg2FlDbp6pckgY9o
ta+nPXpRPRUGluV9G2UbVGs3Sjp2OaldNLRqMUUgMCaaBLZoRDIaMuVTuLuvdqFD
Oqt4AxHiET76OwuoQavODC1dQw0KHr8YWknyGcKkcXcO/0sZUv40VmfjKfqvRJXq
xm6izNwZL7O8cTwH/ipYsLlz7XHJRK4yUkiXtrjV9WaHAFq4FsF5ilAARZavqsfp
wOQzMsKsfMEW4IHv0UiOoGCqC5EZbcAC/Q30guwSCARe7MuKnOLl4CULtWK6qw2e
2zaUZwmHW8FHk1LZrkFWDcPGsVGo2P+YWfwSp9aGTaqevR725OQ/TbG1kBSkU4Ay
tU0Wq760rNLsSVBOrZGbXT9AeJwCzPNcgr/SfLeVXDUAIP3kZYajvtADBmKLjyCQ
y/hxD6GD5u1WVSNgcw2FQh68XvG7xqLQ/cn2LjbQgasePTmAnZeRc0hox34AnfCO
ri7o+hew+Q2jTUeKSMldl4LquPpA6KllTGCeFDuGHIw4CIYsf5rNe2prFuaF92ZF
r6YyCXmKQrBuQz17WQUG5WW58owCewk/7jf294HProHMa4YzugJjBX2UjcgFPFn+
y0wVVZCV5KPVZcQn3CTMXU+Yl84SrXbW5e32a2K4wDf2hVPCEqYEzch/A6Py78jP
TkK0CRnhO3AWWLLDZhPkod37VQQHBLdHR8Ff12nQCyhMAyFRZMBMvLipq2p9UZUb
pb3Z7vnceJGjcxL6EPdWrhspZA29IPO1sf1dLnUQY2wEvNN7tIOs6Mz1qQG33CTh
XMIR2/fO4S/g40f6i5NkGJxsBtMqKyNY2v7pkmGQzu7bzqzMxyxSOvzxe9rV32D1
TdTtx4+MWmHOjLrsZaq4Ov580r5v8ChY8+616ZrzA0wzBt+HNHmDpKY1EEDbX6XA
vhJPh6kMG28D3BJFP+8clAFRn8Nkk5agCHCM/4IiUGwnejdo9UfRzJI5aAAMwTEW
5e3//S/YsQWc7NAQK9/AsCEto2esKlUBO2+FOcv4PXA1uWGcPBoYwjRo3tl2wImD
LvEDiJyuP0pXq2sYdPE6aUaq+VOeAb3fnvpep+dxeaGroXSDnt7gsGDqkrATs8Y2
Sbn8PDqrP06IlcrEer4P6lNJ05mxjtSjvZr4Al/xtVOz3rYwtaqPcJp+Y2oxPR22
w1R0SNtxd6CstitU9+7So94lJ96/5y0pG3pBvxozl0cX19+zj5WwgTyV29IThzzm
H+NamVaNQpJwyB2in7Ptbhuh7eYVmddP9/HjcLdXw3GpmfJ4II1iPDEKtZOnkn0F
0Lt8rWfapAJ7DdIFtwvid2XtczkmkkW2uB5YhF2y4rOqgNblbpcm6S8qZ4ykoDyO
FAQ143shWLr9hX1G0SKcuEz0j2TRvU1sB2+Fji6zpw53YEJtUz+1Lcndeoxooo8T
epj4K9rKI/RhzSMi8mZtRl6tzDlpTusuudmirPtGuy0k0lsbhueJfr1rlKz37gSx
yyyuPIHTlFsEwmDvrenNMFfMFy0ia9PurpoFN1fCdSfTHRaEkjyg8iVvBNgvRl1s
S9mr/m9sanZOUKx4s4XI/USH7A0n4SV8zW9256/zQ8/R5NWE+xT8d42eKgv1pHvz
2rAL4ioydgYM+GL7i7jKBYCz43CN//MetZn0PSDxTsrF1h+yIE5640+iRPsLJLUv
QW7OiI3OHGBSVLv6rP3tAKhkrOdI/7lerCyWqdLw9HTBbGzaoUisC95WqqtQQH/d
ahLvT4/+twU3/i3Frc+NJWQUPxlcdC24mZw1HSnJY0V88QIMsLFCqkB4yu2QnQJJ
9dI3a082xAeXO9kbIUXbdppzBOCuX4up1PbCTKpJo/e15ES1wHzhSa4d3YEPdZoI
3MNYi7sYmqIzzhfXKecyk3Q4Tsz2VjEo2W4Jz+lBqMxHLmmJHsSwS5pPD3D1u89Y
syK77kll/0snEFScEyfw++ueyYt7b0btQ8mciWG2e3zNd9BBtks8RrSn9XVJpda1
lOLLLBBi9sB8c5IhLAfUdnZECaGiatoYf+87GQ9Pe9LMerqO2Lmk7k7LnWVh698E
n9iwJGRCqI0RaG1qrurT2tlZaEbioZH+jiAfTOcBzDtgWV6PWruHM5Bko5lGeeb7
eEurOdeZ3Sd2Ni7+vKI74Sm1+5M3ZaXh9pl4s6TPpukK2OdUxQGv/2nKFrdJCcBb
lu96g2MuOtbqCkUvfS5NQw4SuTwVvqWCXMz6ImJemjSVu/9kNF9/s+zgrMLEsQoj
0et40BV3LOxZdussxN1aGIjMts9NgJ4gN91CyyYIbfh/LH9e1WMPFBe8mjyRkDkM
FUH/NvnfDNYGEQKFSJ02gcJZVERM+/QT4qHDH/rNIz/xkYvPPrv78rf8W/Y/ysbp
WWoRXuZPgAmhXOy1nZkE1vFNI2QN+Obdag1r6Xl1Bym8uF2HvDK4yTkut3/eXoyd
XlZUz8i4aNQXeNshz4KDAE+XPW6WPDY3SRFA+gizDYSLKeSQPMUZxeP9FaYcED+P
l3t9zd+nF8xMCW8lvVW0wtRlq6X6xZU0PeKY/qtD7Qx9dTUGkIH6ymejdS0aaFA2
DGxfvxViyUaDMNeRx8XS2nEa/1v16QErvfmi+r9dR2aBspijREcpvWGMv882xXrL
saJPoHyvHzFP0Kko9nDr7u3WE2rPY51T/j8AhZFcLcRnwv6w4fWiHDAR2hIQgPY/
jAV1KiD73shmNcqdSJ2grWyYsjQ0g2zcVS6jlJuOdVhdvfeRnWTl8ZXucVCMtuFc
lK3ZG5ZOZEifwATC6p9kTlize6GjOm8bH2xChQ7YmhXHhL63Kxde4P+euXPzTN9f
DOZQb9Q4JcL0j1Sur/s8rJG/lEAwS61bS9++YeTqisUcN690Pd3lVBxed8MArHwW
wbn2fegQt+fp5P43E5uV9+R5KlGr8gfDhKC4MHVkmrbMK71AeyNUL45ZDvBodHxT
B5IPLC++0K/LxrISzgu/9vwBRjSmr+7GBaGQ6TC99zJNAK00vv4tMFL3hJxF3juu
jH2kl0yZ9IbFvyGVlaHU0BlNPcK214Y7YoYZmUBwXYShucRqHhQpE4GmFTJpzPXX
N0aPNCd0Rf6hjmqBoOloM1+K/dP64t9LOqehW0aDlWARVA/Kc3WbcFhnd6iyxf6x
eb2oN/yDL71yuCNiazG0VguGhsM1GhhBE5QmxWLULU4PXzRoiBfSEC5MeNb6ZUnY
N8tXCg23p3oKY5zSPKysCZlfNumB3WDBJGA+TU339/ZyA9uu1/QNiYTxOa0jUosc
Sci+ZiEJGzwYo8EAX3Jez90Kqol9Ip6SezGSkUt+ZO8+ac1NfQQut8COlwSmdS8k
tKuH5BzBh39C7jgqlKo58otQzAc1M8kzr9+tMwAE5PevNHh1+MlWNkkJWw4txB/1
ppCB8ct7on3IFhQMnl8Zzzj/kQaY/LkXgNFdVfv0DRJTiXEddGJnPkwS8XiyXXJx
IANLs7RZX/pu4wiWYh7yKlOIeF2LwsGfAdYOLoLL3YbOCpzlMiHqAKg/jdwwkLtQ
HFIOxjOzLkjGnlBZ9ywzh3PmoO68OAOiyVueYoJXQuWqyYOr8xfws+v724inDLMY
Sxv3/O5h3+aEbJMWUTIrNsgfp0LKuVISMJ8Suj2Td4ivzSpJw8S2Gjzpen4KNbjt
AJ7VO/tNDGbzrvKy74pxn8D1QlLRLLko4zlqjU8b0/KUtJw4iCQlUq8WI6alMBvZ
1K4EhnkRNkYv8F7JPzDiD0ZRjzAGitn9G+EZQ6PGxu8fO11gp5kxrcOu846O7XLv
ZIJjJJtpJwok51jMHRXSqsv0TDR3Sb596jEbRwJgIsteybg2VNAFaO7BlM6P/17h
k2H2119iFB5XoSO5YaatjK5YTupT1SywccH/oShfBuxN7hKAL5NEXT2mZnqvAh+w
NoyxAo6jVOkeXROaZpFcBUl60T3sTXTAa2jMHL4AnlFIX8ScOlu7s83lljOpqa70
fISbNeInRZtVdEe149ZeMBqpYmdWJ3IC2EPofOwlI4v6lzYdVhEp/gBKj9xS27Sx
AeuHCKZ8cq32tVRMJ88HoAmkLTnfZ3Ns6RIiUQ6rcsnTJAsDfnE2j46gvN885zCo
1oEjy2Onh+H5Nhe0qW66JrhBQal68QiYu0dJcY/YDOpPuInZij+1Sn5f9xnslxsU
7V8PpR53fcfA0UFTWYqCgCYTouDJQGfNP0Rt5G7s+to+kcpo2esS1e8E7mXp/Ni0
cADanKory//DAhg2g+ecBY3avtXmC+JyzpR6CcnSIiHYXHj8hqeUEBh/8mZoF2pB
ytao+qhaeXBeyI6RHDSaGuA30BYze1H5uUlbiJXEA/0UAS0dm8kMAGMxPsj4NCQB
AKLOTzes/6KRBjUaDYqgY73lBTsj9L0DKxRRRDdH4ehuyXeCmnKLR06GLBFI2A9Y
PbdjXrc24G8AfbBoIMrV9/hNuf/oxvKZQCouqYGusGsr3qEENxGXZ+So0v6Fdod1
FQ6MBDW/ZU4Mh1+oXwDlX4uxs6BI98xNvV/V2kEuv/T/SuB800C/mXs3mkWWp3QL
lmniRfPHz4mMoCW5cyjlG1yHTUHQAB5v5YYHKz6945krRCuahCcE39sT60R+zqAy
FLjgf5hxqJJZe+xzAkrV1cuFCjXOHPqfZg5N3XC+MdFxIEu3hBTSePFjNKz7vlZ7
pVXeZK3pzddkvV1aLmrZOF80chF+fvCuuXMH+L46FbWs/GR8LQDVdPgrnddThfWC
4qqWlbgOWJ8JyITlj1cOCSUAhiE5xiga7ut/sIJ9j3/F49yjn9Pg9WVaK32F/ZLd
c+7CH0WdHDYjnXhNingHigQfDNrs/y0pCc+g0Crd1GggPLWQfTcg+8ZntHa2zzDe
9RTv4WLvd0V+CoXA3D+eCLtB/z0nDArDKZv+qoFSpZzYq6TfdkLHwq8vjZ+h5v8K
FT9ckxJML0fNE998Dy3jReaIqkwP1vHvN5ar3rdRNm/KZ8pMqngDG7Ip803eLQol
mD2Ym56POG+4LPE5K+RIstlxwKGRwfPJD4p+TuPzZ/P1cWvRkUlLjfLJcbRrtZNd
3UNXgpgXVejN2s73jBcEusvstc+1VEHklqOIo62uXWunxLpnPH/IVkHHUphMsP7V
gHdXwe0nX7IfETTjzr4brNhia4uRy0MfMGP8MfjseaZPlHOcGFJXk1Bb60vDYYul
eMQqsd2gn4U5c91dvVA+AL09szc9R76rPE6zY9oEKpNbvyESsjlFMy6P7PT6zvpP
PrDC4iERXNaUGwyuvu7RDNE9sDK5puGFFZRTt3zG4RfgarqfmAatcbWjWOVGcEp2
ePPkXSkf92lEvsFBfBABuh8H+0oHm+n88m7YsN21FQhyGN+zKvqgsu0hsLMIeaBw
IabkCD+JA42vBOjI2QXvSB91FSeQpOHxpoMm2JVfsshBPxQcf+TKzGwPtxDHiapN
UwKKc8zLAiTr87ONCo17yHNu6MboDEDrj4c+u7WPohewaOPRgSdLjeKE4nx/P8js
fFKm+1UDdq00h2jyc4V1x2qa73J4go0RBj6vJXOCsLmBG4cdKeVyPb0ObY8xVlr9
AXSwuSZYBaSnRnnuDpm+aCa8p0caJlprvEDCP7sMc0e70w92HFuaaA//qH56wEGb
BdfRohtMKyjEWTKWEtgu4TdY+n6hFOLrtQZzrsdAfiT+ukl/qurxv1e693AlYrtx
60PvVydz+7NhRQp5wXw2TK2hw67A5Vd6C8Q1HIg9fyxLHA+eph0IxxveJWnPZxnd
gvv+DVAOPK0pZyrIDHqtAcdNl4/U4fhaI7c5IZLo4WuvGHGY6opz+KWJRtKOqV9F
pFjy55T5N6geWFmwKXsRzKkLo+geWDgyvBS+oMWnTzPQ6Uu1xTMZGtj7yv3qD5xk
Cd4UEzK0i7bC+jkZvv6hbr6lSgsd9yCb9qIic57n6WXi49Q/juH4mHizQVB99d+3
Ksuxr6zWtkzg7EJrClorL9+jLutCTOgYdSq1eUdD/15t4M7NPav1xE2m6WPbUcW7
iIRqo647a+ivAxGVr+EwaGovDrkEBBvcoWSA7xRS/JHx2r9Iv+UHd0Vw6TYSST9c
CuP3LF8lHscKSyzGI0SgXiPMDjW8tBTy1s4lGoJU+2sVpre+ZyqG2KnLkqKCfz2G
US9EHiGhmMbVn7VxeFpHWqVoOmiXklmRsAZSlBy6oO7inKjPuSf7UVmawwWBDkZQ
0Fi/JyUMx9P0jhcNV91b6k7LKTEg5UblvIFUbeQsp1janXFaKKTrZc2U+qqlg67q
6Zj4SMSif1pw8xP7sxm5gPShOSXClZwGEqO/E3VyUJPa/opXtHsTugnYTavyKSir
`pragma protect end_protected
