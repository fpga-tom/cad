-- RS232.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity RS232 is
	port (
		from_uart_ready : in  std_logic                    := '0';             -- avalon_data_receive_source.ready
		from_uart_data  : out std_logic_vector(7 downto 0);                    --                           .data
		from_uart_error : out std_logic;                                       --                           .error
		from_uart_valid : out std_logic;                                       --                           .valid
		to_uart_data    : in  std_logic_vector(7 downto 0) := (others => '0'); --  avalon_data_transmit_sink.data
		to_uart_error   : in  std_logic                    := '0';             --                           .error
		to_uart_valid   : in  std_logic                    := '0';             --                           .valid
		to_uart_ready   : out std_logic;                                       --                           .ready
		clk             : in  std_logic                    := '0';             --                        clk.clk
		UART_RXD        : in  std_logic                    := '0';             --         external_interface.RXD
		UART_TXD        : out std_logic;                                       --                           .TXD
		reset           : in  std_logic                    := '0'              --                      reset.reset
	);
end entity RS232;

architecture rtl of RS232 is
	component RS232_rs232_0 is
		port (
			clk             : in  std_logic                    := 'X';             -- clk
			reset           : in  std_logic                    := 'X';             -- reset
			from_uart_ready : in  std_logic                    := 'X';             -- ready
			from_uart_data  : out std_logic_vector(7 downto 0);                    -- data
			from_uart_error : out std_logic;                                       -- error
			from_uart_valid : out std_logic;                                       -- valid
			to_uart_data    : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			to_uart_error   : in  std_logic                    := 'X';             -- error
			to_uart_valid   : in  std_logic                    := 'X';             -- valid
			to_uart_ready   : out std_logic;                                       -- ready
			UART_RXD        : in  std_logic                    := 'X';             -- export
			UART_TXD        : out std_logic                                        -- export
		);
	end component RS232_rs232_0;

begin

	rs232_0 : component RS232_rs232_0
		port map (
			clk             => clk,             --                        clk.clk
			reset           => reset,           --                      reset.reset
			from_uart_ready => from_uart_ready, -- avalon_data_receive_source.ready
			from_uart_data  => from_uart_data,  --                           .data
			from_uart_error => from_uart_error, --                           .error
			from_uart_valid => from_uart_valid, --                           .valid
			to_uart_data    => to_uart_data,    --  avalon_data_transmit_sink.data
			to_uart_error   => to_uart_error,   --                           .error
			to_uart_valid   => to_uart_valid,   --                           .valid
			to_uart_ready   => to_uart_ready,   --                           .ready
			UART_RXD        => UART_RXD,        --         external_interface.export
			UART_TXD        => UART_TXD         --                           .export
		);

end architecture rtl; -- of RS232
