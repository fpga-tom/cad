// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TupQS0dv4M4aRkwiZ7xnIwMVz3u85OoITJUCSLt0srDp4YmC+/FHMDBPQeaG93+b
KzWNeJCTQE0ZCp6I83hfoxraCwt50Pg5kTOhVdHkNEH0cOfWnrp0Z4VZcXVOwCH0
yKkDWTwwLHCF437Zd+UgHzyZ8skWEL0QoZzXxUqDsVU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17984)
3E2BNumxG6GLPk4+6CJSLhieD4stRdYEsjTnryeGP1Du7dFVm55hXt526KASzsZu
3fQFkS0fpBE2W4FZ+NPyrSRMyEGLJjMfw+tiEF/L9CJP2WJKVn+9TU7Q7KcF0Ks2
Z4UbLRICXryLT40BgKBI1dwRBvnygymA1IxpugBNrq0FpdQgtKUto2L50dj0ji/d
1X3t+fGQ4EwIObEBpqQrYL+boSzaX2bpSfMcSqr2VxYl3tUlAVU5SdwHOIAI86rn
3UaU4CTxoOmr23Jkw5NSESZeku1ZPateVKr5/R34gp+oXyOSXPXs8/PfUJ/GaMa/
3nw5FCqlwEHlKTkkdYZdJmnIToXeIAHN207tUW1FJsWRlHkkViWWFiGSurabW47S
VATy0Tws8gdHAXkPdIEwOsnwmgyE6xH22ar3mLxmdznXdRRXBrg+wZO6dTqs6iS7
AwzjA2RWxi1p7IiLcbmC+Xx+F5ZOhr1kBL48+8mY8/7v9l6dGA5YuZqBfyyZJ7Zu
u5NP8G2iH16TV17Ga9G33QWewWP4M0DHXopMfb9zEftd1UELrSmLSlGpeakGdvpS
yDa8QvOhDKBlG7VxuVhCcEuohdf8B2og0kve7OEd0IN1wUE1LmS/fVtwXNlO8RXR
TdQK14MNN8plT9R3LC6AmXMAm7pUJqJiOfy4wLB7K+Kn97jCInui3JjX1T46SdQ9
cOM+JGLCpwj7X9U/FXY+OqgGnfIKP9TGVeqwZWToGKEZ6MOmQ7iMKRJfKAlbEd7W
x7ZcTvOZFXVnjnHDBqqU0VH4TV5+nShke8md9M22kgOcHtjBz+ox03iTtv6QNEkY
i0vWXZzOWKELz9dUxVQefZPhq81fpad2Qd728CxyVdTx9da3x5KzUMqDj+JChB9+
ngM2Bn+m77KVONzsXc5V0yKe6GGq4m80R7izu4gwybh/Ya/iqVru42yWR5CBXKNe
xBQFztW/+hX8k6YaKlaz7buEB6pPkHPgmLUQABjF4k7mtL603UOthvUHc1xAyfT3
vqQVy09lNHr4nkcxdwfive8wc9gzKhuDo7stChNJRx6Syo5Fb1Ii0PEqoXtpqqGt
z+gud9AyFbsX6ULX5feD+wrjqIRAKVnmokFpNMYHIKral+2ekqEHcXUWVgJPGg7h
lrc7KAs2pqHZQ+B4aIj5DrDwjexIHXLtYYNipXqS0pY0xev6/5rJjUzWAM7dIoIW
lsV6zVPDblWISDCIilinsVpFvaHZRIcZ0S4HShL6dLff4FX4YgRAoFXIYXKH3osz
Br/wVbUSmnnDt48IRFGX4Ixq//JT3ZMzXk2QtgSOEiPLJQ9bWXdyQhONr/aq5xnJ
N2cbZAQRyLQNmJq1/a8zT67lvz349iEDlR1xlLKNZvX5DOubc+j6npo2NZ83V0qv
VUewdVRN9HF3+UcD3J/OnnZ3sqjWZB8iOo7csClaFUvCYD6Ny/ao7E9qx+LwKrhq
O0LRz/lcxZEnIFrpiIUGWEKAF5P3LzPJINMFG5DXKK/9qLb1W7ima8k2gpoLx4in
b9Zso+ZG3mmxW+4WgTcZwRgSVxJALSiz81d9QzA1RpXF2DnrDNsM7fmr1hd1VTN4
MmmQPo/FK0RWBiKsIVJ/70tFl2AHDZgvYu6h8M3w/f17soPh1azLiXk3NI5LqPal
9wmo1VAYQWadKcHTHvo+4B+NVC1M3gfFpNEWN3335J4c5pIZhJxz6KllyJvXafU0
9Vt1MX4T4CKAG5v8/ft6ZTCKYZKqrtt1YV7TSX6rg7dfaM4kFmut2gMPY1zMQzIV
sRHs0pzPnkAQINBF/b9T7CLVROpUfRscVxn09AFyKmlI6+UQuZIfowh75+OKvf6N
nYFhj1a52uzBFkZZepc5P7aGY3b3AhVzDuh32x7aOZgSjPSFt8yvC/tJa8NYQotC
6BPSD57O17UO+w31VWwEuNp8P0CD0xfdOAnNifFLw5xqNdZDo9DiuE4BX2O1WDrs
VOE0ZlVelw3OciR/n8Y+KGofDmD8g9YD2I+0TNlR5RNTHfVmg11rDo68SFDTvozs
BToqJGTOhFvYiMAYH7zEuoOkfRGOcmZRQonGfZc/k5jSqOglcYNtx6Ywz3ZfCD/Y
IXjfePcJXfrFRZcaPajjdsLs75qsJqEI/CVDfSNOtU15qPChcpzhJZ+A2Bvb09k/
zYoe/bY/ppg7UHBwFX1lCmYBmc/CfsFfl4XiHAIyDzj8JiiRUKnaexd7KYexvUq6
+pkAK8GHBOA8FmcoklXgOeZR/YlA0XzFgMMlBu3sgjrc1RgSC/H44fXvtYDr8cca
FnLGUyXhvKA/8l6N5c+3+GQsV5ehGLgQ8MOOpW5zafEOOk/e1ysjdcbcML2z5Zu+
JHlom0x5W8bEcqdcYlp5LW82ZrSJqKJJ7UpSDt3jPhAy6C22RjaxDOfB3yVaSXdE
OV80OU9QpbNV3jrTPOPoBKzNR3gRXlLfcXi7hb64JuQni6X5jilqYt5vCVSLo1l4
lOS/tQ0ltPNG6IQ8MLXYv4Sr8SqQUwS9j7xdemZHGl/gU+9dNNO4g6uEQ2oWvX8P
inRKvgEKKrKM+0v+pEdpHOmmrT/3wUPWYzyHPmawg+ZxHC2AP4wVEeSDH4ackcQc
i1VxtcJ7KbWWw7JpdwWjD97jq/VinccXFNxCVFj400GQBHrIQ9NAZyuhZ4V96iy6
c0KHfwgqXy0Jzkb28yDkkHBFqF2kk4Usno1WcEjuaLCcYTuT5EJkQ4UQuaRATKIY
AogDeLNJi+uOmPdlhkBveSpnfUfVlNHiOLqgwHJr845wmPXTsisPCOfDmjdagvRI
vlJR5BCaQW44GkQyYhnMInygPnL3DDH7T0j14dTJN/0PbNLzj5RUtsC2FKFSJAdA
7cxgUAiMk56IDrzg0HylepA1qi72u9ZRnsnRv8eIW1vthfr2WPlG6GKOkPldKblt
rq9a3XToC2zYX+FhLyyO7NCL7OWpNO8QbEwBRr9zye6KXTc6+Fgvlc52+VMCqvDJ
b9cf1PKpjheGC0b583xld8iXb63iaVRPnfTeDb86vj2ETJ3e6sIJZQmK2yFUeIn/
IFbx48rSxV2edmQc/2pK9BjWOkp6daS+c1mF3g7WuSUkvaH9EcWIdHicOyNgmIln
EfJt5mNdubeAhVDMCkqWWDAew0x8s5yj9Bo75UzdLqykoN5STkTtJXYZkN/hXiV5
qgfXX3bj0e9TSZzcTspiQPUYXF2BKEOoa5BJIRFnWPUW+LuaW5hxInxNQmhrfbVe
2PxkmdQZnMh2LbBwyXh76FjKwfzQz6dZsEn2YJ0cHxaso825gkHz80M7DjoVDhJJ
3IKDxmcqYWAB9u3u9AVONcxHWOBeroptgJZbM/BYvMp2PKnE/nX1nVhEAL4yOPVA
dE9kFnWQBsOvDDOC9DgP7L0mU5jl0z1Yv3e0oYi2/vL7HiX/TUOqUBvVMbsEcfk8
KUxQ7d2CfJ5ey/DRPgGHM8qXEiR+jCY4TR90OSq/u3EzhQfn9p+fiVT/PI4Fa1b2
HchTlNCtaDT14ThOZ8FqnldzgeD471lZT5GYVYOnRbgzu/zWjnO0KhJXrIKbtQz+
6s7aZT4cELmli0JG0axF9t1Cz27fXZCt7qqtM+PVsk3CpYOFd+Gk3zqOyfTi+0On
jWlfZfYCErQq8lrIfzLJLYCPdSW65BXhJ3uzvKtN/ETorB9XFtO39g5lPG8JDO8j
HlEddQn5LljMlxJ3umsostziIrqGrXP/QS2cr4XmWYg9BHdfbzYjIpW9DKLkvY/X
8tMQpaTJjd1GHpYmOUsw9UN3/6rp3K4Mxots+outH2ttlT/zuOssIIp308K9se0O
BLNhqdmWgV0gSHJP7GXVwJIpyMrdtTzcgTNGtCwhA3R902sjrHmk1pH0ASDmadDg
8apeuOfl/msCp/WonOBl6QI8SlwJRXEQuKKHFiq0U+WvBT0jyfps+ZDclCoILp3W
pBWZCKpma4pkod8dpyFHzLKkUemSFTU1W1X2DrVlRXhsQu5LbAduO2+TmwXHfvaR
O1oqxlOonfcVIm/ZYCEkXhIT9Jnfq6E6dThrW1GPnvhCljkkOVzu3TUXzA4fXaxk
ZMtv3oQGhMMB2/eN7D3wLJdLKH2qUfdfgISJ0A0nqilQ/28a5tEIUJQmIufbfVlg
zBQqXN9Vt3V2n7Jl3zYfiuPP/7OlhE3wPjIifIo/kE3Rx6J8ztMp9gGJZqaPmKsS
PO0K89iLLOXrnjcyEsZbNbExdzJwbd0OUAhWekEb/ky5K16IQ33vUpeTZWqlkWes
jMuXU2XRU3z/mghojda6dhBt3qaah8mJM+TjgmKCbqmvnBp8g5MEmck+okQPSfGI
8/PB2uL6E/UB2UoPVHJ7IIEnPpbuN9uai0h3S5J+sW8J/lQGeMTOOuODKEFto47M
Ejw8Z4QXL/YtsLLNQwUXGwdD4rXmoe3VxT7YaBIkpxeYtTz1OQ+Z6iMTWGFhs0V8
5lBbB/nUkzWTMjaz1v69t8GglgrUuXTsIl/ZI2cXveQXcZu5ZDS7RpAaH/++jNE9
8Ou1ps4kRT1lGkk2nU8RYcKcZxxUMM8mkaHIk/hQZeI3lY/kusFeSCmCxsK8eNY9
nobUhV2eh6mcX3p71j2HtGNOh0aNjgxecFnZXXG+p/g7PaEHJE9d6sun/AQY+03b
FbhUUZoTkugOSkeGLf+HycztqOPt0ntEjeMRn73tf3ZQj13Y43qWHjKvlB2QKN4y
K31OTVRDAvL4a3qQ0IQlfAwqYdLReP9TjhVGN+kAgREBluCPznyNDiGUscnAhZ30
K9njVW1UAM8nANYI6Mne+f6w7ldMPT6IzPKfiRch7GYFVAszi9hZ3g48fXAdr2Qa
R/GE6AIkA3+l0A1/pO1DRqBsDibonlhoKMXvdrIN+jAkO5fMunT4GhSe+qpikGRg
s1i9IBWtyno9tmCTayfRxVFlLCPIjyKG2GI+WhnG5Xq6+S2xX08WWFTlWUkKAntd
QUuFB64PROSODX30MHctrPygggft7n1LkJFBnw4Bml3R85AoiJgqOaPHji+6nKPj
scEZ7nn/H6XEtiLBZQ1VZxFDUXAklDNcmSDX17J2c7zb3Zsj/cUF/ESOZPwlzOno
6H7GapaRW7lNfEMVUhV9EZCHi3tY5R//ELD150ihmMeUjxttLo6vgUlZXJP0FmyL
RrphEPWy0mHaONVazdjZrvoh9nRO0wKmSb5k7ph5FCm6b0XTQ9kwKN1Td+rQ3iZg
QOnO3UT2sIcznCAPOjIPmOGAj9XOeUU/fsUg8a+MXbKIllQx2JaVvtL319GlPPgZ
3YVVtULKH3YtaUpiJuQNycUI20dx8rRQJ35w44Cu7CvWEAYGgbkJmtTqFcHWdYt/
YsfuhiaN4EGrg8HSFZgOWpZUB93/pG5CXk2QHxGrp/UbWRv9MnLYKpOsLhow6hNN
ROcLuDmCYXkAWL9sjZZM6Yab3+zQrqEhSk33y7T/kFyzgN3T5jzA2pFq6QN2vj57
yWkmOmzb5dCgWnVekGGT6dkURsJnJsbIRHs48/GMIe8m4mtjuvU7ahyvzjdliB8K
ZZM6ZYrGwvwlzVhQ9//gqt0U3rgN5aD0V/3+w9i3XeCpXV1Ef9myv8ZVAqolG6hU
GIyDVJakvdHxKLyi5W5DOqeew25k/wN+xfrfwTjClfHzS2cvXw+65Tv6SyjM9Fpa
8XaluZsKeJMUg/w/xQG2WdWFQ5r29dSMr9atpT+p/MAiTGLXUPHokkEUSPrl80ok
17LlqJcYZruCCR16zqf5KvSW/VdwusoOeisei3NPxMct5L1/Cj7h/boXBCd9WL7i
gyMdYa6el41vYdekW+7agPCZoXx5uJ+qWXH/5Jx2tW9TrU3DaAFwHsnpJBuqeAVr
t+FlxESaIaVWFmizoDBqg79oZZLkmlpPtTp8cXgdzrhXxDiK0LXgoSzS1XQD/yjJ
w6p/sDh/ui0FeIBNAXiteECsn07u8ennDMWNZSVOYJlgprl+ldnkoGGAmNf64wGF
n27YyNPU6Jy38022rzFGQviXm1tTJdkddApw0jC7HhJSAg8ua9KClRVcjZ8s2QGk
JJS9ZZLT6tDxDQ35LLsUB/yJOg5vfWZAEfhUBJ4XrRk9ooPcviEAd7f4Pt/mE3qg
sz35gvVsVKlwkWwo5nZKX0a4OhjdZYaxYLQFwiHlcPEy0KvIa3mbV1W4cOzkkBDE
sBmBjC2BSUA2LtoLF9H6/MWropSqlJl1mxxE0IqrOB9NpX2L73tffRovoU4ullPP
4dPZZvI13y4cmnSK3z5DnsEEnmVWseW6MVQiibY4U7NFIC9FWT+xTIExzWctUbU0
7tfpVV091RaWI4LqcZKJXZ0OA70fLPdMEtfSsAyeqpyOHN8/Bb33PpA4EkzDQ6OC
MEKKAtLzpF2ZF6nwFM34Dwd5MScMiO16QmWePbp8utfBJfDTW7gHXJOlrPmd+QyA
IZa4m6B8McuMGbVmxS1ujp0MoVCu4IMUB8wZ8utp6GoXk6FGNTWsZdv0kaNS9ERW
XRc7X1eoJ4NNqpDJFTPuS2/1G2OjGNSIKPGlWz2PnorEQY2HjIFZCgMq3DA5tR6y
o5REOnq/jFqH+qwA3XKzQsyvZ1rfiCChwtyaCe8DnZ792qUYNKPkb5Ri7yZ8EfjN
TQVTmqEDeHpt2vA3MZ+3W+CDVgv4S+5bsJIGDdxrn+BUuCFoNoqHM8k9FxNWeSpS
+kbIt5/Xu4fANedBNOAhN6KshoYxxk+1L4Jdwr8GQ8ZUjeaOUyQHtpBxyYzR8TIh
mxNPa3X+d3pJDJeci+ZcHHtM7S7ZwVvH6dT0QPpOMF2qx95Cvs+fbEJWeSakbeew
ti6KucAcIyHvyVdRFXzO2X44MPIQtucCcKLWhGVxRwyrBqEjtho2WV60w2FnJ2iB
k7az4PSp/ZHbS0ORWTLJC+szVuUTzd+hsk5UiVwuOAKst/RDVAgiE4ppAxD4X6Ei
wdTXYEzfFOq+KSNZ3YPnOg4J5+pW59iX8dUM7E5ec+sxS0E2IHTHYlJKRYeNMoAn
MDdkmdDB3GVXjoCNNSudJjGmXVRXF4jRAiTZUsAyDXyA1zyqtNS1LzyZYMtAD1AV
Fv3rCYk5AzLHSjbNsO4mPY9Vp+wDANnGAZAZ8l0mB5cWneG6qq0mTGyFE9KTuiKU
2dQemzm8LyJKXjD+dwL+VA5tQ1ssGrd9NFDLGmGSg5qvgynhyF/P9ZhvxSJDR1Fd
iv9RwzkhJH1dV40yySo6r+6/5yC3Ir4R91oN5vsSQBANRr0ZRSFq9vq1+SzJMaVd
HNPQzgFUA5FqTfeUFPGNDNblKnrRZSv0hQjDFqRhZZ392ZzyF3BXEqsN7lXhKrdj
Jrl4+AHnN0rdnzLZfY7EuaLyiIFN/S/RtRMLp7ecPMfnDSSV+O+Nrlp2vw4q6JMX
qMdT+cUR+vmRHL/GcwL09vcm0gqbcabPH7nCGeyG1yiXwclbNhDGivZ6ZrBS9QrA
YmqR/bqY7RBGo+Vne8pdu7YRGu7BeagxWohGR+IxyR5ROtv16nyPrbrWkW+Gwsxx
5HUYZAzgghS2oeBPe1+Kg19x+ZnQTl1jS356udHPf5ZMOiGtAdGjXqSmsTB+5mUX
Vs2Z6lgt7AFjJzVZrk+P2NFC9epFg17E/JNjeARHdK9jLELHlWNCCbiATwupdyHH
1fp60azK/EAHLk6VdgVlkazi/+kFk6QOf//nWqpBi4Z7wcHkyeshrX1KB1elrQ9J
dZzN1EAwL62t5BsbsrPrtx6sfbO0HylKZmSBaRnKklUxF0ANWZSEFnuufU8fZ4ba
F/vQy6SrlSjjJ2KdbebMy2KFMtfjXGIL/8vf0dHY6Ef4N5LkEBT6ZUMR2YDnRcUf
cZyBkHAU1BWBizV7o++W2cEokBvl7T+2vkGvHD4E5PFQjgm9uRtwFnlq1JwT2JEq
jf+bPCZ1HIDS5Kk2LtfqWdQG0UNyPgUYBHebIpLtpJfJrMk617s8NGoInEsAc3TV
I2ZzqWvECCg2VxN4NS1wdCI0JD2GVlLABHx5/isIfxkSIWd20imnhMbDGfOVpsEX
KhtXT6iYtAkSSTuRAzDcECE1sdQ+BF8y9F5tiYEWRi2EqrSyAu7u1LUtxuhZUkhT
eSvGoXXkkn0oq9aP0hcYXmWHCX0EQ4XtwNXIMVmvigJ1y9bteIAimKySnA3uFh2b
NL2Nw0O5EGdUev1Je0/BZuTvInjf7TboQMbKvI46UTi/HbHosv77d9M+7AIfO3QC
oLRui62G5z89Xw5XyWChG8Yr53xKm6cnrgrm9oo23RiDKZY3aaix9UiNkqIGKx1U
AuRdLoPgN1UtEltW3H4LuLEg68+o+1MpssVTgn70PZdygPYWA5RpyTsDC/j3G10i
6ZqjpDqGUsr+z5VunCiWvZG8RmsffsDlfv9DLM10DnkbPqZEPjMIOmbHtqs/i2Pv
npGzQh4jzgZD3NAwsCRt7gd+/AKi6aO5smV9pmzcQLoqA3v4wGdIiPsZaM6+Jece
NPdK3IGtjrwHWCpbGirhzqXSVtXa/M1UMwOqiQwHr7kHCiyFfjFmiAEwCooADFZn
lKYo4w+sIv+8aFcqc3R4Qld74okq+8SY2P1pjwpp2634O7LL+yncY+RtR5+Lzd1q
uUpa3o8Uqn4mNlBoFSkpSElnzxmmooRNXF6TB9KngjILS6W8UkbfEJGEPy1mGpZt
ipm2pI3/zd1fjsqIDayrix5Wzaal2aOlFK0pI3cdn3l4JMEP5g4EX+v2cfsaGC5i
o77iO9mrP5+2GwlETc+slKxdT4nK55Uza/4dmiJ8LoSjDDUGks0ZoQjViWQn2JbU
Q/j/tJHkPOfge+OaBtlL95MRtuWXU0KzNXoetFHkXgITXvyMShycPXNHslx2cmOE
v01fGhC1/PpQnQ3tgWPJQ4BbeMVzbW8y0wHg06zdEtccvY5dFQPBmSSnIwDZTvSl
AF0Tvr4ahkOGNkQxwRsc0oOwtvUQd3X8nGoKx77i3LFQyVGC6xBBfRguxXzr3FS8
RiDAeIb4grYtdI7Lvx3DopmaXZrO5r5tukCbInaTIIHhp0X6Yk6KiHoLBXYjghTC
xHrKky9XMmoZx9ulmZRXH6hEOUOYxsQ2UGdsq3HHShZ77EVmKTA4F3bjNULP7E+L
o8pysuxUpk1rw3UCo6fm2RdfOFdlsdh4lrGD17vAX7NmbonYmmVbmlYYpTMGz6d9
/bfH+lUU4kFe6we4ezeBT7Za47/4llqzBTK73mPL3hm+ZXwMVRMQToZgV3TvKO6l
Ly0Z7pLooJrr+Jai1Ot/IlStLy2sLt+oyZ98fk2lkQL9RUfeBwe2rnmmh9KwScPR
ikra84qq08Wb7Bwl8I/mQ5JkPujHURoazDADGMOvAhdM/lMZJKY3Bb4NUorstAEx
nXqcsO4cLPF7Y3vUhNEBPooeNf+R1gW1QL6/Z9Uuf/JfkL27LmUybCjvYdiyz5I3
4H06gjlFNVxe+T6XPjHWblrpgETeWBzHMzUq+NDgwFXAle55myP8qbfHEDbZVVC5
L0Rx9zzcQ88BnsnwjROStJEkHR14PTjUIQo8PhXaxEdD7K5c0gVLidyV1XFYyFDw
WqeIzIjim2BfXLFvTgR0v05wmNY9cPSNoL8RNCxRmVwSZdYUqCdZQAHXPPzF0K3O
Z7kkTSZXR5NKbhsMTynS6iP4jVDn8Ubgw6DmpfT0woQKh3cBWmbJq/Ns+mMd203L
ZRq45p+1B6EvpLeHipAHChuBiCQKLTjCHbDyrMqaoLYikTB8fpWYUPj6IRDkwpgT
P9ytrU7HYBmBTCb+x2odh55cwfs57SNsZLNqK6lI31OtF+zqzxCx5YuNvF0nSXHi
xWkIdWrjfS9eDpA9tgO1UxFdOvCEn7KG+gzlyuZuggzVu+pDlqs/FOT0oi6nkx+h
C50NnozIOpwT+a2/RuaGjoDFx7go5HRl8BP8+y6RwrY7tk4C81JOIG5VV3cJQv1/
8Jg3wDkua0PNsV+3YqpFN0GsYbxyagc6pFyeHRgytVdCBlMNnG0P82tdjRNY4NF9
+rB4aMZYU7JKvU0ZY3eYylyHyoAtK6UZtqfmCXutr57eovJGzzQEv+mRDcH+jMLk
nsqgksvzR8QwCPi0aStaNds+IpT6DoH/7arsuAuoIcV2A36gfr0nVB9Q+ImTrjJN
jC55uNiuFhIHTDnA2VSc893/Oj8sNNPgmVCIPZ9PboxccRB6kkfkvSligzmlGSFs
ZGwWFqDEqxzHXsm2Cpiuuc2DMz+yix2/zzjqkOZO3XNDHLXyDa5t7MiK/540jZS9
k5BfU8I6puOJQO+LVpKyRAVdZfr72PU7PPhri3x6oVv8k19NbFEqiagfnV2JyKXF
8evH65b1ohqCxTfLZ5U/YW0hLo5AIt1WS/b9u3WS1T/ZLPO4+VYEXPyPMXBmewdP
hVnHi1aWmvropJwhTDOg5qZY/xT6IEJcN73a/R1kywdvYYmP54pUYJmOdOmhd03G
EnDc/NsxYLjgvTyY4Njm5Evx1sWjX4nyPwCETyAfoDBtOaH7IRisc0bFe58r+BsL
ULpDZcbzF5iRIRt827BErwkQrAKW7DG40cgOjAEs4RllzVFNNU4kJwR4sN9DP0vL
00BqOqzqiyt1ZHE9zE+PVEp7WzXArIvR57f+BRFnRwx61XD5FuD6JGw+uiqMDG+S
Dx1Qa/J/m10R6/zmrBpBtFHgj2ZdjfruetPZuTYHCjDvAoeiSedEkueKlanyAIBq
LV5o81MYooXcRFTDaCDkB2OEDlr47SsEntrUQ65PDlZWlGytwrTJxXqK9LwXSXxW
36ZSbmylTcTqUQuWwdSSSwSPrtuHY5lfOvc614A1UJIpwfUbOH++43rwVmhQdnzD
XoNnhp5ASG7lVqcSlc9AlK9wQhTIhsMRfZH1c7NlbatYaMEv7bxUe29VT92LiOxh
2+ul4RfH2NN2hr+d+Ao2LZQb9pmqsP/XfNFvrGQzQKtID0He9YN27bblDg686hD/
0xJ+DPlrqySD4hMnHOgC/cZwT565EiAkxefcKvv0JpUOyxP17CFgthUg4NOznK5D
sZ1wsyjQmn5CaQzw6i787vBG053lrqAE810mc+P5eyR00vLtDW9Kk1fIfEoykAzl
Oav2jcFJFOFwaS1I1UZsyyaDs/rpgZD/DNDadmm253RTzVbyhw66Fyhr+qPvlvEQ
p2Fykgpwcu7mJyMO6E7ogbds3SUWC3pDJTwBV73lDoeBAkSZGRwO3kPJBSo9epqx
QlhSmkubjr/biPpojEOTgidl3yS4YS7TpTXplbyFHFFL/AhhY8uk3KEYQQYer1fj
FNuSP4akfuyH7T4wysQcsxDhvji0PaDIBAwrAWDIqhMkrm754Tk18nS143QrGeDu
Pqr+Q9imCFdDKtqixM6uh5RAZO3SwCR2kquaJVIiSKOzY8oVExaalV88CT+AACKy
Fome2hx+0IXTD88WZxnHsaCKT22IhA9yhIjDNtsiaUnyiX0NZRxepizFZY0mvU6s
uf5YRKt25xQyWS0T5hob8BTb+zEDpUAMQSQuDY836AlpUkd3cmWkrZX+hdYE+GpQ
fsFKkHIcXhI0kjuBnkHHbkw82YUO9DTrK5WlDYHiTO4oTZ8G83/ZYLkPtrId0kv/
vX4BTLbvI8ikt+0nylCuh7OhBY3aBnquccAuNFUrnPuvdHMJwBxVydq8eAxM4Oro
mZEVz+crEKYimAAavub31Lc/JZ/2FCaHJ00Uwf1ZhxoZ9h8RN23b5B06kOLMtzkg
DzKXOPNlSxVzp/DHvoH9PixyX4BtiLPkG+K17QJaKE3vpnbMZ1a79pVubLswYJgM
GaKvKbLtOe2Rkk78g91l3goYFyBvJiGio8MjUKsmyj+qisI4twXqPK4KxrueW6YK
ZWhuj7Z3jaNXTIfXlCdBkx4Y+TaWSvP3FSKree3OfVJyQ5IzFCrvycabXKqU5ysJ
w86MRBr1kDNnfT69yBR9En8i4CWhqx2TWGDuHZ6OlWGwYuaI2gFOtOWwT6ZDOzKi
NFxDpUuO/ZkRokK975TXdHElQI381I2ASbofO535NjaFCf8+Zj+TrpnmxyukhCkc
tuzYaC+IDdykq5T3kU4anViYNBOjj0oyt/ltx1cLL0f7rIZ6Lvjxcn3Fr9tnmdFC
kYsxpSjR4FlMHO9zaeFRTQrf9Hel+sPDfqdLrM6UNmPqbUbE4KEgP6wgFev0LOUS
WZnokXJiF1uVxemFm1hmHMzZVuCtomzhPLh0F1zjLkyCqhJLW+dHJpqpS568kRV7
klCjrB0WCS56hT+hHAlKsQ879VtFubeLeJxUOwaEToK0UWfT/ONRS8qmwYRVU2ax
OV2tQXiai1R3pWYGoF9OqzlPrHxBWAhWM9YT6UpNqqZyX0U0eyZqCfzlAzkYbjWs
/ygX3mSGeZaFflJapfnKPUPMkhxUYmbxLhI1jnUnZt2RgEzcEp/1BjJpClxBCppW
RUxzGJkxorJsiuRCVJmi5x9m/oRYb0Z8CZXlsaxdDncJTRJVU6fRnDZXldBt/1Hm
desfl5g0sImJz0AgI1oKdPzR3Ps5r5n0uhWvAf34olddcfohLe8u9ro9Hzo92VII
QXeLL0XD0vWeirxrBw54qnMon8hgJ4Tx1PIglFRw6/VaB2jC6Eu4V8qnX+83GLes
PWCMkAFlC6dcFYc7ogzgeQoqhPCeVPhbNS6hhaSVgoN7+RMlM1YvPA081sLOWXsb
McYAoe6Zmoocs1QVA4ZxnJWjjnpPGA77M6rmqChdzuDahOdUHT7OH6tgEBkEWbgC
XoedQuR10f4cp0D33nOiysBBtZcXK8rjSSgUGeeZAmthVNYBPZ7hzekXrDMyc8fi
OTrGFvAof8n9i3ofnqMyixVgw5NeltI1dIjyYRUNkxCTKqUT62idBtdg6yoZY8cr
GuGTfTkLOszTRQNmN30Llim/hxyLtpmRCJRqlxY06HzC9o1ih4eIw476kbozHjhr
7wC4WT2I/zRDU5et6EYL6jLeP42ZoPXfQyM6DnXfx8HV4TfuHmF0FZbnjpFJK4e5
Sx2+UL1N58bjSM7H7VbIIjcz+qON2uwGestlqXBWTdZTrJq9R1vMbp/S9lbIfO82
P7hkKmGkPcgisrsNbcbVr6+PWTPl8j0nZd2K1gbUbaDycGPXBXRA0nfzS8uaNDJT
HOG39Jt4X3qikScmYhxw4TrDIqEn55RjUDzwsw7SJBSbLnbN4h+6NC3FfhGWBOxf
2N0P9KMe/jWM6UpxoTC/A9ptLc5yOD/xhcg6v+YVzJd5seI50ldxhfkrHX4SDYMr
bCWuKCFXzRR2cZYd2BoJeMn6ejngCJ2I47XIYIpUcxxyCFQJdu8x1Ovm+LUr7i3M
Ua3+zxe4MUlZFj2RGLtJ0bSnVdqmsUJOExkXRnSulw9Qn52RqBrYxQFfLlfUkxpk
BkgAkibsz7ivMnZpH3KTK5LV1xAYkvctSMua4Tl4FKIM7tlOmvyZLr5m1Lx0xKJy
iss9xRYO5mjoHnhSnR2p+W1zAyECpW78BQ4D0gv+OIIVgfIH00oBm/6aoDswk0H1
DYwcQ4Vuxe+b9k6IeK4tcpOUj6se0Gid5puHHGBCxpl4BuMbSHD44ihGPTfY0sHJ
2cJk6GXLdZSe2r8rMVOgoIh1XjFzWae77UaU8iOXSoHmPYb93w/u37L82E/A/7YS
CPE2b7/Xs5swOvhQpP1C49DnpvMprNPWxqGmWAoLRm3WLTKtby2tHLY5g8f3Bgw6
4ECq7SU4JjjF33heOmZoP4O3++k2dobnV3GOyp8DvS1abQtAmYc9Ll8lhViJ4/xF
ayBbLtlqn9Q6CZkHyMLhrWBLRUgrwIN8QI6haWv8t4uUj8RkW9a1WOzz7XT1bf4C
BWgza9GuvHDlxbH14zicDfXEsBZ/ZRraeax8eUTpd3QVTCNMEOXoZBa6UhsKsRY0
KVaS1p/FbvqnKMLUl8A+ukknwRs7svg5dvOcsLXdQd/7hQ13UKRLFjr6azUvdh4+
4Rb/BpvDm3gGe888/Qwfn5yQSzhz0WzqcgzDxbVB+05cr/XYBtrxbhjLLRI4Djmc
fOBriO2Vg0BB7PePFLjRbM4MSNFa14mAPzXru7V7XNGb5CitPEOhTLkwPsi39dus
j8H+06iMzWp4NcY6UL2UK3xHHndWxwHWcajqwIWSlYQZ2OZjDu8/JhcWHY6rB5Z+
0ayrbPhsWhX9AVz/FbtrryZUi6SK5li85XkeSQFuaCkFffD0ha5Sl4XnACBKisi8
N51Xl2l33S2wME/oZ2r3VDKWZHO5TAxSHXsYTqGNO6im3g7lX6xOSGB3YQ2SZRZk
36MoYxEeC7UJ21GLTaIPyb2Qny5VmLKatBQ+IfQ2kF4w9Y2d381P+aHhOL7JqXB6
Dbc5dHrDmDC1fLApp8R90E1ypTnBp8ur6oi2x2ZitBAEUIaRPf8SnRSbNKXRTOcq
nzPCNtWKF44feRaQWy7On6rNBvxbOo1aLeosGavIAp+KXVO3bH4GyawY5Sqo/9iJ
5XYEulHu7lwJ6SFr/knlXKYzFVW1L09/+11bvyOobmEjvYl6RX3OjHFVaZlcbC6Y
7uPfRGvcWmVrhb/uLu/C8G356QxEVD/8HmsV2BNR2q0RDUZhgk3kjJ6k8golXCLX
UETzzaw+usumOphnw00Tqi5ltz9ow62s0ZGBo92b1BbnkFOQhO4YAjOKpDZtCpUu
BljB2qvJizrSMAu+XQqUlO6FjjMZVWYwrip6TUJ684trnLEFoXfJ/e86L4zfa7nv
Szm54N3fbU7tWTX7/Aa+pWAJ7dooXVqevs3PahGzMBzxoegKh+mctzdj9BAcn4kd
p9Hpa1zAQWeTa0b90vwq7tQhM9sx1WjgL0+nJACw5F22vNBnIGWj29kGhISFlkB1
rgtR2llBY2XhIeF3D9S5zQ69nIbchJV/9OmcQT/H3vGKv6dZbEDGSIZWtN8eMsnz
4svgwmy6bWSuAOvVrNLqGfzQiDSjanJjxS5LrRg+1LcsOq4E8TctyGjoGWmM79dp
9Qpz1KzKL8qaInJbOoGw4+t7y9nmEuw6O93iDF7KaSlxAsc5ighSV1v75DqG4yM7
aaDXuiqxt03LB6Pf6BbbbFYosziaBp5vhYEeSog/RaYk0aZCAv+nRIAqbDZDUav0
nhI+D9LyqxdE2yJV5kmjTPgytDqRandggXI3GAua3S0TjCvGk3cys5LA0sXZIuwc
f2vZIkmqmL9JHSmQk4yNKgnyyI2Is1QICiVT4+L8RMEqZwz6nTeKgjafPEROZLOj
rw0KvL4OnBh5X2wrstzM4S8Z+gkKZBsYH4I5a8CR1wJmp8iz9aHnyzXkUEG+VnIR
e3b//AV1bP3uZrdcoyS+a8l3zRTTBj+Mq8Te02AshekfDeAjvPX1IB+w8+HkiV49
/8M2rt+fAFgW7KuUmsKfjT9qCW2NyCme3vodZAnU/cCuWUgUkozq5S/8C+/98BsG
k8MIspmQYcEZ067LmLBdVgJfbOHaDasmbPpgO7ksTMvic2TP6ZKnVVnfcHS/XyXP
ZlAh8MQL+sNdLxTHXFV2/L4qon7GDHmf4cjJTzthoz/ceoFFm/IbOhpTJifjtLge
JhN6+t05c+ZTYpjVUOtfzlNCJMNMU/Ag+SBkkGWBTR+zThXHDCzwkBo9naEZX2iN
BXLPyILJKV75SGVLMf3rxgilMK7kgLKg7jw+JOShXuqBL28gi+LoxyY9wYkmvdBZ
ZiEW/GOwO1MXTQP+YwGD4t4iaTk4FotKogCe8iwnhFqWJKbQKABWDHAEITw2JsuP
IA+PDRFbd/oSHDohhNj9CRkvVmAiIWj9e/ndNJsQ9Oyw6+0Yxl9CbGsqbjpiK1vx
2XF6lks8WNHV+RYyx22m+mbNMPnHrInB16lnVCoXI8pXoY5/HJYcsYv1SpBt2lKY
3gTXWNv+EABmwbrDSLYr7fPcMtTeqA6Ca+Pmffzw+lK0RKRz5HYDbQx2HBaOdpwn
GYkHcwUxZHeEClKSXL06I69hfZV3IfC9e+7YzN/qDZJ9Iqn6dvoGMkGUI2sYMKf0
wB+gi3y3eRjL6elURuKw4eupdBtxE+m83D5mJQnfzR+w5NhGdUNr9zvNx0iHYWW/
+UIy9rkEBbbCOR+4Ipxop61M9Lc/9+Cn6AkzZu/N823sAqUhEHuOsaPTCo7sb2ZD
KVW00w5/w/qZVVPC1Igy1RmeS0P/vkOpF4/q38P+116Tc7HrZtByDrubU4g0xfOT
ZEAxV2fgh4uNe8xFEzzSMBsFghA73MNpDcRGe6K+w0fnu0VPbqEGJ5fQd7wESTzR
x2S/yAVOjIgnJOImoDDGud9hjCmHjObtd3rEYr6fGUtbXCuowKKb1FKdi4IO0eQS
T7GkFTXmc7ys6u7/AKDXxIJioLTqf2YBwpIjpnMhpZ33HgQnE3cgLjBUsA3eWWGw
Ek4tMypJa3SxE43no4MXz2cLZV+OThArzmiVAM3UPkbBQHQiAKbLWOt9d9Wc2oSF
OyPpFumEg84JNstJl2fT57C4ENFXAipipxw8p9YY7uUM7v8k2OxfyMso7XRgDVN3
yT57JKy5QPvxIjvhqJA/rfT/QSYo7L8wMhyrzgri7z8XHKjOMTTIRGwWlt4ytOkc
VpCCWjYQ2raeEutmNIu3V+uRM4UZ3XUxU34jvX7cT5nPe5sNDRTcyvhWsQu6Hbmn
9Y1MGCPOQmPZYT9FWGCVxAiSQqV0BYxEEHzULBZdG0yEYrqP85zQIR3Z+eazwfAf
UUnN5Qn/+ABKvRM1WqT9YM+gH6VNyXwKgbOQ2x4wg0p+LWTcCviqAbvUuaIbOFi/
t+mQnLB63TU7O5kWQtIGes5WXRZ6YWwxlsHCndR1Fq86jSyOft/T3BhNm5CXGbSJ
BKmAvDL1eO+nipeoUCTwwWBYHUVs/M+Q3qhGliWM8P3rQA8FyzSfM7rkSN3HQ4at
ZBDX0m6006NLFbVNXbrdOITpXKDA4tMYV1C+vEaYB9tcko7AEReRdSgnBNwT5KxG
iKloEfGG08CAfN2yzJovBnoHFntYBirvEzcgW5oTx8aiT+uJ3oQtSJ0PfWbADnDK
YQQ8uCNeBlYbV1jNLFrk+0gadASK9lHCQDnBenKPKgDrLAergRkXlQA/7vqHRm8A
bqjSMYpwg94MFlgiwNbNHno3g4lJPznPbGhFeP7KAT//DpG7ZZ0P3OU6pdvLZd4C
stenAhYjj8SQ5Bl1nK0p/BYheoznV6CYRJPPqol8FSQxLZjjBhA4PVcOFKlIBW8D
clDAkZ+oGhHih02tg4Rm64uXb5/RPP0SHNXrItpWMHK6giVaUJTcgUtJ/MT4RgKD
q7DPesvWe5+bHe8OA6vsmuoKOY6xXG5Xr2jmLAPD618JIu59E4W0qPPzjmqlQenO
et6+BXi9kY5Ooq5A27tMIUxRZSoTRK0VSMKQqmPs4zhy0MuA+bxBVrR3DmPx/KC9
4fXrjYH0Lhm6GU42qL2imHoyo//LSg9xGMgv1VmusFimUxjt8cP04QCJPbR0F6Kt
eg2O51omWNLbDNSoLaT2VDcDgeKpRvq9DmxWWnjcBApOxYeTryMx7455WIXZkxjY
TrH0XO21ErfcIIu8kmuwmOM5YBPxoENij8qh41yOZCrXHVR4agSe8eD3jSEI4o1i
Oy62fWfh0ayArqwO1uR6UHmZS1jGv8vGgNqIJDe3K6bJ980iPt20fg/Nb2C99YEX
i2UkaBDrcOQABRrkcKy673omq7my950A6YXQoXdDnO4oA9kIyFIn3CU04Mxhoxii
qTy51pIj4/KpFiBCefJkLU7Y/b1Kf2DLyopQvU+E9aPLIhYGIF7UP9cJB5Yoxn3V
ASU/bYp+MlgN0lywyZ7NASclvs19IBLDLEiviu0z5aQE0UDjvVY60PoanaCIRUj4
Fr/haQ15zlkD/nSnwS+GUtHfnBSfihC6/6mb3XYhowWfiNO7a2ulIJNElt+z0NK7
X4ykh7rMPpmKSPf0QXdc4vgIWsLlkQt68uC8+5Zl4EnOXcLtipH8Wol6kOSZEQhc
IORw37vdLJ3SAVg08lTnwgCTaVBzofnLk47g7gBQaueeZ8LdEQFYidg2KtUwLGHd
pRFlhj46JtEJ2Wrl5Th5bVNZ5+rZ+9I1iAfGC/zkfUI9gNELxzUN0Y1t/WpBUe/Y
SwZaIA9desNTQ13HQcxiac+oJUakgSmQq4xOP+/krRe55uLQj45XczXKSY025Cxs
L3eYlcpa3ykSgiF3PfFqVmNgFoFFp4N+iloVedTgp2x5QpSSkW64kzMnQUPAJVug
HDOgjxIBOLOiik6AITvGqFMt+1fN9gLLQxzuNLudq9xsVAV6nIfc6Ktv6HVad9rz
mI6bW88KiWY00s+BgrxS32TQcZyId8w7qOz2rbHTgwgBAQbN3+iGF9NJyYZNFujE
ve09QWSWG1nYpA1n3PeMfoXLuboh/aMfTcinlSR58Jqj6iDzBoXwtSwoFpHiosDi
0UKqvDU5pTITlPZR9YSpV68gAmDTAlggdneXsooT0IORrOIjCkIGeswGa3bECfQQ
aZBDgYGllthCyTn9saHGkaSDTKhQppD3aAmczK4TkQd9TcHlMcFwPs/WDV1h/7Gh
XhmW4bMdmMIvLAnceus2m9XSiz/V0q68+2WmGVlRaVVJkMcmFKQI2QGkFA27YNQi
Pd74DVJ1atP+2BRfL8pdvaPjuezY2q+s9YjbVdgXeKUSX3H0BYFP7wo6P21Lg3gh
6E6n243yaBQTXWXMbA0tSBP/Smgof2Dils99Yy5wlARAXywDsKSF5If/LObmz0Pz
sXnYpDoNHg6swlBjVgMru/O7llG8FlobPYSvS2aGPQQYRNyBfMzK0bjFbvrz2FBw
ibGgTr6S2yt381h7gFnkwEQzuwAqFpKhPLKP8nI/dpXRLQ7gkUvqnqxSIMIgI7dO
Pnlk/0ZU7vGFCi1qJqULsi4EuIHSTDOvRgwJz1U3rQjNmi40pNCRVUKau83P5X4m
6coo3JFOavFCpamht5J0CKJcD4AKm0ZCaQf9zRFUAIUE6GwRx0Gn5M9jmlyrADjT
4CAedFc5iphD1ePS8ycqAHDeNpOjy6ygkuatpE3RDdhzHfr4h0Rl0cE0jC8B0PwZ
G4Vf0B32GZ0fJEPg64ZjyD/e0SxuX2XZEcCsY3SRWbBfGfYhQUtwBh+mH0DC4PvT
2BIabqE6IchH4cd4suCDIgKPuyJouyhg6xyivomODn/XXW7nY+v6IvPMLHrQZiYN
8WVVNMj9IqQ8AYXqd1D+wxUNgJSi3WZxhxuaFMkvccPJfBVPQn5aT8nx9YP/afsW
7RkDN+bcoxGybOGKHMettiSCBcg51mFf5Jkp4LmgbSGBbiqQhgjjjBzXiwkUvRlN
N/J11SuDQxfyhLeMvgvzJp9jgs3lLS0r/Ej0DUoPBUoaokOghQcYz6IJI003XqPC
IU4L7eOo6HC00UUV1ySw4ou59fbE3OcguA/Pj6kqq76Y453C8HkMB4+TS12iFAsI
Exs6CFCeWMDd2HgsPVylU666DqZykJ88Dt7rNRVqN9IqsiS7cxoo9U564cz5HGBR
MxYzTFSRcqLOEUtuiHbW7komXk2TAIU8ngxvsMSYXFEEjqbbgVUOBMDiudd55a/s
fj7h7UDy+Idyi2qZZr7YV4fO/dMi0DcHeH/UxOxQU1HIB4twlB/K5TyuWHQDtOUx
K3kZZCxTC9Po+Yd886PSxCsAxhq9W0da90d/rCOPvyHQByEKsvX3JQWTYPvST2/K
ug9dINFOl3z7SqzBWR6/+GgaWQO5RqCujPa2v8x4V4MERs372HBVZq/BxdizWhkg
t7nW8cCe+hgBS8qxEXdqPRoiccgIgqCWF7y2+vLNqRosq386WeKfTbHBnBG1tHci
euhjt4il8RBld80Z06LQrh881Nl4C8/NEtsHAMeATSIpSpjIWfEOgXbqs1waANlh
K4bz3ocLziIHApi24XNEYt6f/qvV44a+Q9H+aC7gRrW7gBBIIk0ceOwkXKQ3PxEv
Rv6yyiTsHvgVYcanv9zBtBOdMMj1K8atoIS4VhHXAeDAsDWNrs+G4DBzu+ZRM9zN
CDP5xFYSi+ZyM0kvyoms5mTWNu7IW4mCRq+B3N8cI21moRo8DfA3/7WXVEu2+70B
xmDGKRTiDPuBGwCxFHKXAN+/Lv+jv3TO+LF+ie9gTeaCLxgi23bOjyUFVD5BDI9Y
JSXfv/JgQJ4TFzZmbHZErHC/2TP6t+9Ap1nOrk1v0BxDXePFTWRhhz+FqODw8avs
JYWrNRq1zwFNwW+CHmDHtpno0djiBaz2y4j877LL5HHEBOGLGLvtxi/QLVN0+7fM
Ths8oLL5CwCKu7+lrS8KWpfuRD1j5Yhpdx8wkRH6EuRo0Im+iSDFHA3CAR/Y459m
oTQHPQvi1KaRwY6jzGBb2filvxSEVf5mkGMMymZt9P41jpy8vk5OYowfZPkl780a
Cciy4OZBCp4K71Yz1OnN/r2dEhzL/NB9Vjet82hBL1hVDwpHCoCbfTnggfYt5mcN
SQkEiEy3QumQzyml4v1EaPFFpDSvO7bDRH2W/YUUY1KY9OKyQ13QUA33UyVGCDGx
yrP5x2w5MMjT2STVrjgU+1HISTqjP6c9cYSINxfiXVFIoV+2QI4h5TLDFwcEl759
g6OBAIToK615bfoFNg9WloULfjummPvFcJORyg4ntSlkTlDBWolFtQSeJIcapCB2
nJHBq+72vvqXh8Lj3mWkSfy0GFKn/aE0pAYuphSy8AsNWXaZiyLVI50JaM4e7RQx
GNwvY2UoL/vl4/IT690pmmdD6ldWkyZHtorPI4WBh+s1bT/U02w4dkHORWLQ6+RI
bX9JZQTVcF+JEXJ7dymR819iE7M65j4RTWoc03EqiH4A8+pCsxEF7RLB7MR0YY6y
uxV+QxLaa/ZSEtlt0Fstl4XxO/qV5pFAthHptBkWdHFVpz5tmq5/6K/Z/388Hjxu
iRMDvamI35hp9YHDHGKZtCLTM7IbVdI+YOzHt2CjMI7lwZn5Oh1osKUn28TJPC+k
1vCMWsJdzpKaKPncreg7FHN9DpeBPdMTllMjiOsnuC7E2rLq/JY/1DDiZzDr5sKp
C9LpeM75N7SF/ypzPzQoFKAFNpO1S8P6zqV0WSWVBziPCU8sCkr1Mmr9wePLNq/P
Q0hqR1gPQWNdZhQvmTIQ/r/2v5ezZi+43R/L8VfBGl+/JJlZL/B3BOMSk53aqFi8
9EQJxwZ7iH4aIMqnWjZ0QOm1ZSb+FT95VdqGE36005wCEIflJVo3ifKjMWEO/9bf
nD4zEeJLxwnZwVEYaKHBMiwZfaWaFFAOVVsBakCdmluhSxC5LY8u62oSAv84gYMv
Dsfol3eF10dCEvfMqhNsg3vOGRI6QnFxEE+fYIxn/bPumO+jyBccPdVurc4v4qzr
YL8rMXroH4HdfNY6XiZ2KdWTHDnXQpLjdkWe8SIkx3cW5rN2vCJTkxDyU/RH0rfq
bj16Q4bMeqiIMhGLtSbC1dow42chAKPKfEDzyrvKn3X1cEoCnIs+cNumxzO1AyV0
27xCVoRlOMjBwF6CSoa83Iy8RemBmLzJuDlRxdxCLdwL+TduwhfJzEYNANfarjxW
tVv6p7rdrgD4m83QxMTEG2d176sXzdINfd9YbAyI6CNe9wBQoD4lujAYc1DqiQBL
0s8KXvaCBv499r983qaGVmmzZpBv+FGZwi1YGmvIsCX8b1bBH46lLgkgd575myjm
MMd/I1B+cERngq01rcOGPXyqLt+2yPsq2googWgVcoywUO7fstYpT8f6PmSFlmpU
DrHuYKNnwlOuaRhxj0xd/J0CxMkqLp/wGa/K5P1uZknCTqwa/s1sJvbp0xD3Sniy
0dOQc45flelwAeqyt29e3MUD0gBd4Gwlw6wdGC7Hw6YcQpqMoeRHVCuKX8S14SJp
M1+d6GJYgnOcIf6jj8kgG4M673w9wa/hsEtvGIttBaPsL3Sw64Y05vs4Zu4afAAh
RUzqbRP1SSa7RlwP/1sGAu+FOUZU8w2Pny25LuCR+fHSd7eb9VVXlzE2XTesaNuj
CSINVGk3XKv+aJK91sa6FRTgMU/dnYsN4OJaHBx9mRRGtT9ygRMRIV6kWoSDgClX
oOnSHMQw8M9wTx6o4IhCD4pNG3wSMNlvZBx55r8+s+FQMoKmv6fCZoNE+0Ty7Oga
8E6h2wEG+A1q3ScyG1BtVS9f+hEXj0GMZuxVO0aTDQ8DPQyAbgWKR/X0OuzhEVff
SX9bXYAVbgPjrLtVSt12znsouseNK97sGb5i4mc1OeYw9EgxlLqDVkEj32vMZSvX
0Wdrym87DVJYDU5BPWra0Omo6dfcl9fZF4VCNA2lHyiCLUZl0fN2C9KClk1twj94
FJkQNs49H/yyVK8VujuufMNAlizJnG2H41+YSQgBilWDWI42C22cXw7U1Aq/dCRC
1lVc14+xebTUujcUnR24J3CunBVZdP5f9O4Ba8RbRXVPLaNNNFNykcjKWP0Iemh2
mD7yVbo4fkmG3l4u+pTtHfm+02sxdlvwUK9lAkstu32N3VMjHjWKx4Rvrvh8ys+4
UYeSl/6BW61RGnJtCalYsCWojJu1OT+H/m2aWHlXa5Im3EeZ95xwDEqSfeW+0hEN
FHY5Vr5+Vsbp7tg+nH8TiaskgYiUjV8w9IqsGmDeeSbZeo1E2y9yGlnt5kQkfwtG
0NxsQDNPtkHpIaw88jqr/JcJ52K3YnhyXHLB4Vdb5SztoGwz39PzYdpm7TYqDUMr
dfX73tobR3uliH66XTeWtgwcLTdHoXLHP128v8wrfu4AsarA/CYmYS+LxK00zTNK
tzgVk2Odc5gJMXTC8uuxm5cYG3dq9SWjKOGNCxOxxivTXmmyCYT4o6c8EgmQxyXY
szznS1l5+wc1b6hR3JJfzMld6VqlUSL0SzGAEsWD+7d71bOWoVQi3Nu1XwGjPJjY
w9aTUFEwgKEDo+qYvm/+KxJvYUzrFxXWFIFqHSShg5he42HDn5Tk22zroA/uK2vi
/SeYmw9tCwPLNyrtrr42lNehcJicbkgCubf1cI3QDqVDuIpiXaijclHZcqbBRLAY
j+BL7ICdRBws6V9rZ6PbgzR53BGyb3rJi0CZsvMKj7gO7HHIyTi+E5Io8w87MfoW
N05TAZeQb/66dlQomwZP4pTdVHVoXqTlpmv1GTX7I/wTX9QoqkIvoCmbaLA0yR/D
N0n51EBSCycJtpYJrFIFgYS5D546d/fR25FFTm8mRoxQ2OeQN3F5v5kzk0+LO5nO
wlRUqIWXxdZuF45smRC+y76Iq5rhPOcSkYg13Bho5cWiIY9svar9Pv+hAsVMPFN4
kcO4kt/t1gP+t6kVL7DdUadGKK8MAsVic66yQrvUriRyx/DL73esOAb92xmrNGRX
U+27vBQDY01+z4LG8RGxeFfpmqxQHhh8NGLg2MPgigzGky28q6bqxr01NW/8y1Gh
U+Z/ertXLF44gTGBN7rAM2Wze1QeRAtTlDJ6YbrYOtpb2GL+0e+as3RspmUVgHAA
ELm3XxILs7xLtoC3GToq+NAqXhRn2bSPcvsMIsZ4M6iinMZzvcteQD+ron0jeQV2
CNRXDC+MtNCgXO608Sy9Jm2geuNzWzXXvBwBmU+exApaY3T3jE2RTR1rycea80FL
bij2rgBS7hOyT8pj1Rufdou8BwRjvV6NhIHiH0sQwyeuOeBegZHv4FFKmzGKReZx
jSyhl80Bf+fTRCRci1YOFDLfdo9SKObxZ1ZnE5dqUJluiNhoyOTKHkoZ8L+ONqGn
m5ZKb5RFpDEAoY1xnwOb6pK3/6rcujKB4zDYwFuVaXe/ThTs7iSLs9V6jqnfTKIr
aidZZZRi70lXwNu3Or7bUhlg2VYFhSfKs/NccAqFpEwm8jsMQO618npT5+wxkw55
Jlu7s3CKlNjJmC/mkONll5S9VqraYlC1r881H03J4zM=
`pragma protect end_protected
