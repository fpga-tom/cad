// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bLgAvBjkg8bJUpaXxkeiMtqKz7MHP0SFaUmBfK9EWnWzHlNQqXEq/nzxT7tJRDbW
8UwAczWuy8NKWMFyiaubbti2mBxdhrAU9CZHcqUS0EyFTdJtH0na9JFM1/Bu1+5t
b8xWWK33xJKM0NVkR5Dp3/d1OIOGL+8nUoHX4XuSIEI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33712)
/n9gAxP7UCIBBD4OlZIyboTy6o/PLzSZQdX/pfHXtIap69TzxFwa8mmGsQZlwMvP
23THgJd2lc1VCRiPsM9FHN4UHcwouLBvQ+UJm8dpmygNdJS55GRCwyJP7letJzO6
YYBZ1ZoD8cxJQ7Eos+/MqKtSodkU4euatvBALff0mtC3Ly6eKvlnZUe7cFKkUG4N
odT3BFXscnL+XQWp+wCpmBYtEUzYaQ0o0jKeaFrzschonYcnkRX/2jvBe6LJlDyS
K91SnHji6JgMrLdnky3Osk6UQOkj5BLY3LtUyb5SU2tOyfB+r1dMSaiyxek3yktQ
SnBRqq6NIGxSQ7mrZoKTiXIET46TDmyq9gUNx2vr1MHk3iLHz0Z3DKd6lGNmOTmz
Y+tL3aeIt2sjqEoGRKMc3rxibqCP5Ff0b7tNJ0b0aKsNTYcnMJm2OeRU1yJd492Q
DUBDeyvlIpupYT7XAm2EWzMH4xc/O79/114Rf5D9DnvF0hoszFdjuK3SGN+em0qi
sBUT/MmUdnnUAet0v0Aftv0WfEf33YfFzBr7m+uFnSNWasKPE7ggLpqu50hB7vIJ
hCkCtLht6SJju2Ej65RZNvpEAQn5LuETRhWUDxQZ06LOH4t2N8u+GnkehF3P0OfY
A06jLB14gJ+Lx6NLWBuYrAMiZidM4wGZ2VhKsXXKF8eFI9hcY64jrqzVl5fSQP1k
9hE6c2ZlaOllxXEX+hXUwTLcOEuE3g3prY/JyIyMz6V/9/a/6ptqv06+cGtgvFbX
6VrQczio+0k3x0ZSGiKzXp92URJRSeikBsNSj7wlDcUuN/cy+1aadZqzqXvRpOd0
4anO1tEnlvIS9PrgaZGC9b3HU3VMrKDKnoWkAAVZUPUaznmK+hvRSak1nX93ztH2
uMxsrw6KJz7QplA2TYVjRct2QY+Ktoi2LgNdiZq50lbwdSsOEF1EmwtS7gx8/Kim
UO+bBBIGrpUN1B9nk1IPcZyexxhDrnO3RUxQKouZQflH/RKwSHE26SNbqID07u1f
q/Ze0NAGh3G3LbR/zz+CWg9yWLuHgnrV608MCvCZf5SP4pZG4YwzUTYSU8a1FMSU
pwjB1UOBowbLo3xKNRI3l4GPGiMliCEJvdvlBzdzMD9kYNtp4f8jV1zk0Gz5aQJb
zY9aBdsmxcLLTBpOCa05caHmHsJJlH4lM6d7piS8L35FJa1jOsnIl19cImhAvXVA
2YoBgDChwh5DZ70sfTrOYE3+KeoXWkPjJaYI7WSoUxIukNgS+8kEzb2Fa14YVA3J
KoAtMzh5PGCNa+AZyYLSGWjHfgtyu1D6gttMusYXITvjQkuqkC3Tw4zuWN3J/4WZ
9IOIkapX9IqrUGE9Duj6m3h23MobkL231AVGXPCCow8tgJTx3UHl4t5G0aBy+o0t
9wE6B5tzQfT2E7DcsNk8+AXMLBXgXV1AyZGppcqCEyJmg3+alM6DNbCWz9NrmUj2
j7s+L1IMQ+r0gvZhrqbQHyEMWFLOGmPSNUXi6+bfwyuBIoeEC2mU3LPB2x3yximD
CP0O9LajUr6JmHq5Q7oaJg08ufMO4qTX8eSNRV+kQsjQE+fYKF/WOpztuftU7mO0
tsdUMiCyr8a5f6habwBRDbfKKrWeaaaPfGIqv1+dGtv9phQBmJ1FGWZpsjan2nuI
6LJctkTQdmJONLJ+bQmwKhTbFY0dku4eGkG5Oya3itjkKzOd3es5Oey3qJc4lysP
NS0nOqzJ1lbzAoB4erObYrYndhz+1CLNxN/kuICbfBQf13v5bI0hjIc1s0AK8arg
nmSJizTb9Tdj+JrVgnPUMgsKRSg0KHb7babJFy0RdgLSDIwWEn/1Qrl1AGL1K56S
IjV3ksL00oz3K+crAqB8phhnbd/5sN9qjVBQqNioODe90uaujNJn6JogxJgHG0DH
WJ4RY5QqJUshYBg7zJGnP/p5+Zb1C4U+lKq+rAGRkqc1veupZtXGQ3GCSCNc4NCw
6esrl3tvJ0DrH4mwTi80FkrDtJByYqg+J9Angqgy5mKT1+LMUkN2PRa9+Wkcf3hd
KutXNeiW2b9L+jE4/Zv7ZrkVnxH4miDgC2EJoNdOjcfbMD3jLnjaiTcLBEUzl6y0
85fvSHUwIUhxDhaAKwa84Z+GA5bIMxle6QFyUBy0EPTpgMGJyZR03qKCL1w87jcu
FV0nKBOGwXUrst4xnKuo9UkranEAFO2SpkC/ISEyCSQ5P6053TARrcP4diE871vL
4I+d2nNEC+mg/SPKsn2dSyQVBncOFdahjnoAtONIK4AVn7cwnnYd3fIBPX86GhEK
RHI0oo4xrqo35aRF0LIRpNqDhNgkuUy470tFPvD1lIqqL/QcSZbeatrKbgph+Yqw
XskCL8d9ylE/JiX+QlKybbOhO0ndAKs7XVbnJ7mLc7+PpeHdss+hrCbAjMuTTHUU
AgZUgF+ZxEfloks5+p75lMYajKLsAlzDCsvES/zyI6UeQpuLFt6NBsHB0UUbhO7t
kl9p7IhV4DwyO1TIorPCX8cwtvCYIe67xsV24quOCYqmYYO1Udp021QJSOY92lCO
FU6gBSZt2JU954XdMu3H/KrDJgPUL168d4dIJYGoYrUPjjoj4nvZMLRvLHfpY0xs
MVPjyxPLnjZ4DfPiwmuu0X3S/S2K27bKxmZrWHHyER1qy46DmYGKCW7SzvWkP3Qj
mgfSzYp7n9KlvnkzMC7y8L8d0F3taY0DM7Bvo0XXurqWPgnjhQD3s7sU9WVNrRHC
7vir3uEYhmlJS4wBQTymi/8iVA3fqHI3XQii9KzVZdpQStISZk2HC1GNCYJUhlii
2Qg9dslJp0OUM62RecoLCH3qUEeeV45yH64App7YEoRtaBdVezKZ8my2GRvPiCuL
votVgZudSE7kJ5+tKjofkI7wyi3VkzNqB7G+ikjBFDGENy7bGBQvQCEA/txT04xL
22JGHxDPW3kvT7Btzm0A31Cy157KLXOIS3M2dPuY17csmcGFWlg7GdtoXVGSlshT
jWzrpGqXtxrVfYBd0+rK7uvH4JvjJbW7dL9aA169PG+7QZ+89KBAGORmNb2ZMGuc
dfYXubAWLUVAsbC64hPIRrNxRGky1FOpMe7oS/4uGQa0ZrkdS8fyG3g6X1ncWcFc
y3HWR4gMv/ZAbkun+IWHaZQ6WiqIcaPqyCCYZAF/jMg/QHzrDCno4SMsWmnOi/m9
qYvbyWwyNVQgAqpC9II87S/Ur9guZzNGwTr/AHTMYdeBnih1i+pgoMLxGR/+jLwT
Ym6rBzrWfEB/nkGsfkLBPzAjp/RqxAv9eqEVkbQR+6lRYivLKVvwEUT8B/Umz/vZ
N6lASy3JjlgXQhnWSOPCWFjZbVCKgbG9yMWSelFKs/uONKTCaH9yYMUBw44wRyPi
ew7ZxfuaJCdXKEeCHEjNoxz05Oq2/pFUa7tQJWICupXE9GMW9g/BeurrhVyHXmii
NREgulADzqgioYXcsNENEd87pOdyw5qkIG/NTaRlKy/dJOPBfCjsUAcfEoJGilOW
kIY6+C0QY1fduJi2cUJUOgqnqXkN6nApNUlwER2xKae8Ah0JqnBIN8reihnnr7wF
ELXN0LVNmVM+vRLEplJWXSGWpQWFnXG1b2m+pg67O2o0ku7oBFULpPnyoXimJ1JE
KvfgpDg4cYjFM9kjQMSuSy4MH1cjmljmV7kQThDMPtr+xbbrKbWiVXLXuPBUjaUx
/ADiolO/t72ZTnch+BUAltVXksB3XEyuCrhzbrGRlSvIAs/qsvfySSPefsVx1z+6
Z1qXygqeifFHny3A51PkQvsCNhXr/HUjHGuUXutytMbXDmjUr9tD1rfgMOqkekVa
8J+Ugj4ajbA6IjdUDkaXBSltD5PsEAeGbjXLQo4uz0hd8wNpD4erRpmZ/Fg9OVfO
bW1tIaakhNHa2ZKF2x6juHIYy+iVCi7NvOJ8KlW+LWx47IbawDaVmdP/J7eL5Yk7
ovZb/chZWarwLKsQwLJX2a6N9woeDm+IpRcDhbRdnuXMh/CtuMP6zx0f4jJe0t9m
1Z/yfdlnENU1cdzkSl4BTmH+pmowGcjmCQ+Hp9PjPEGV7CZ6Cmm27dBwNqdaW8ec
/VBYI57INQdo4MPYZQDG66+4Gy5PV5iufP0VS38Pz9PE5oqZFen1vUKiVu23d6cK
s34jEhqzniZSimWIcvwtApQ1BUPPxnxfpEuHy6Z0HjFviE3ltcpxLL1TUYX133Di
xyeDMb6/A9H29Gn0HVJqc/OUHQAW2Zo5osvnYXSLXwKnwntJK7uZyWbkU77Tc/X1
Ke5zoyTKSiSoqSul0LmhYIRk1CeqfM3J0agT2QC/prPpM6rHMjNQFUYD2U4Sttqf
6VWJsSAWluwrY0Y1WDROl5MA+TzzIY3nYiMUvEV8gFLF2gQV9ck0fTgpvqWmuWmn
6Ssu8qf68bmJRm6qOBvvYFFp9ULZjxYp7rEMN9nfV59ArVJnTLzlek1BHJQM9C7i
yUwLXsaEXzuHTmMlW6Vuk+Q9xaa0xBwCmg7u3HIEn6TmIxSn4zHu+UEhtbNbR2Pa
33XrHroxrEPzmqdnE4TAif4ERG7pCTiNmGBXC3yLfVNOLW6UQlvLlZHoHx+VlrvT
d4PDT/fN8FW+w5TZRoQYXM3QJDdOZmmZZ4t85pNpdMsBsZniputAbJo9KNnEtDhh
IdkPRY6iVjesFpsfcR6a5OTP2h9x3l7vbPrTUcK3+jzjxbrbpcDoohMxO/Istovl
xL26mKPG7zoNntQmL3OnBchtJv5zh1XHICL42o5XSxgjW5JjFatqQVD6dATWSlmt
a9q/XSSubL2mPjLBLq/g2ZniGNxr0bM2aBE2aTqltM8B3vJs5VfdsEuw7KUtfeFM
hI5vZ9Hp3drXcekgvMUdgYfolqI4TTILqfmlCKbKYDNaCFEVnswxANapIXGr4Hbc
9F6ijsw9z05Cf/Bz4zUffS9VlZHWPgIHpNDbQeU5UqoSJHwl0fArz98naXCctZDI
tsuOy6148Jv7z+i4rh+jgRyg8I2ykAqdhMwQwdj5yX/NSi94UEpkh9XocVpQD1o9
BvW2OKkU9z38NbkxL191V8hl7x4xe3Qi9G+Ftx0RxVWKSHfrBN2qT7CKsR5wkc7Z
Y5y90+c2LSTDPV1YZty48m2fJm9+OHzO21RDRMbGpmhza9HqnQ9TwKK9WTZaeWdV
LAznzZVLDxG+b0AYKjx7LLaTNmuc8j9fk7ocYITlNi+q+ViinAyWGGGXnA7dQ1mZ
77eI3rqbt6RvL2wNmU19juM8W32222lxpquIESYa8HyUrOVcZHx+nwGr8+zri0yT
VgzApNUVvHM4CaWPVaw9FHwL0N2RPL1PSniIaCmrwbJH+BBK+w9meGApXtYN6mCw
cpIIY8CHS9NutOuElG3+q6ZfkFS5kPIOgn0ORAXWIlLEO7oHPQA11EbY1mTYcTwX
FhZJiHRiTS/1wJAn3Crdm2ta8951tyD1EnNceDztSWR1DbVxbBApwKfYKZs6vKhd
KKF+lDul/zIQzK2JdWtNSmV2IYVqi1tK4YeTf244wp7/Y1stQA5XtMGJ5tMaaNc4
+5zA5Sxv26WZICDwLRU5ztmcO9yMF2qCuWoU9OdDjlCt4ddj9+x3J8maXsJcdC5x
GcR4G7AimsNdNEy2Qk+d0zzVTgtZaqJKckwXT0rZu/SC2b4Dq0jj/e8pLU6p/0dC
/w6PTTVYr7/hyJVe+nQYJH3Ju09fpQsTYGP1ap/NzsAzEdHlhGR7PF2b6/UgPPTY
ayvuiff5cWv6+BVnNCArm5c+N5imDzj60S2AdLW4WyFJIIZTqi0b9tMwEjFuFN7K
OmopPvsqoK3eeQ3wit1O+ceTF/f6GkNJ/AiYL2BtoRnCx9Pz/6r6pfTvK7Vh7QM4
R/qG+luKfgV8jMcahf+1MYREzYRdbVyi6KVF+K2ZHWKqZ4p/FSpoZ+aJ/4kzg+Z6
2NHcA1zUeRSRCIEQegAML9cTpHUaCNggMdGOFb1G6bVCSs8byluQljtD7Qty/YeI
5vmqLF3lLxbwfaRDVrJHNAz7DouVch/VWFyEPVDqko39mtCnM8CongfDn+s8DMeb
9WniO1YEs9W0LtDsx4NApqdXNrYqW34GfHPhJtWhFDU85o0i0lybTfKxVS3zPMNR
V9UE2GcoPzNNAdVc6KHN8FJZ7J4w6kwpO+s7AwTW7rUcWWancuogwg3wqJ5Hmixg
55c3MYbZX9JZcbYKGYIrWoNEkvyq0M6iBnC/AKjn26cXlvNbjqcKaGw10W9bnYEZ
RWddpb45YApaB50vAjBJmx0C0z+lOuneONE/G3ek6HAJnSrPrpb2tWjMi7spvvsh
+Bf0IGq19RXpdW6BFvymzz9H1tgIroTcA7CMiWh91F/bM/ijZXaw9/rvL8u1yDNV
pcZwPvdjpwsE1ZjGj4/X0Nb1O0h8953+g9SZ/dqBWxbDizQAwm4rsw2NMHcMUT4J
yQNQOegivdwnH+kvfLxK2mchfd3HSsEbsNSNwHcIxM+DPDjLgs2TuZijz4WBwdES
vUWYQJhMb+UI4HR64cVs4fMEYMbOBd3zZ25KQBTNTd9DpgJmawC4NT45yM4vbVuy
OWVTeSMY+9lXDZba2VHCJvHwNORAS5en7/t57iK0YgmQJctRZ54Rj8NgFIFrnq+l
8CMT3QCio1qBE/tSOKpkvFEKMwmZvZNYsJcT7HAzOHanPy7DTTdhdTEKIjXr32ZL
sUasSebeLAReW4g/feqPYyHHrDtIhbGxuYEy1YTR9OsJScgZgovWfPKU6KWMssle
zcG+qs5PTqQZURNQwESYDbvsYrqh6X047Y13VQjrN3SsdVGW1ZnQeUIb5UyoBoOV
w7ajaKssC4gwWONYha3uJQP2V9aM8zPFWRDrMBMYs9WWNeDGcQP2thg42TDmf6p2
HMhXeKbTSIDMDEqOUVi3EAdscYHi82c8Skf5orA1fGc/ttDa7NtVA85eQ2OslFF4
lpp32sctct2PO0zdX26FzKe+pEUhEMskAK/MlULahJIiOoyh6kjHQjLfPDIEAbLk
aHK0FDrSx33Z0Y3280xwkE9MjDJ3JH6Z7n4jjC9RSSntjVnMlGsPtSXw5v04OxCu
G4tjt51BDwe7gblpwg9eGvq3B6b7IVnrWzQWp3t3cUHeXqzmR9tR5BvZ59oPPswY
IdsJBOtkZGRyKG0u4H3RC/qNHUJRgQFsy4MJYM0wDetGQZtiN+2f0TwAu5tz9TPE
qCQ8OYso5MQv2kPJSNLXrTGvDkkWUvuYvRObzbU5HrrsdSAPZJ1UVVQbzWrqXPl3
wNzCwqwlSR8v7iVQwXfx4QxHo81elLx2DTyq/TzAT9poimFf/HcNkhRFWYV9Ohva
WqVC7LahPOH7AZtSTWUb8+7Ktj42SZ2BkbBYqQsIj4GA3mgWTOJtqHhwPizUwxom
UAvr82qFrtxlt2ok/I0EdNmRhGZ41xZw9SnWxuBtqJmuRrR46YPagUYGC1mb3pkp
dKaKs2zN5TZ9LWCV9nwzi67Ni9mlhqvGEWsLz9YnICOkQtTmBvyF2ChHPBpcLhAe
n6R/G0430NH435/7m24PNhMBSbJmNadQOEYwy3DUieNfYqsHNtr7Wsx4r8CUNf/q
IKx7S86oIqk5is2aH3qRagEBkDg+G1ZNtPxXUMHWRQckH2v6o8MOewGtyDLQjWJR
nEZ0rp9wQJBKLwftRPqjYZsJNG0gMfp+aMPBlIRecGXkZWYaSZ/z9/IOeODBmdQc
07UoNbiLyLSEimOzKc6+9ZEu8GUOEuUoULZxngaIaya1Z9BSrvXP81W4JisLVSuW
+jDP17OSE1/BhBvOjdRZ7MRva3uYpC/fJfQIF7pkun7TfR6lQBNx99mkvRpW+EmC
/28LRDIaRjrmq+uCtxnDw68uh2v/tHBdaj9cfcUz0nfINZPMtmqz+CK8r/wDW+9Q
z8sT0vJ254RsoAdjNcFVMVejVNLkZeiVXWgkofI85L5MhQdXkxLPOaU8+Mh5pFW9
5w0zBXegGNJJDgK2DCpusD8os01sV2wlpjmguZ4o0YX2tfEQdCYn2AsUP5zSLEbV
mw9WUhfJ9qiQi1EJDHXlRwok5d4OCqB530gvn42PwUa/iJ2+jw0vmT78vT1RYEKK
Wk/gAxPiuEhAprxK4lgegV2CzQ9VRC0ZNNs0huVq+arMNfChYQVeNl5iHr7RHryN
CgBJPW+laHi1NgiZ247fbRmkGhMpiUlQyuhnNApnClmI2NR6OlpAQvuqp2tawIiW
heYbxSX1I4KxeLmu3E1Fbvj83c1/SmMS7Mrq6qnSmQdpUyEE73NgpuTDAmlT6agW
4h/dP7O1sybAPTX0vlvG5XgWfPBeMQO+F+YUvjiFj+ZiCGkuoqSJQxJtBsN3GRQ7
vOWDNHhKI5rypRCvCR71unxTdIy0ZY4JmfXbnROAz4cp4ASbelf43sY6xyWgdFlJ
udLMTXy/kp0U5KvPa/hqBEQ9eSRZRC7bl3/im9fQsM5ZDH5aEELAVH906+j9TXgD
wIkD6uFZecgnNPCdWHosAwRqUoDH/bJcagQdNPL5PlbLUnWIdrflPrlo3E7LqIFe
Zrw0/GAEUcSbqCkvre7g2XWqLPnFNZF6EQoENuZsJJiuUdo0Wuf9f5CESwl7kUWc
mpRTejZ9bd6mpi7m+tDVN6YZlwgxYCIwvVeLLzZ0+4h5JkMFMDk+5xYFBq8uJq39
5KToQgKi9stDn4t7V9/mltunmZPihQZUfMurfFLY/Qd1WSkoRLGX/LGIfvxPHhe0
YKUP4fA/WwJJTPatbc1pCrUm5qe4pRps09HIct1AheevEx3sBeg4/gPyaY/XKxjW
cGpHPL00mKXNSM9TfQV1V+EGh2lDPtuCqXz6i8uA09Sk8lbh3zCsJ+iBGFjJWAAb
7hR481WZsOsWDFPdCK67N05cofM9ShrTU7UzMfUw/BCvkIAMvbd+2Y0KOYUSEXOi
dCQP4QiPDaMwT2FKTmoVID7egqsI03SacdmgwzuP/u+5+Ip+rQqQmAzeil+N9uBH
Mpm8xdwNZa/+L3M12bl3sRDWKgF1/AR7M6X9BUG/Ux3QND131rctOWovmetigHVm
AYlPQYevxY2EPiJZ/M30dOC/s5m0R3xXQv8SMEXU5I56Ci0QQJCsF7SHOsLHSFRT
viuaAdCJB3XZF2U7Xm5zavogrwvymok/9B/1DL+la6VdX5XPpEBnoEpSzR7k5lHY
WnmK1PcRFmBvDAG98MQNuYacEbj5SmVje4vitIOxntGPFEGbs0TaVELWPiujTz/S
DIEDchyYyl3tbVc/jXW0fMyUTGC9oGZYaEKxmPti55GI5FV1wfFX3av+457yh0SN
xGAiXtvG/B+889JbZIW/Q10JvFKAIwXUCrheA3O4H4KJXofYnoJ2uuxnAUIg1XfW
iB6IqoorIfSDkTfu//R7lZGbi1PKtyPBOC45g3DXDlVh4ZlvTVk+C+7I/0Y0AZof
tuREfCI0E1JaVKDhSMiB6CUog4oU4oWlueph+MPsSXitxrKimPKUhMzBF0peGqpM
f1A8166AF86djsMClepQ52kmKKEtRspGd0ee2xphY1G26AxW7Mav6nea5++gUuxu
zFtT5hT5wAUO736buZtkktfCwDgpMpd290whv29wghAtOvQWgCbD09XKJQrvcvdK
l3x7LrzeDED4VsJ0rLmfup1uPdflBGfM4rMqRWnnkwxn2zL0YrSzhexUnajx6E8q
cplxxwzgBXtwUuo+k9SDoHJ1kvEF0mlFa9ywDLld0BHQrUVwXy72i8gB7Ynf/X0m
Dk13eMe0Q++vcuulFDSRYOP3e0Z8q6LEIfNYVE+nlBikqc6q8HYvNzdpKPAkHoDI
jMuhGcY5XsRHh5q7mswN71FpYgb4P3qhckZwk6W1Z53vGjx0TrrD/tnS6vCAYT5z
FsYqpoLqJzQ67l5END+IwZRNfCJZF9ra6FMIqwGG7cMhFt7CLyQM3i9N6oUFr8yc
q+TcRRyomVuOn6LgJ/fup+6O6HLeiK9afZM/3updR3xwjZFft5pbUayHWR1PKphe
aTRUtfhdc43y0P504jCYCSpoLAvEQPcq+Xxr3ZbBXKZwhoAw7U67ZjYvJAINL5Kc
p51ECrQQkvZwjVSNwT8ZyTwia2ZhA2rNhxvcaH+AOlTmw9vqZCLz+MBQ1o3sGTBi
RJqCNGk5SUrmm345MvbKFYUgtd83drAL38P5N3/ZJJ9e6f47aGhfJ5CmNmH3C5kD
FU8hQe/JAa4wmcVPaeeNaROZNo6LfWR1xqG0grzeNBhN1JY8jXxw4A13PcHNkp2Y
kYvmPRDJaQ1Nf/AMi8yTOzyPhZMTivtGFkMVNFOisDrr9jFSDM4wjaQRtoOvdTuy
wTd4gGd69b1LPi+E25dWowgv58i2hKry4wRNZmID8aTsepszDzWUoogyiCTJZ1rU
KKJZ/2mRRSmL++by0Xm3HZrKiwtCNUiRswcBl9OX3TVS4m5D47HjMRQNZ3pMZKw4
sJpx9FI8wPHSEV3/Lx7iu6qNWKu5zYfJE32k7Ln7g1sWIFIjrQSwjkR3UVaSf5wb
Nvv74ExCVBqMybe7b4kkV7djKHQktJaQm1y+tDvLuaa1iZe4du0aJ+S3p48j2gQA
xhWvWAN6+NHFmPOPEqI57klLWTco/HSUQVOKicErb3Wlx8okIqUMfJyuGK3lVxK0
tcPiS7dsDWDn9awDaa/j1lJecNmDanWluoB2ZzQKxBdc6NmLAyUD/UHuoVm+ihqS
pavkqyBTJlPLqmGS9ZfBw7/WOuLTxSB0757m1WyML18ZvUWb5qKuwPXetksqXHkU
hBGz+4Lb4oGUbaNpWMjJHdK519EAy62MdtHfiLkItAFMhBj/MA4nJ2nMa5dktL0J
v1yVRyN1rqkoLpcMPhA8q8tQFCE5oFtGoTaj1K4UlgfgJRlG6e4QfnXJvUb6hXpm
qWMJHKPL4OGNTCh+16Zk0sua6r7J2oMN8J5L+XvbtWPNHlMQgLgSN0s+X38rdDRA
1XnEgGu23ykLc1jwuYY75uAAJTBS+sU4Qs/3s9dU4lR0pc8DPf1bZO6TmTPz3qsB
x1i1E+c5GtX+X8bpZctstrFJySg9ZpEB/4KgtQ+mf7t2q2bmX+qPRB6UkDVanHrm
aJ7PZRK/E/j8rWUr0ve7Lr/U7eF3IQoW4uA75DTpDJQDEh327lh24Z5HwLLq2Q+L
2vA/bdTEaldPXAuBw9uCDCJAmQsbxDn535j9Mks4pvLkYsCxm3QjPYSw9vtoJKV4
zYeWxwWSIPgG97DFBgQqN28ml+Zszal+VYDR0cs0imrAL+GAzevtIi3LMIsRoqKP
Sulai+W98gOLo5c4EZfdQeCI3D6qVz2JmTDpkamIY5VaY6pPykg9W7hJZQ+duU5X
eQafGPKFjCmatWgAp0WKh590/Wl3wEgvlfqOgV4VXuoCv7WbuXj05MrApdV71QLA
SzaYJtl0BWG099AIWnQo0R58XlNlT8wB32FhkTrtgCgwF2OIxOzGj3PTwxfpzR0W
M51//2A5jvSpVjwDdLZuNRODRN+EIMYZmzVMqv3fNYlKMMg0H2He8by14J/4p1LB
bV6ZpI/t2HFF0fDuCa7vTSO9KAtUitPD3mV3vHpE+ISl4bCTm+MfWaYhBLbWDjU2
WIZgXikXrVkCcTT+KLa7VSuVEYx2KzTWX+yFRX/7Uy4NkmqdbPuJwBxoCjlK6pfC
hc5TzzR71XU6PbBai7f/c7YvE+ZUrn8k3V30f8RdBXrk8mRszecJ1Yj1vLQ1ELuq
GD4eERLxf+WJpVb8RptrRKiBHE55cum9XY35AUxpOO1nIuyDs1iqG3Y7u4hmUSG7
3ol3oAVvJGDqOWYex5aTBktO4+PaGoFF8rVDIDWRQrAsMe0fSqNFCU2Yv7XChUx8
5nOrTrPBYsHlVbNXskQqX7MQJ9N5BtrfmDVVVpL8wW9qKB0MsiPu+xA9YPYpX/7S
7zzTbK0B0NjSXf2QC+ZXeiUEbdzdYL/dYKEXydMTK04WNdokZDKhifjXIq2hXtsv
UPhiCu6Waa454m/PbT69EdQfNMYnHlud/7hqljr07L37OTdTpctNmed4F8oyN9sr
I3DQFLsHAP7xcDzvvqEJ3hYhul5UgArypxF+MV/udUZneaxlVANJ6X0qamVQE1kw
XTLWEShyvqk8/PSBVubTRZ/Wkq/y15KdXVkCUJ9CWWhVL7oQ9mI3b8F6FXilu0U8
qaCh/HxRmF2fmpJ+xI0qHBd+V2wQworgUwQDUR7DmNmwVzyYCwrW3PXskYwqR3si
m/2YEeXGPP7e0f5SG8A8kdVkjGu5sa9PhyvwdezLRKxvFTaFhNfm4NIFpzCngi3F
9C72cMbr2AK2YyNLFShJdYL3WLG9UrNL5M5UUXRhRnHk8P3tSkg9VOw3Ufh/kNF4
6dBMlQqFtYcQKenvyfEqtVjS2If4RGTQDBiKe+PgDs9AXAUs/nss18qh1KMbBzen
+6f7DGA5Jq3aGPMQv1tIf2P4e+rcN/H4WqcSk557hvSdew55MboFtCW64byz2+WV
uvIza8Y8nAuHmrs8EyAbPJhd0yf0X4NPZuZScoFUe3WeF17/ahJxcPreV592B4/9
Px4FahsxwEReXXt9AkE0atsc9umdzO52/12+ALSWx/QUEKZXIo8jAH9/e7Af4qpN
m5kPIiej0eXW3wKjHnpgakDOqhE/MgEBpJVlSHBNAwXVWer9fX/WszRMcYP36hMa
TA1SG16UKT1WrqVORVV27TDbRJmb6ddz67q/X7TUtItLXgCSnqn1h72zOSR9IfvA
Jv+oTQklutWjeIBx4WJFpD3ws8DlX7kqQKel2Xa16i1zAovqHJpPdx1mhs/TblMI
5deFZrDyN/CPv/31ILrRKsVox249mJ+wVGimw6Y/cDuONIUn1RKSQyNAlOBt3YD4
iQRKkPYAL20ejwqMrzJ+2PuyDP+K3TJa8qCVF6bKaITrkfUdcbePtDrqiLIRWWLj
A2CdI4c38YUJEsJpSKkzYUv+bVKfEe5L9QIsAcZDvt9ZY07JNujOWx4Mig9UrOrr
wF3YZpi8UflUNa4BXlNV3L3tE9iuzb+XLDH/Nw+Cj15Tt8mIKPqdCDaqdLebfhT6
XkFC05ou9lwpUtHFPsGoB5XY/NusvLT/NM+N5xaDSFEt87q/+IEiOcJ+ruJ0QEv4
rDBWtE9qIVkjIFSiry0xmP+IBYaf18CoHJkrHr6XsXfSj0I5Ra0j4fk6LCiaMcyU
AN/soUyklzbn42OVlDtS4YkYQLBvfYnrU/VTBsHxzDHG99lrnCxxwdjgdKwtsp2F
hXgKaUT0P2qJG5sByENqPBb9SKoWvX9Z5+2jvTcZJhlcNag8S+MajzEyigN/3pIQ
qK+OmJ8cZCy0C7dmxhpmhmhH+6jSh8WrgoY2fa9m0+bkf+QUMT9JPqnCX5vsFVeF
wZpBI4zh8NxRx91EnMWWh4WfXtypAuPR3HEcCV7vETtnaYUkRqOZ4FZ3vGVY7p4h
UCVr/ULKlhxcCtGYO4VYgVge9IsF3lAwjwFPgu4Or7i5+eEEV5rLU/b2AfQbsgfF
vfFBXaWpPVpIxxzf6OGK+oBLMofHjIS9BLOMBiO3hfO1WTK6IFEIn+o3giFdGqwm
Q2XqyuClF9kkcV0rejY/JK4M9Zt2vtkNsYkho5AWYY6rHsV23JgyYKe0l4nQ2YiA
hphIk7LfuKexm5F3520Ge+tI+xK1ijcR3kI0yHJdOfAMm1bXNIaUfIo8FhrmCVYx
CZmFShJ22GmomjxnVrxXGlMAbaBoQkCqqRKUKp4rkiHtz3TjrUWzsnzMERXpdygT
f3MsEZqxjUqAIX+nhqMwZxMgqkGZn8eor9atLTzEpLbzGIpFhNdkuskGSlIX7vGx
s3jaAiLEG+y1IpoalrpcKjV8seHGf1pBYUFYovrMh4HRyOliOMDH2QJT3qBV/WQj
74IJDsjbzu4tr52mTkcQR07KYezOba9T7Cb3wtyMaTfHn89gYalUH1+wohoWuKTB
BDivgFmpw5h7R0WZEZUsODiyTL4sUODDhs2xRF+uiqfNCAW4lPKH13YaMoHs5rfZ
BbP69fOYJ3H0uf33bT1nunNF0aThWmqd35qF1fzuI2p/V3rW1Jr7lcRQZ4J7VW2a
YAqnin40UmVUKdcOEvTVOUr2jYrfnM3SUibo/+O0iWI4Tv3v29eLmwUtlS232dEp
wxjmaiavaMptN/Uo3VNoQImPRAnDLsDhRe3dtwe2WLpIrG8EVcluGsitUeP6e297
H1bfigI2ExbuuxxeAuaauXptNiFtXt8vXQnC1dc9drhSyW4mX5XB68pH4TJ27YAg
jx8r8DDqbjby8E8Aq/IkIpulvWPkvjbCl1+2tKcxsIMKLpzLncp7cWqEgY3usIUg
fHP3y8KGf5JrcC7r73XvcYUOGZe+PTkYVWSGORkV0vphBqZP1go+J8moi/GH9xhr
ni096in8syBjTVDa5XnkJTkP67v3f4eNOJ7Rx23Becnf8yqjYBNyYg2ufVwSoaDR
QQhmZI/3AXvkLAcHESwouCd05BJ81P5xLsd/VWvrZd9stMPoaSfR8s6QnNiEaTND
T61gEtcTt5flPBms6hYUTkZYLSRKOkdrSy+LJhtuqR3T5ClRqP5eK66pkQtd6Gpd
HjDl2tnFyDzyyFPYPXuuEqexLPGcSY7syogUnFblUvAsG5Uk/0+HdifHYb6h+5b0
SKQ56ppzD9X5a6jMoc1Xb5ikQhJaa+5RwXgVDGe/a3JUYeKihfAUvuHRvDV7t2Dq
SZzF/wyAup8zdQbwb1o7B59uDWHM5qUQkckPBhuGlAHWZikZfhPuxxfpK73XiZP7
vnyDNAYTcaPrrbVyKl9cS8K++roXlTJjt10UFyMf47LWozCWbBibCnGWHiQlq2sa
AlhDwHv43Cg38YoYDSAhwrAxJeRun627tPMe8pulHd3zcviOt4Cwe+sHkmanTDdO
hSJbM26WVf1aOW9R/IpP2TQyfpiIujxHWpbfMCJjMP5JzvI8TOLoBWLCGq16mz7j
i8tdYeR32cyG0dCY3a0UZgWGbHzwqgXIViHKxCI4t3/wPLf0lzhjfT4F+H+1m9rq
q6u1SM6pXvqrZxDAv5iIruU55AkV5Q8HaTkvCf4Vr23wEEt9ORvtnSsGMZXIZrJL
sEgCW3KFUR36vldOrTk30cy1PrId5dRYTElhpefBVQpKACYywH9vOjgXBylY1Il/
sRf3cGztHwL26+uAa3jkp73alt2yi16r3bz1uGZyIJBjECZgu8WpVkLU+exfnqaR
PX7EoljO3DtenmKwc5Rsnr1smtPDGmanazDemaAIJqnKv+Qw5iuXvfwbtCt8iykn
o1p2oT0584PZDM/FgcX3sas3qZ4j8X/ANt15Xl1FyvS5awO7hFM0QGeoRvsnFbvj
QTjoAdchwB9ssEJCbNEfhaUGunANSGz+Lj6PLZNAleM+3mB92e4YIGFyl1zWR1ym
NCSUiy5YZt4jsHU+PO9jB1pyc2glQWaYouHdTxCFQElcsKhhRPGpd/bFi2bt5dPY
bqMTMsejVl4GUDZMADJsKzYozJmYi3Dtbv8nmWVQiPvy6BRMHqqO62zRQgaifCmN
YxB2XTBzPSxIJRYzY+bPtvX+p++hx7fATQ8LNxmVuk928DZjh2RkhR48CMsow6c/
b3VLuo2RHxyChEEVdj9nJeW3ZkNv5ohCF1ogrP+3FI6eclOo2WfoL3DZbOpR8Ayr
oTV8jrzuoOfgkkT00i9fhuCc3XD2FPoZSLlzpTAlxoxHcY53TEM5teHZ+AyQqZdE
Xwl1Sw/Eun2TmhEIXAt2xftmlRDdLMg2PS+wRXPqkxksExpV00qoJbaFXIVViQnv
EAxu12pTXKV4HYtOb6duTPa/1hrgLgfQ10HgWdFSF70qwOShFdAz7Do4jpQsIbio
WldkDcREbngMgdilWJS9hfkcZ7Z1PQuvIZ0eDqF06kIQxozUztBPWQBU7ErNtk92
86i/mRXAcXcSMsAqZ0P42JDXtx/oP9YJrVXLe/I+3xF2i32ao8SaGIth8XDWIg+7
ujXT21uBKuJgS9tKJcZJHqin2CQ9PwqHHdd8i/wALIuNzmHKms6rrZRiuRkPOR7L
X2SgBmBiUqYcS5WtlGdG1yVXigLyX+hE8c2Lxxw09B3NLooSB51StG7s6mzmtAZx
C6AJhrpRuQ+sUJYT7nBkpX3gpWwscp1JDym9POhqd9zAoF2kN8flLWcWoV2bAn5H
FQJLT/514hZ/max0C+T4K3FUGGRjmHQFx1A2+C+WkB2/fQL8/yk6PqbQEia/F1zn
pwi4HtSOu02dGsMWBDGQLrG/LyBn+Dt1J8vcUWlfB9XX7G809c3zSau9FEqqfvTQ
dkr/HvfuChAV7esYlePvlSYDZWo+CUlBOF7ywN611BoCW5xNm9+Ac1ICFzLhXSbh
q/YR1luqGn4fn1DgN+4IMWwL0SKXxx1HkJR2HnYS5X3v598ZXfQx7EsgZR37QaZa
5OfPbYDmdJ/5UV03tpVyK89oLpe3xVrgVrPhhiRu32OGXDi+xUDwWz3siKGEoBUr
XD5aZNkvvCUEE0SxdCd2oVVcrg6yTEEi6sH8jOIPdfjOJby72+20e7/P8LwsBeE9
+LjoBGi4LOJbjOwoK0ZElP8B7ggJkDtKIfN9stxtSjHK1csUHXZnxhd3eZx8GqHa
LExAgqSTQ+2F2Yn1WrOgMG4jWo8mnK4SYEJs7z6mIsCkO+f59LCqONwcsx+X4DDO
vBtRGzV1I0gbgTvW8I6KtRmohsnJcLnGO/5TfVxQCVwlfN+7ThUGEnUMfmGnb6sa
SxckYDGI1RJP/ciGa5VXo65OJalBXidU8s3dLBRvl7oCH8laXEBh4ozLE+/kuEkP
xSDMccgl63+O2dY6OUX4ql1aI/HWBMNx92HGH7pgvq4fWHpfH7zPZq0EjZ/p+0Xv
mYY8dfny+leP/XJXV2omF7gjDeAGANO5a4GVXg3yZcfUyfUpK8a9HIfzBk7ZAxyR
pZzN3L6fV37LAtGXL3Jb4KK596sRI+eSSzy3Gfa6dWvZnTYhQnfmqZA0zobIoAf6
dEGiX7TbqCCNRGPy0sCaDf1OAjMSvQaQMK/PyCm10MzLbHap/1noBvJi1KLb5fJZ
yAMlv5gemCGGu4Yc5f3zTBaOjzOFl2TmChr54v/fMIQLzvxFwKPeUxAyEv27qVPY
7rACPeuzSjfyuVFimwt/TLx+ebIrTTmwh/phes7RlnAFDXhX5u3+cBk57MlXWjgD
16e6UrNMmngDSKuMxCi2cFBHanj3rRtBgPmIwojhlaBY3XwkvTirx1EVzkrUvNUV
dAaUV18YIzVsokSu3FsZ3++JjItClNIzoyixyRfE1ciG7/p7EjPivRc6qhKuS8AU
H2oFgbEUpuTqfDp76efkPKalaj4gyDI0BXNmusaJOZJlX7pLdXisbMUOl5Ll1HZK
337w9d2Z2pf4M0UyIxWt0Qw0k0okvr63b0JxtEULtmr3NtHDPJ0UmHZPev9oebNR
Xmy88rKvlge4X0kb6sBPPZ2/Abr/DK2PGQndcSbDrPDPF3SC5mGSVBAZO3o/Q0Y8
FkrL8UfZkqypocbvziDAihneWEW+kmrRksg5RGdZfqNoEYAQ1hst5m6vGIjvBpmw
wW4cGlC4jDf1OuWW1jc8eJ2Epd9Bmxql08zk/VetrZdnHgXQI2cIKJuF77zL1fAL
IcI+GWCL5zoSyDtbog4tH8yGfX1eNpgs5VLKBdgb+Zr1SALtjZtRGNhhjRRCBbuT
rt/N029oVGLzCVkTqDp2nlOcGljhhSfF2ZibzIIihmcpUAYDG/7gbdg9Fl1uf01e
GLXSVnUn7zq/7MF1kVZgQoSmQKmrxcz11E0l6L6/avVH7pTte/EHGvn22T1Q89wh
lF/21p0SrViLS4aeOADMxqV3DVKYNqWXxmD9rQRKjNYASh/2V/Q1D/eO7S+81dTv
1tRQBDf78IN68UK7KjjkG4xu+SUt3B2aTE3tmmQ3+bjwjpdMvsX1NG5jHb8+vp+U
w/FFB8HgvaoOtCbSYqT+Fwv3Q8oUkoLkX6Fv6z3wuFFiikmttt1geZKVvuTGa02C
ZvKSzz95hSVNHkOMkLQdvKicpPQOAT9/zo17ieOePibUbvDVz4u77FodFHbeGSJN
LsbEsW+T3dJwHEi5rsd8wQGJmKijNtuHvE3xFSM18jAAZPBTZ8z/lkteD7otlcN/
Cv2GaNs1GKb/oz3FD/ows5OjaHYQpniYZzPsoOguvoECH/oUvH2RbUNu0SUik5IJ
0Dx2BpZuoSIz6y/C58Kg/+WfX8DquyhHidmwvpFIqQz4q1QbOFbPedQ/3YvQ/+gR
vIfOuLNuA2hvTyCg14wLpC3jvXy+wD/kMQoHHCoJk/v6bHgmqKC8yiaPBsL9Am98
agUQnJDV09Fv69yOJwy332mAvDmzu4zk/SQUjFOC/pMQddUlawtJARZF0UKxOZEa
3u6P6R2FPs//Ux/IOKxuGwuOhYg2/qXnbkPltLbsmIBQxupJ80pOmC0Ircrl7E8Q
S4ePKHTxPPuQ/lSWfUjapF9nKT6X41LRTfbktQi+pXEWSliEFPuKjP+/dUTcO4c6
EsiCG5CfE/O62CxbU9quM8M2V4wyOjmh2eIVZM0zpaeXsMB7BWmQs1kGOQZ/a+FC
STBTdiT46Uh3s4wFX83tEZS9+86hsiWY6onFwkqf/skraJ+8nxmZzC8JL10epeKE
SS8/m9wKG1RBDpJc0LFK1T2Fe/Mv1WAr+qb8Z9TphTO4yU5Hh3rSKGwbdTTffLyz
Ua95N0ZebeyJYoIhXs7Y+M5uxl6U+OE8xaEKro9Zv3bzZoQhIddFS0xicLem9qkp
GLWKeqK+mEIUbEViaunO7BhlCkV7OJmLvLGLHTLmD9B/wGikT93BEZbcmaT48aEW
gJZQH+D7dl0X78SkRMjGxoYOMogdD4RTLO/+SEp3/CqQl6WSYE8qjPCNLaiJp4qj
jdm4r95yQXxprNMiFcrs35Q8MCKw5866qT5HC5ouFIOt/r7sneCF0fS6Qn+QAICl
PYAQBdenWwmQedX+6/Qfk5gC9OX0RrXCJkYQ/1TqmQO06wxsTurGIy11c3obITKQ
04iIWCLh9fs50Fuk6X2HrKp5PxbdCeNjUWjvOV6v0YknolxMsy11JbkPL3jPFxYB
ZAuDAH2uOi7UwFr7Ecs6Jyekts67XJbYTHTAM2km1Yyc5wKv8lmHJ+13y+hGTKIN
5oDXUSfD4YYLJbpi5PBJs0DxNi/DfiD5LIH9pX2WkOmlnvPizrGzry3au94sIXNu
1FEhKOLzIZV3Li8JjdHIBqUyi2N9O+M+3jhnDEmOSJRVbfMOZbR1zqRGSSvOFkoD
dxNo3XGfkeWdSSdcNYBtCGPNvcLuKLGfJ+vr8pqsDz332THYXCU1kVkGeu7LNhnU
TEwFpxdSTLiI0bnn30AFLQoTYcwOQO3Fklk5Nl6R9/eKG04ROLjmJ8X+znIEjqxa
FrTpKpQB7SbPmxJ56KcK3DIbG+IPLhlOorPn58NN2+4uqY9Q7lHuT9B/uaJP5u8D
7Cmd5JPKm0JaTUdLefEOA6P5u6wDaghKPccozNjUmNhbzId5tvn/vyIpZjc2v4iD
FnYbKzETfYofTGZ+UlyyBKJHMfSgktFG4xxg2cSo8B2DW6xFJF3MF3KM5FvMMdca
vglQQh3Jur4ikOmmHZnysWp0r/jfkA2qohE8pamdkFDU/EWDcS59OHjpWQr/0QpS
/h2EfNttXuh27RIXm4Smr2wEAW8H7QKq/7nILrvWevmn1WCjiTRicIfrJCfzAPp2
CZqev0ymIn3CTCqTr1wWMBKQwt2yL0dTc1C757TCMy4ncmvr+WrTpclF7ZG6kjyJ
Y7O82YxMXQwuT5WxCdFOifR89o81UXUt+Td+Xx2XviMG0yWAv0kmIOU7aU4w5NBk
06FupGbVh/+IYCZFlM7hUNkadrakP3ZG63tuo39xoVlfJlRawvsNC4MZqTwkJktM
Y8AdrrWwDU0dAu+px0K2VecSYls5/qu7SebuPOMjoe6f5AN7RAWNOFBAwJW/YOSB
+kyg2lmaCG+my1OWd0VvRuxZzp6n0TnMzIu/k6szjy3t7gtY9uT4McZULJPibe/m
ZCl5rayngcBoWoNpF8XbiY9s8WcwGgV985Y4Z3YGaev/mo/WAWoyQnv7oOG2x3fY
tRVQfwinAt7KaLnORa/6AURzIXmNBT6foYlSkfqCLI+v2tPIFeUEzZl0ey/9sGT3
EDzPFHhER3SR8JwNqTFPONaM455cEQ2Lay62oD2NcpBDOPxImoUDUMRsgnBqoUTc
3JNhvMNaMpL3sjNC3Ca2kfkrAGUyJaMveyyjh11bD1eyDFtdUcu2P74uMC1owBab
Bl8xYEo3aVE+2WWNYDVCnbZ3MTzNR/TyxZe+UyDhWgao5+E9D1eSrhj0wZv8lXww
OMhuoCV6A+aKlVZ00U/Doc/VLX2H8du43wo1HppoyKp9jtnbah4zBgKaVPmTQgw/
yY7U9+l+jkG3+kiXTcrJKoDMFGEYiE8jzlRd3+j1ul/lpl6k9lq32I/tSQVaeAUb
oM8De75NKN5oXXXKuyXc+5XZZVONoLBAoJhc4koZ2DF5n5MI/MzTJBxb9Iy4bjL1
hGlBIxdMKZStk+U/VBtg9P7cFOPubfNcelz4dMsmUf5JHEL4kVzzx3GWQZgjDt9T
EtOLJgv3TrKz0NqrgVLsgwqaTPm7E5B2Nv0n8kCbtx1V7JDOm20GTKB9zLf7mkRR
R26U39mUpqU2P2Bz968CTAWdTiiv4ugC6CvX6X7kiUa6Jujl3SbpccfWH+a0AFSN
J0h7gi62fieQD1eOCFhmGQQnJW5kMKdZrx238YEwQ2yz4OjhshWhvFghnl7/oOt4
PtWOVY8UIRSyrwvx2m5Tj9uwyylMNemZIVpJZ2SJfZ1i1nZbQj1fL2VrgkAfDvzx
f3Aazz0W6WcTkKxCoZsu7xow1E6sGZvyKGqPwHVGyPaSYpDxnDdsLPunDWAikQ6E
pE7Df9tvf/NRGeLhOJ2T90oLzu0BA3c0ajwMTqDGRaixJ6euxAlSyjGP7ihUcF2a
8aEcIGuqFoJsFVG9xyaNkfKPVydvVkp63HBg9Qe0PhuwWtBm2VIK2rd3C01ma6TC
l2pCTwSq+kRd3jP7/UaVP1SBWihYajatnuEU0RbU3AxP5xt6NJhsZAPuFcD5CnC3
8tLqoMzX+9X1GJ5mIBL5+6S4HKSd6qL6a2DC84I1EDtvtjNCFiJp4q5HixaYkHJp
V3vDeI/4Bw4f1SvJHy2sFYEf2CMHA6d65QexcxmkLbGClRsxm0IS2bRxblo5qvo5
JL3Ow/iMCSWdcscWxkJ2g9FxumZ3QV9OGGwgSn7fftUwhsGhuCbDC1+wrwbh3clM
HUzp2GX3Yydyj0Dmxm/Flgd9mhrm/Y44ArjmELMFRfW8D971vjJus2Zk0q3dHgoV
pudiHnUD6wTHzVjwQKVamWD8E9WZlLb8uJVMo/hCIaI/iRJBWW6mRRF03JZa9Aph
GvuJ9xWjC8uQQHabSB0FqzUudC8LmKtNaD4w2MqaHldTU0lVzLxRIiS4gAjrAGdU
ageP1+pw52+axk3K7asNnN6CI+0vQ5rcZBGLDGU5ccDCj13d+U8/sIpVRcFQoCiK
SES7w6PK3lLutMBqdX141jWaFWyw22t593TqZa1RcACldK1+dVPQGq2brUZScstX
xkwOzDizZYcCD6ITeB5I4womlg3c0MV3Wxo2690lihQsYBQW3rqGq+Sik1hl3kNT
/kxzzfe5vOWhpm4+3YlKmzZGn6Wbil5xoMTJxaDAF87YHz5OtjiWyKx07KbrgGxH
x5RpugO+exvVb04TG0bCXnpNOoHkokaBuvkVhPiAszulpx7ZYlzS+v7U8OLo9C8N
XvXnIX6Z+QFS5MR+IHccG3B1JqIEeiSjZJ0X5lbho7wNTYixiN8JetWIOAyM9tqt
k3MAtAITGPPb/NEzG4cQeOaTLbMXxboJlIyMufJQqL0GwSu1+KiiHct4jHe2X2jJ
KEHBLBhZPCWbNmhAMOwFU4dhuhi9e3PiFc5wRSJ+JmED+NXOHzdgvw44EzR7OV5k
AL3q/wBA1aMx+HawGGj97VCNUHxCWab4s3SA7luNaflfIa86fKgRQu3l99m4UQRw
VqZFVgBnFm+wk/Di6di8VM/1Est42T8giHFt3bQJtMMEucRSqXy5craQ1B1oAV7g
OsoeFgUDOUTjvghalXbnoU3++y+lMVrWueLE8DCPawPedxAmvgrHo11fdVkcm/ER
GpXxUIZdmbfpVAumRWcVDuuUAvkT75BPQlik09zSVjUlUh8J4Zpdog/cNE1avgPw
1gOiKgWyiGBpK2kDlDafmgPrOLWt9Sh2uI6OEOlT82SYh9X1f47LOjZi33WIVJLB
fmj5SKFtJxWovkNVTesTwMZ5LJdL08cM+PyfpSXcKSxztTTScAMhMSiHEqxM5MUs
mwRSob+o98Cdc/TMvoMNsSZAIQqzlGzkYakJGOEvKS8U8GWRRX4BD7ZM9hAQ3ozB
rRwdmcetNnk28PYIcOp/4xxssKnPVeXNw3dfN4OTI3Pxp+ngS69tkVQ93jQIbfSy
OAzevpo+M0TTvIT5O8q7J7YxpQwtZSVmMChUXUqlF7JCVAzCmDOEblBja0r8W34o
1crSJGehiF07R63pk69XlvDSlQgJNnWN8wEe3G4mCclSOmkUQjr0G0CfqlbPT+1Q
l2Dxhy/Pbu/dD9TKkbw1sjlv7C2NfunBpae8PNIP1OPHVe9x8hgigTflH020+urB
TpEIjFpyS1e+k75S8m99/u/JNTp/w7zchK+dyDFW2IpKZT0MH9RT7fjWenIAm7bE
zmfiQGD6hSVSE0pnUZS6Jecs/LW4qofp4DMFfRh4I4VyHlf5cvMogzoTOyw4eIxL
vTEv+2uNK9XDb6VlbYPw3J1kpkdRj6N2Q6AaeG94GMB/k54dXDgC7iqHMcjY/giF
E4MTf/5WfSHsRfThUFkA+eBYPHeM3q1p7mwl8nDhBbOlkeVe8SkzFK/gTpT3RMAQ
tT5Gm6tfSVEkz6rUZtFDX5Myx9vyMwPwozmIq2rMSZ7bmy9FBWAfvBeX0TUnjzds
PZgEySrHJhtAGMte83zZ9zY2ykSjGB+ZO+/CczXq0p6VQjHy+dOKX+djAttSKfw3
Z5/zvFF9QmkFz1Zcmuxm25iPb3QT5kx/Fxj1cmfhOr7Qh8eGmVTpOT0oKYxAzhRy
nyACaV8vu4v54Cm31gKMdZozk/HPKrgcJJOlGT+m0CcMODqpaZL7QAyZe+yJxnD7
KIVLTGBedJ+tJGVmQq8XOFGj1bCbwLH839tH9F0aCU55q2Cug4rKdA+HBBHXCL+n
pj8XPQu7WOL10cFoW1KhY8wFaD1cHTacHLulnsUUJfM5yhiBBvmBrEwcuoV/q6ra
jja8oiw1gXZHGNfYmW5g5qP2b/4CqHscwG6unCoqN2Hj/rFL+lbOlzJ0/2DEZEOI
CqZYpnpzdMetPsnJAJX0On94E+nAbvw4UjMSS5casRnIhdR2qmfEEll+oWzIX2cT
V1Xu+1NkwMvAXOHacvNbNgG4Iz86k8LSrLpQIl+AOcUeZuEZ6jOdBEdjCBZVD/8O
G1apuSVUP5TqDwhg8yaUwDWETj10WrkgRGNmvutWT8zrrqLrax7qnZpZjNkeYMWP
dZ7Y4lQlgjxiFxpOf8ElKAi6K5uz2ODMeg9eQjb3skgA33EH6cVc3wIm1/sKNQWe
y0qLMvwPbBwAxNuZk4Ur7+aJLjgpn7vyWWwV5gQ+bLDo/opRKp7X+72cqc08QgiU
YcSUiMLlMhW/vwczsIto9f1bsf1qQWylHFXiBxRpY196BETRcQNTGxCn42qyoxX6
uuMXdtkY274HMGg+xx89BTaKD0DrsSKsEHaMfqCklq8NW1RiRXHTD6/fWtVw8YMh
6tQ3pbLG3P1I1s8c/uovqRbdY+Cm8z2D8aBkJoc9L67IpjI1bfWzjEwny64aIIsC
T2PCHMljX+T3OnkvxYHwlHWw8zT+KJsZ950MC44cW/kAbSoXevTIcWQMEnp/PHVx
3Q/pwF8e8042OF9HBfuzEHlDcnO9Ysroekx/k+LfMzFcsy80DwZejY2O77Yi/2I4
K0NEBYXUmUkWejS00176wc/rwHFX38llotHskYxqFUqjjwej6t2ZCpPJpVvCR9i/
viJciu2zWBX7ieJhO/HKzIJqww/ecrBTzxXO4ZVo+TNfrTo/SUzCwEOceg5fFlTS
7bciAfhqlvJnMeKBxgMGtRYwj2dCEDl0S8Waxoo0EzIqaFa3y4s7vdBgNidS+seN
OIHlwALYLOAlyRf+FpMZEXl3e7EeB5DJbVmjKIeI/IvWvmNNA/kFbGYYytcsDTRu
1AE8aZIh0Q2gYWeiJ77QfTMvLRjwFWWjqHFRE+gcI5yluKl+L+my7zI0WQp1rNyF
3Pp+jxM3vMK3eRAkCUc7/+2CZCvIs4NM7LaLH8tQYBImLkiaXuEkBS1xUdSmNfFh
NiNYlkOXyLNA8sF8pxyj+vWKlNyA2ALZwIauf0kcENjPTa4Doo/hZpMFE30JqGWx
3+/NXmYGoY2p8fycX30Vddh6Iri2867efSnzbAa9wzXjsRZZVcAvxzM8/jfk7XNn
+n+7LGLpmpUZMLmwdBSYTG2enVxhvSU8FoEJemaL0pMMJSRAteJ6cWNjehC09u2I
G/q+4+1GaRGxzPX03LUB29TWqdHILdRQAlNYeeDSO0zLW6iCNqJ3bb6hk6lOEEho
ieGfZOQxmlis+aUJRlEPLP6c+RR6LodGGodNoC7r/ziEOv/BNp5jAYyl1PevnU/5
5lVcMJ5Sk429nIH5zZUccjd1BbT0nPYcJm2v8RWKYL1l0K+986/pma2Kd5RYnICC
7VduGqJctdM3MTlppqUB/np+eYe6W7bCpOKCul9a6eqWnMB6uUtbuPnWiDLVyye7
9ICsW2VLJwtexKq3TKn71F/R4cRkbawapgyzfOlwk7CkXQD5mCxH412SzNDTASUJ
s2Z9MtWXh7g/mhbTmq+4Ove24JGlAltbtGUP7EjlAZ0mRYfQokrbcwvFUe3dXGWo
QWgUfGTX/W93/Pjmbzkqa2fnyUM8xQEn7Gyq7+KkpVUfL4F2hJOkCwW16pMyRf7v
rgEc/FH9WAZGDAGpNjXdkIf0mrPi9bTsMb8N9d+sLOAZ8VadQ6Kytqaf9/YJ98M1
5BT7azpgL9+kdnk+NXxaimsoYQAPF/eJGf8YdmYbHfrfd1HwPqk6jRxr4+CKlp+c
qribiNizRgzffzi1sv4iy75MDvfNq9rrkK3bVbalpYWWnM8RVoqAlUpXrJEBKa4Q
2Ty1sNrE1nL4STniBjVPqvRLXHgZ+6Z9ikPwkXiWBoP7xaxux8iWFkueyDuF9sGZ
g7iwrqFBaJLho58WvpiFb5qV12iLn0+V53yEMXmFHVMznVQvqyiaINC7y3b5CkAe
r5uqnIcLjE/TFabxJ7irmbpUIwGo7F+mebiwSRlDSV/5/8twanrEGkCpHKu0/SoQ
vQFQh6CIEKa0IEbk3ZUMaAp+Bl0D5le+FbhJL598c9PT13lKjX51DUEP9FaCfH9X
BgN4IIeLaRqTQmQPjwg7zsJ3ZRTmVCOxam34ajoHbgfX/WZjJqThekIPT+hTqSyl
ZJtU8LrXBz2J6tZ+GT3Ci6y4GMQfPVhnJGWWsA3l3b4eFwPPiNZQYiGMLISqpqAc
VebvhgvqXUhN2MKFAovqWroYzIjYOOWoEafql7tmYPdn9qaTpACSBan3akC/K7Lv
+np6AHmk6851iC30iCIZuY3/B+V6YXemJ9XrnvOTgbzij+Rr8T+gKJM+7zbikX5o
1r7bB11WbW8wiR6suZcB43x9zeuk+I7EuSv7fUpIh+cCdG7Dbd68SDafFNFGj3S+
uRHeGMEXrdbEDFYsgEV+u6RVSVLC02183hDVi7eaQROBJzUKXs5DPktBAlQ5BUNU
B2HRN2MpqDMoq0i+ySohmFMKF/OmmBDUKxAjIyGjy3F8D9O5XTFXTMMzJXS85iyI
Dzk+eC/C6FqCLA27rZGJg+IJRlAo40Wz41VbTzfFRYw4qRr3TZZ+rfGqzfsMkDtW
p+5ZIyeFWnWI8MJUrHzWrYu/R/XGqVV3DME3OQcf+9QOp3qpTJ7uHm0XjViPrdTH
17bSlpwlY+eulpswGvYZ3sayl+lngUG/Ixs77Xl5OZXn7UBdzwXUU7HuzrK7kqeu
7zaW9va5/B577rmnLFL/Yjxrknr+uCDM56RoNnqfM1MzjCuq/OoGrroib91nBI5A
uJM33AjSnl/0XQa80yOMrKEvND6NjywgEUo5TtStErdPjV4cLh5H3GsdmnfOFB6W
KoO45FCH9YZYceCA9nXF2w8KwOhh5phkCDi7AOgXpRwVicXaqILDISKPG6x5rsiT
ZfkIkKHQJRfZovBvV6rCEb+c1F9nu65vy2tFi2fiC3on+eOTPCtoG273e2h0gveV
P4TTtclXVW4+057OmJkjC5XMZ44nY7zCw9GJnNYHoPzBRESVETW9PLMTPMF1ZiA4
YQ/PNSsnUGZr/GuCA0lKDmJQdkKaz0Ief3phdrQdz5VyGJeKpVv+nHfIj5yxoIgu
kShnIfHsb0qrXtp464SDhpKLP3hlhzXMOT/009fW4Ne9aWFsF/IjVlZ3dP8phZcT
9g2/YMCD0HbBgDtsc7loXR83L2mr8hE1gp4LheG7YxJZxCf5RFke7XXhRvr9oWgY
EP/bJxzZba9YiUiUxug0UP3hq8efLeDb1HVUnJiZy/62q7c9OPNlwwSurx7n+qwE
ShhZUq8KQj6oF5rFRAehLPnO7cCE/uy870+ruPX9P+AFyqrUAI8qX1x4iMbHqhXH
AfhuCLwT77mPOd9lR4qtHxu/z88cDzj29t6u2lkwgqP4vLavVGSVZadD9ND6RQjU
cSO5xpEBFWlMTapkNfc8wNwFPLgsKemkzzk2FjgYz4a3baUExBg3BW81NRFBRvUq
doEDFG1Xe0wYMaghr2ne7ySnDeJqFP1otFfk+N5ktBexikN0w/YAtbJ6h5l2SpNE
nLtuXgb/EGRrELOP7Zg5N3Y3cQ1kGePoKIm3Owpr6HHho/Zu990t577atUVe41i7
gWXf5rOdfJk5UOiVQmzVqRmKwnbBo0VtrtSmXB/UUOysx5w8TaSIvc0jcynrkMrS
SpUgMnS3yFL79YDixFgvmL427uJHw/PXBM+AMp1C7/pJLG7V0HXFMyrWvswnp/yU
qaW7Q36qxvT6wxhIn339Y4wJw2oo8L6akGjRnbb07txfVJbG43KFuLTlN+RSJ0wx
BkGSh7NZxOYgNmCD1/h92hztRI3GZ/82h91ga79tlpn+ZingWGNf4BUk1ZB/E/tG
O/L7phtoGFdH6Ad4fUGVxILG7oaupkzisxSXic0kMbmusXoCRDC/Z/iolOohiEtN
MB0DGZysW3yYmD8CweXIOg0S8ercNlqOkhOCMUYpEBUk+AxfDCQitB4IHS5HkLi9
b6TUNeqplMT5lnTxkJhNlUlt6alxi7G5nu5HaDP3KujqOLOMMCTIlj0lbgel4mzF
VaC7ylwdAx66bgAY3ihzSfaXmYXl9t2BoVHBOS2o7wxzLdwNrg3RIS82RZo/kC/K
NF5jSUmPTiY9//GQA9tnOLrxXQoD9oWZC/MF1tfdpc5g+wP+h8/MHzPR4etfC6oa
C9FeWJY6NW4eoeq3UUVlQKUXX1z3Ptutbl32nL4CjsEFSjM1hXTRNEeUJVDnX92U
Z64RWTwDNapRuKb0D5/HOUtFl37shr8iSNF2OTkFRbN1yFhAXIpHQqDn5BeK7vOL
uViFIzX4qGO8T4s1Ep1AlIb1psBwYT7wodTkh5debPDHe2Q5+NxxM3jqeW2qsMrX
LzU1j08eBSOptgGYWRr71y1MRILyxWz6Gu+ldPxo4cHSddNSu55DOnR/gCFXQTVD
5JW6mjcGIY8ui/wCe07Y8aXTNGzENwOkLBu0zIQrgsPaYwRukrvH5Z2/6V6naoyq
HMh4/jVUCUTSx5xyEfgBdW4qNmxpV2cNhWKCAOLKtG1912+UoWVVCFQgtUP+0ryy
lr5V0HKdBlU3gfX3kO6hVpROLxA34nSfX0TAJZZN+XBec7yg2p/APd8DNOg1KJA+
HQzn19X3cax0o4aeVStnQBYDzaaG1Rpx9LcLQvpea7RSnnLjo4I2aCxlIzeeClfR
0BCUBJPc2/hRL1ncIztNbiYZMiO88SW6xruI4lu/kPyBeZ03y4bwt83/KbyJCaec
RFAcdxNxwGynJB5wV6UQThG8EQpv4emnE0Fn9yruaZO6fMUVhkSnm94WPCX2BuCx
i/kSyl89QMrv14b5qhRLWEcyd2HY5ZiUSZNvwFTsyymKfvuFczPcyxcWFW8c4Btg
McN4gZuPFFf7vP9IjgkTDhqmOI0hLMdrQv4fh+/9XbhKk6TnLnanff/eIh5NNefQ
hKFuJYyxiQf9uXh2EImx/xzHzWOPOWQh8JIAPx3yse5nEIHmjVmXSxQDL8LU4Sjh
9mJl/849ECPzORXNjgWAnJBD8e9yYgHov2sOoli0KWKFeMVQUKYyu5yKxqf+Aax2
L5Hv0yKwuIoMNnETYv+rlmuhPowneq5tYkKSEK7WgZEmf8foim4zFyTtXC168sBz
d2BVLhv21VW/ZRneeU0q3If84XdUshi0SB7H823hJn9eBRTuuNIa/DX0kovHTu85
i1wkYEqw9DfFM7j5qco29cbj/pri/d22S2e1Il13Y2qp0h+ANnVw2h3AG+Ylq3Ay
+RwK8zNxzg6Z+LC942rkSMMZZ996Rtv5bPTYQNeeHGqDZG3ZsnzXwvOP3zaOzogb
pE9m2i5BKFqdxCF3Q/skfkzsiBgDnzRQmMp0k/tfnR/5qh9kEckdJ+n05tDea7nJ
Xe9hZTrbVu9D5lnLb6BnHcl8XAOKJVIZYaVusMpcJ0JTpgeDGCfnwp+8CCcCkNuf
ghPBdPoDgP8PekSL4nB2qnddodMUOwKe6Gk++CON6jnJLw3tDvN1QebPOmazDPSz
rIHa1tl3vc1elVuOf46rbqC+eCpN9wV2hHq8crnHG9c3zLuqPFfmdBZjHvt+JOui
H4Vaxs0v0pdHo8rXzUF0YflideoeJ58CaoAzEeMjy5wz0WR9CNkwQvSePgGxQsIx
QQMcJZecOFDa3u6LvtcpYdbuXOWlvkQGApVIFQ/JUqKC/IX1ifehn0zB46YowUYr
lAakQ+Y3SiJh3uBvq0HvR0ASoZaZLXpTR/EEvC7XkFUwg0xb2TSJz5B/4Ilj/5B2
9G7PMSmFK+v91NOvydFfC3285Hbpx6OTJjKjxm0+STj9AHCLR7+IZMrT5zoiM63V
q1P7R/0pmkZr6xasg0TQK79jICT/JaouWi8JlGlxOJXInL0BEfEW/vUMCJoaSA6U
kYz/j4KxkRrJeotPptnOJjdZdoLW6ciGSVSFKfuq5uHREQS9q+KOOw0GMsrHf4Mi
qhSRwsCm7uOxxDaBWtV282fvZcXZweQNArQffLaUdhrQB/eo0pb72pZRgLNN++2R
aJ7v5Zz3eSOUMMx6FNatO+etoXsvmkmny4/rQEooElOvi5qaAOkvSb8GWDhYYgYJ
9U5FsoBI9wNZlN+5wxKhm0CllIzBvJRBak8tiWaXBCD/D5e4ppTaDVru0OVu77BB
3l+GFfBK73+iYr8n2pg8eJMA7yRv3dHVcysZsQMqPqcsaM6Tvm+VBxEuL+56g+sA
34YjO8dLppinh5rXb1fxUWAnOygNHRG2KWBGQVUV+0R55fefckoIT8mMbdXceMZf
iD1P5SzrK4/HsYW2bCRIxAMiCvErSCKYK8yHGWXza/wcCkXfJNc0w4lB+L+BqMGu
8fZt4g3hU3VLt+xcqdm1kF73mfmzvayEYaCWjbdxVk4yQrLJFf6vskCEs4/8R8Kt
grdRYFVdcEVTUAeq6POK4pykeXMZFIFMqytV+GiTKPISFESEj332JafiiM1Sr9QS
D1W3JthvrkkwRqBn4vZPWlD4SNWCUHcqzQig/P/ogATOiJ7ySmQ4j75Gkm+vlsQy
o11TYYYUfbxVBf99gNJ7VprQwPN1s0YYK6xafd/oq/7XuzG/5JZgj7L0fFvTvsv2
bnopJAQVItVYJArwpyC+4bOfhocXkFq521XVfLEaOSddryxC/Wxm4dMPDpcd8obe
cTrgv7G5u7OnbJghdxI6wq7oncIUazKC00h+c1S+t332M+6TPKDMLTkasY1cMnQ8
7uKvLJn+Huoz6e1VJLchWmdWdGPF+a4RCavzRWzPT0JnCzwL3aeFM6ReNtnpArFr
NcXe03a98wp59n9kf6bkxqstaWeGmRPeKzeDxiFqE8kv08Hl+Oy6d96t9BQDeMyR
5UpfxUNz1xMS8VmfTNSgCLlzlvB9uweqM2g3UbcOeka9ZCA0/jNuULyrj+6s2C5X
jEjS09kG5c4I7deWCsjXSxp/hbLk+St7V97aG2OGItSzYmtY5JWVmnIQqeLXve1e
UuRIN4dezv4RW/OyBunByZr+KBFaPg26YQSQ1n1EJk4X6PTUFg0MInobpkyXlpI1
OmyTV3sGnouzgQrlgqNby2+Pg5xxdldppZmpPGJpPDogN85eBjdtoctTg8Qc6VWZ
QLa24eVWkSd2Yy2WVDGuiAb4oYY3t13MciSalZAHtauqyr6kA9bK1BQfSZjy69/0
ofKCOwcNMhOqAyjHym6tH3D/BfiOxBkx+2iiyFrXzxEd5oMt8gJyGMkNOMUA7nTF
MubUUYldt8c3Rpx50nnyngMbaKxGJNSn0+gbb9BAzxn17dpzVhMV89gA4H3absz9
6eHJ1bAfuXEOrmzrd/NXv3rrsVDKZygO/S4UoKQM7AleBsNOd8XwyRySB2ewi2oy
dA6pBdB3DxfUoYgRpZvZRUhBW6alWATgAFGNoQtP8BMTu7RTH7ofTq9V0/VjsrPS
pe7q83jMC8NiKwMZkKqFn4VoCd2sirWfnIPZar8pBHcdFgDzeEtrhRYy+YNTyWek
V5tjHbV++owyH0dqrVZv0Dg+kNvKKxIpBTohVBRtw6z/A6doEiRVtHHNbUCftP5/
eD3l3fLq3arm8wBZV3aGTzP6Q+ldQ23oEkbI7zMU7+IVrerAl57HaXNBUhTPTCDc
up+OkrAxqyQr6OkuAgfeRAmGZ6ASeW2En4v/ieVHpnzZMJqSe9TIGNyrt9ScCrMm
+pyk0gMS5xQPWZCyVL4MGU+U2/BSEiNZEXUJrTuNLqwG9xDU+bLp89dDj5Yi5IV3
aeSVMLtPI2+s2Qsv/xWkhXbvPhvWVb+QO2tl0HrJOhSSbWawi6j9roPyYMj6fQaD
FZ1jIzIWSywMx+UKJ2CoJAmF0qWlxgxkZrCG0Nj+jGD+QstQs0wDuhdODbONZAQV
RtMu1ALw7qJIMQDUS8L6w55RVVVch7w5lH9LfmNposGLHxCqGxRlvIsrlyRwszox
DAPhsgbJDl1abbmStwOTy86UIs/Z3LPP0gwYHo1+InJdnfBZfwQc75TPF+3st3+s
PkNY920LiBGX4tD3JsIJcvYibHjzYMJwH0H02qpV7YjKdb7SSUNogBwLdhe3KQ0T
Pa/bXQgyPGcoGwiVoBt/bl3PYt2fFOMbw8E9n8+9k7eGSS1X5SHLF2M6eUtEbx9g
5UalAluypBC8NMN2aEqIhDC55MEG2s5tBjBIViS77WDE5qvzfATzUP77Ta3E6CEG
mmy9gvrXQlQLbRPBQKllG/hu1PY3Ur9pmLKoaNk6sgKuOvrp7LDd6bzCd8qyyj3x
2zvj6UQ8Dj12GrIZ3sSHoH5JdiND/Vibzxhrg9+LNSjLRcMZDIGK3zc712eeLtja
nGOeI2fKGS9lFBviwf6Tdp6vHpXTNv8ZWO+KYLvZ4yBVcsEGHNN6NFogIqL/yqXA
ItjjgwhqWUoBVjsCDDwevtUXYfUPfEqXvlIkyLQIJ6F4JYLdBMqXvnIOOxqPYaQm
PrjJUNMkN0osi0p+sBF/WrToG1KUZJIfzPzJ3O7b6I7iHBBYoHvNdrixmzjpQ3Dk
RUYvbpYTEzbheh27uwH+xhv1zrPKzU73AbcD5c+OMHbTv+0Mzf9SYql0ka379D10
2XY5rz9eLTBbN7AxwXOFBLu4eHGEMxd1LaG70+bzcGhMXnEk6gbfFtLxeExQPOtH
1lWDOeWaDhv980/Ea1G3pYmH3zYOgc195vWm5Mky3nh4UDOzJPdKHdt8CPlAnak2
8pZkDaWIKhC1E3mi/NgxpBnJcppl6ngJ6c3CXq+ewXQtLKNxfAjlY93TV7Hajy+s
J5Dv2UoEm85ITPkgpwxVYLRMAysf4QNfMoDql/5LTRw/A5L4OQEKq9qyQsxf+mN8
Q5L91Yi6+aJsiYV+10FVq2CPLOeZM0DN4zGCnxOPC6dzUkjdmNXlNWNqz/7vLRdR
8JbmwNqb6ODe+QADpBQyy2a8tT76xp8uqT5V2IVkF9orKZb0tpqLCzJvApPo01B2
crkD/T9xNneA0wzYO73Ev/J1Axp1BVyPdfs0ik7GCYFXMH2XbWuw9DUWUtN4IKYG
sptmH9k7lXaMg1UqQULMVgwbfnxq/luyHaGakcxUV4LX4W0gxd+2VIJv5XO96sYu
E6v1anvluql9JqZK0v+OUVYP162ePD92MlqfUaWFBZ9Zi6qeVqfC0xnKi+KBnMvB
gWkniYOMhaOkmNLhl1qVbNYtQYyMXs/4fpE6wJggJd1akhFo6UZ8fAQdeYrnNiN1
v1Du3bVkjfbwKdmSIFw63k38cfuKx0WW2594dN2VxC0MiowyCENKtXUxqVG9nmSA
JLvb6tAEf2HDtjUBuB5UEZOM6Ym6gOd0d2IXxHJxNh4tBjnt8IH8DEH9IltwHRyM
nN3RD1/hvPS2mlYvveT/vpfXXNY40eYZlG3ULnhmJi9ZyScENh8a7LZPlg95lhMa
r0x4ssQDbnaKH7LlbDj0tYXtlBa+fNPGxijotIxJNeLqvIQEbHkgKnY60frbUwBV
Fh1xZ2AqA63/8k8Zny67n8tJ2g9+3ZO7XXtTQwjGOG4MgwQXJpCjni/vnU8/zFXq
vdoezrG99CcERML57spU55jdrIzquQf+oHNmaO9EgKd+FkwNezsEYlqaOUTso0t4
D1sjb2wcmsz/RrnK3NgV89EXD4ws4qtkUY3f0MCpyjcQalAj5rWLP7uAzO0IN0g6
KXoo2DW6LrdgRH8dNCk/3ubWkfZVObIiyGUUkD6vquW47fnoLylLlxmC/m1EI7PA
5rK3LPTBNZIFbSxEY/s0mmqgFbHPKDlVL2nAj83/9VoDt1IeeJow+ig+Lky+SVaQ
g3gZFgKo6QpHmum164w4982JTA2SdWMX9mm0JlTQmf7lD4AFy6tjzUt6xXXZhbgx
dE8rY5Ec/xdu3V50isWhrKbNQpAIY+MWqvfB32h4YOmBBxTqod6uVWwDFWk3lPmj
MfkYR5q6EHugaNrLiEuadfn8cyb5uByoadV61QBAKjv5XBRqeWS8ZyX4yay9B9ru
NXGctSUEtSDbDO9DSqmaafyzO8rm0kzv8aVSp6Haj/Vmc3sa/O8NxPTaunI9qKjo
1xd5AYESBoQWttTgx1q0HDTzmGai+Oo2v8s9bauzcJGF7DIptxwsPtmYEXeua8p6
kTQ/0PYn6LPVLTSEbRZEzgotfkAXkKeGPM+zwziIWbODVRYZPhsdwB6ZPjn4GXBY
H1IwVbYLy5IPyeIvtbzIAPnwGlScD12u1h7rC5WwzwPtf6NempMsv2JhYCgsN5cl
2utIrI0wd7ezh6DPqaHr7aDkkjs+s8QyxUILPO2RJl1NPpm6zWvw20RVP4dX5xc0
9jQqtIYxgXed+f0l3Br8FEJoNjcRJWS2rWsQm6rcjMS3LgfvEltFoNwV1KJoCBO4
tAH5Vz2bEMdy1WTQMnL36zxMa+Dcrujoae1WYBRXQkpFEgm0f7cQuUg/p2Y93cZx
viw0W63aDNCRmNsAcwxhmda1AFO0CrnxGtaeMzX3addsyyVYlpmSod3tLZz2bDsN
CKO1UvzCdqlQ0668is2NcPjIjRxMaXOhDFopTuxy2jmBx6wMeAKRfWu8G4GAVsy3
xiTvGliZjcz5ONzhM+4ARDvrE8wMnUdjby6bcw+8v88KlD9eRTb2jHjnAGT0OOeB
GrZ0XeEAgbeZS33JZ17j7FHZHfXdVHz0yJOCjgS8EacZdfDppLnUoTS7WXktCpWe
0JHqAERsvL/8gWWdcPMA0DG9l98wRitahqOinjZAqxohzCF0tBrobKH++XhXnCHJ
kdAtv+/U6hkq778AFEtYCOY8JiW3WZoQZhNJhskdviYJ7VTAYFGjAThuQX9sw/Br
WpgeJCvp1YQ6rMoWE3+ap5XuKmVgzObRjZKGsiq27lqmBNatdjBuqLKNvrM/rcL5
giKq1znq9sDBiFSqcJG4uR8p23r9mWJOHXrotYivBkQ1faIiR7esVHb5CB3slLxH
dezE50+jw5/q069/f5nGEJf5oB9UCloUjRSQEzRVW0+XyqMhdECcpsTlGlQu5hTa
re0YulwciefF4Q5/J9k9gLzSigNG/ygbRYtXZhT0X+HyOPeNBYgot44GAOdVzo5S
nNWDZpt2xkw/dqXuJSIUMAHrxqU5kgpEYTgRN9OvjxBqP2oVefHAmiPbYccQ2S7R
pPu2CeTdZdRQcxfPjC0Q3znsT3lNgrvYdM86SN1+n3UNBm9LyMxVB5oyR8+H1W9e
GlwiylYQybBAlSngA/Ru2JeE97X6zMTTjVcZnHMUu2L4dFnf8yxALauNLeqKj2h1
vecJESf0XzC+A3X2Sasm+XQdIxuT+rkD2I7L08XSR8YVZoGEN77NUDBgmEznSbGa
LL7cfRmUdJwoa+MDQSxTJk0pDpWHrfQLZFPik9NRckMD8cVCj/vI3AVmWv4f3+lF
2+wE6JMFR2Ot+tklYMw9jaMzayKj5WaGt1jXQQflIg2TCN6Z6dCnf3ZWWE3lRaxJ
D7ygdt/PSKi9sVLLwyd1TbmoD4+yWvlCgtXBAsJLXuhRBeLkgbySABkCIfBu6iK7
/luT0Tpn7zz+PFchZHuj1qOYt0o8A8zYAXHmcjtdeZ+W6SJeO4fU2JYsxCJNxKH8
rC5L2yENIBavogqi+OeXyctTxQcUbSft+Y5BocDSMtvNaOO0iXf2YZyqiRnhP1aK
P1L1nT56FSrTBGgtmWEqPdWnzBSw2UqNkTFS10TNfk7KPCMl2Dg2SXfRZytmoCJr
PEmXWYiyDwQYv5ba9ub6sb4PzVzsD8WggQgS0Q2JOpdhQlcUXF61p0OADj9HoJa/
Dsn7ns1dOo132hww5maGgEwKGdbId/bRpzEF1QGMOiu5U/WZieMs97xX0Gb0wfup
7x+0BF8SN31i+8mhLIRwwIT6G06xEqb92N3Rtf3H4XLzDWtM7IaLEzd+h0+ivIRy
DdCowvD7WA7lAvh7SaP7SSU0HCL4GlcQjA7oe446B6fbkYAQF3LBY2c1AfthBcye
2vWvGOUKed/EiCBIMrL6o7fMeXs3iQaff0p/q8whKKAb40w8o1/b0bNnGjFkmVBM
8Bq/oPoo0NIDxXZbT9kSRoeJVcYUA//R6uZ0LNYnYeSY/9f/dcwsoEFKmcr55kZH
4b/aLVml0/P0iqebVIy6wKASFs9tytWmjCTYd0dsu3tTOG7s4zik7VU8wJAL34FJ
o2TIm15G0Tz118adiYxO5u6hNRt8Vpvp3YrjtkN0xVmc+5YdOYuwS57n4uQTTg6H
lDuW80YVIkrn7FAfCHoNu8YBCWy9Hcdp1M8dSkY6F01cUeIltEScDHCX+Ln9rcun
yK8oWQK983rGI2JIUlEADjBRjOcQPJ86cn32msL7CGvb/78Cl0KogjpQmyzECwBD
yhzw2eijHa355lS3ETcd9V0+L4+DlE76/kfKLKPvfV7NiCEQQhz712F1RImrmpDz
C+EpR/pTo4YQqNTgdGBW4n6GMJCtpy03pydAN00M+b+sfmfPQlkQc0wYA3c248Uf
pP07Oi5hv+RvtiBt9QtcMrBJe5guXES6Za0HIxKCDK+ir77px2cXhdLIIP2hi2HZ
MOkhL2a4notK599ATSkyRxCgYPyrsgmapYP57d5bwmHbMDCMuZgO1U62tS/gBvFT
8zPV2ie8uj2d9yIisR99HjrWeeqwZ5T5cwPKICYEEU/hrlsJRvHW1tqaOMs8VY2A
4UpYgpCiukxM/8spKrY6i7QQ0JX9j+m76W3GsHotZROgYpLTK8pzSEyHCc54UVTL
K/1Pl9TLr86Mw/GX0vgt62rB4z31YZCe2DmTW2xk+QOWdExSVPsvaUrmiq0mA5C9
KGHBwXvx59hxu2wFYqSyNbHD3/mB660GuOmqFIz20gqw8W6cnOqrrVx5OAI1JeTC
aEDcSc+i4PUk9wh5lWBHTFHqIajYsWa4UNdmwDDlebQef455cWOoLMGs6FKLzdgJ
d+N6JxhyTCqGt5lAjVusSc66z4KMseCZpzgN8QItN00yS0PZLEpQYDijHPfJyvIL
35AorBFELFfAFak0748bQETcHAltsJker5020Wf3dRgeR3pnSoxv1oaevFK9Wnqo
4NauioTpyBksVRX/IVq7hQRSoVWPPrK088svPkrzGQ6gFGBr/U3BWRvb4SyP9hO8
SzoJdld4G3RKRENziUL6+u2xBvHjCb3FhQPaz/6GMq0zP8GllWWB5S2a0IbScTnv
sm43jN1gpnTiIdJLTXEF2xrns3VkAfbGJe9+d02HOXP6ASgeW71VwkrsBcLKgDme
biru4K7AKRWCcT+dNOcbgx02ZWQM6FEiy/LBX3oJb5arxBMxFxlammb6uiVo22Kz
qvLRHtNO0cMpYJRfXWgjQgWEf2yvOdWOUpLkW7zY+datbT5kaiR/R4H6CfvVCnou
AN/Lqf6Ir+ksmszpT7kXjDhIVYSsGTT9BqUdW0dY7AIOGhBFjiUDXmq0LEyvzHZM
AsYeO7sShN1jNHsg6US7d0i67Lzf5oXmsbUqUsHXEIiH3jSn/HoWApD4/hzt5cDN
LarR3PZA0PkkHX17+Ww+OGbDt9btvbxp37emM/B8m0hQhFXtrD8FoZW4wyeHqS4X
kx13MPCaA3/I/KjXIx+Jd+VCmHZ0jJqmWgSoyIpAZxbmVMm+W5qvMjLQ+OcIbuIZ
XUucSp8QLE88A9xDiL8M4E75Iolcw77XiTtpqxrl+uo1+2ERh+1ak301KlTB+hPK
ujnwok+U1rNTA+doQwf4xq9VYvU5XuaPPpDeooWKWDrXo/qWyzKe0vNz6cuvmzC0
dfdGplrhyQ4VyOvHOfpURaWQQiFHNayIlKwqM/27vRC37Y/SDVmVAg0/DKR84TNU
niF14swKKYQM6ce++j9T0XL6c3ISm/nFP8QRLRunoMt/f/D9f9CKSnMYa5KvH/py
4qLeqhTqimLymfLThosbIZ7ZCnrV8GzmkMGkWr9Ou0QrLivlDC1pernC7k2icnC8
hD0H6d989v+nCmxJ7jHySJHRUhJTB3e7OXE1cfOV/MrXSa2uktd45E0Y5uNO3Po/
HObNW9oHkKzqQHT3oUwbmr9VTTqJRPyj3l6LIBtZ50PKeEWbnn9vrJqYF4kg3GRX
/XxpLe10lJRULzRnnmXuY8KfYr2x/ZLAv5aHR4W3dl0AtMNwB/y//n1Nb2R/CmF1
PSsJxGx6oq4/f7NL8iGp54HppNOTInVzkFRSBDSzViXeP5o2/uXW8yn8p8QcBEAT
gc9qgjBtrPMKtI4qu3Qnao21cF1QXnn5FepiHYOeKNwA8LJEE+MGHAM3fPdA+OlN
2KBcl9wFSBXs1snSr3qvekmidP3/Yfu981J6L3Ilgq2eBKQK386NY4DUHUhFybs+
tSzvfnGhNCf1nSdirQouRXz+1sdQeB6xKW15PKBYcuSQJIV4R/ou1fvBPFpCXsK7
gmuxReoieFVFxBxEsKN0KmAKi5hcAxQ0eNTKcjw3ncsC9v00ThLPCpIpV6qfyRZs
eGIOerB4ACezvQuribdrurBBihC41aRXc55Zq+7QHEVG9+kgFHx2lAnWwh0IhuQ3
R7eDrPdKp0MIZpVugqXk8fq19I9UObN2HYvOrndk2vxjTFZMrjS4APe9LOGOtolz
uHEC+nICdtSxKiInm5sq3mRc8H8mCt11/mEZUo4ZHPb/5WlCWKNPMmXVvYf/DaP1
6AbN+BIg7sVAy8XHGP1+4tTV1L0Sg99CKgA1V+vJllN+ipB0dYFLlrO/2cowdNyv
38gmBzC1qOj6o201bdA3h53OPGIhtPdg5i6+mB84TvJ183Oed2WnK7g1TOLBt6FI
0Na5tr69eJCjAJr+GqOVmmBe5S+bgmPkU/hRvctohW91lyiaP7dOKy3XoDL1cjwb
1E9McleLl4b9bugD5BJn/lqp7tTiN8W+aAfEMjVXVfSe1ckLcCXQ7LIyuS/TjsoT
6QhUVpznYcBEMFS91R572j7KOAVPNRvfMNi4cwu6adIjJDWVK2ZdbxgFmEmIIG3M
rAdIiRUg8J8DPB/40HpHKzlqFifZo7w4auxPDQvbjQYQfw4VzgPipfICc1B0svz4
JY8ZayIOjAbBORHGVqVvTS4XebyLlLRftBAmuZW9Sw5FIMJZ0x7jlUOJ+NoGCvHW
XkIsGrEOpyP8z2IPLlHv39kuv93OI49Uialx44DOshA51KIEhOyq5MphPUNNH4y1
6F1TJZTewBTrHBzGFoSETbKuYSTSEv8KntkLAZIBfIO/LDSSCEsEz10Pk2DEpKG+
Wzhj6397Cxn3aoCZ2rL/AWNTwqIwpBnRijkhaJIq9/qq639xXNdSHNAXYAQ02srL
F+LHq8CHTyXoH9ESHqU47Dy8jHzQFWjQPmIA+/glArImX14xS76/QcakL1BEw6lF
RWpOSVjSTfXNU8sXdzyT9xhrtA9NsCwO78djbIgn3InYlsZwsl3+WC5n+4vrvVcO
s0cBz18Wv7y+hbeJmmkt9U50NHAO+spTt7NQ5GUlSWZv1ybse44JYJYT8+h4+yim
NIcWgOMp6z6z1zT6WNMAAc6a5EINA4hUaINKC6h78+2UIiC6cbInh5Y8ULkcJmo+
YC7wy8fYBTAFWvxR7JaUFkP14sHouBKOt6OLXuSm9B0Z7T/9dE7Vjlm5k2hB0TSJ
2mFokH+2A6YhPfxreFheSsnHRgrQJawcZwJdEPP32sWN2gckwyuoTOw77DWBrcVa
rvG1MAGNOBlBsiSAhLr0nK4muyVJbbISbPsSCMuumscJe8ETH3/MFNu9CGoSU6sJ
k9v5atcdRxtFOg7/wESA4MlPFvp35zG53NqSX2GksXfZMCjdFQMR7NINs1MYCd7p
djdu+ojPiuei38KyBmFdWGk2rPXlLyZTATYLFgjGF51aEvso9Y9r9jMHFQfIKi7x
eQvor54UJmCG1WYyS+Qm4cpScN3bL+S60fzxD/lV1qznKRaH8pX693PaY6sQ0vVx
zQmyGVFFVkELTqI6bCUZdEIxpkO5qcupNqikpICrsmmWyQnyM13E/wNR8SHY4HQ9
FHckGatEcaGoOoKSODapepq0RhNBowD0HSYKFoXFYBWLlbk2zUnhjzVNXoyY55UA
5RHxdFepLOAo+0pFjV1uqEaiO0ewxFA67NtjkbxgJ7tZBDfCEOp+DR0RfO3pseI5
grhTXibgkwepmQuRg/M4uemvJlYh7KWoT/7eUYtMe2yj+PnRzWdAZziTZ3iDizrd
jsZqcKFv9IURZt6ophkmI9t5VLiUtZIRm7LnUAQ4AjaBZFsStNG8/XVZge9aRjWb
LEVf4bzlOkaCNsXd522Gc96o3RxH6LAJP4rsTa2rhAY0A0eZNfC8JTpIM5smsx2q
E+5kgs6VAho8+QA1Q8L0keN/1tijvBqLyVsT69cMD4XS5ausj1xJDTbLa5+ffGio
bDkak3TIofO8lRh1fyUySwR21d/4SrFjAUO+OeGMQAwvhr//GZiTHOFV8xovZhgp
43Kjbv2TkV/1Z8hQzfmAXP2AWP3u4Kuw7LYN6tx+gmA/Nwz+EkPGkn3j70QEa96o
3AWJYovX/xLTFQpiu748nPGxjgHSRMatm8jVLLFjbxVe81r4HctPCbD7whJeqwhS
AEq2xQqfpyfRy4YoiqsrvgS5gYMQrGvYAKsuEsQ0hY7lO94JCRLlOaPUPtRDMk13
8EDPgDS1SwOYqHRXrvkeM2//hTF9Hb4iCzQhxduCyJ34Y41NrEXKCFDq6ydNNwjF
l2KAMfHRxXzePSjKYo2wAQZdi6CW49/N6rkzszduTE1EsBnHKqhScaj4r9Q/nJEM
9HTapyqQjftTud8te75UerzsiFtmelMx8NNTpySvRfhkOweO8LYDdfe0NApKIwkc
U7KCaNj+JQV0gej+Z7w5QwqsoGfDyNXRTOdUxEFRBfiMssIqR8cMYRrHSWTzd9U+
f4qSF6GZPAbzzeokXIOJ8qHALtuHEvGJ8cIq4zn+UeFszgb266jdtW34h0NFshdP
+Z3MI+eXaTt52MDt+IpTzj2nATTTx7hj54NS0QYyv09yoNglkYaAEx4522hQT2Lz
16SCLFiAVqlsRSRnpiDgQa143c4mrGoY/8H77EwhrvyJ23vc4Fv59P74W/zcD/XL
yrOh543+gsaiz11l5XIi3HiP/hvooihzpOsMweGglUSGaPzzNHXc0Bddn3cUoTlO
Im8x+HASeHskHimIkPeR/W8YOxvhMP4CbtV7KD9F2XkMfU3AwdGxKOTWMZZTmrrN
douuqm7yMJz0zUAOOMyKfmJRhrCmZ6MgMcqnpqPjC6aBcMRx5OgBL3VOH6uetgYG
BPwYDfpPzx0W6NAVbW+0ZVfKoiP1AtfveOQeOamg1RHsPMzai7UXf4V3DMmFI3Sw
m8Dj8XTMP0rIoHKcrG2F9tXdQBcMVJ1pJr0dPvtHDAcvxPfJHj2WYR3uNQ99HDiT
54kk/eqTDGM8mu/9hi14Lcfr5NWdEw28BHILoNKQxDHeQvqSaO9LaOzMTflMexGi
2GIr6laIRDOJfzdxzGgM9hhlC1tdDMPjwHeyvtGXPtxG6M3CdUaRWyU2ngka1Tue
yI6NT0hpw765AvHmHhfzntbNKy4HiLIsdFQiRVz6lUHpfl6Z6jYwd8ka+egNL06H
aI55uOCMY8ysH7Ho9FArQRm+9fk5okMzAAmCWT/nume/VyNJgT0laoWfFTzGFBjJ
Hwo12ur0vJLL7dX1QOdO81sTW/2T8BC3iDdqhcmFqLSJb4rA8jnVJjGi0wkLg8uK
QylWRuNGHx4dqfHIiw1+vp8ZFJvklrbHHNQlcwzFqFydU5nFPiPQQHyinsI+8cNl
23xMu5mbhmwfbxgNSL1DaE1pZ7xEczl2+4RIamejhKCqX97svc6casta0sf/jH5o
/VEfBQ5hC6zXYtQiu7VX9bVzZFEPVPckC4WgeR0UwhxIVJ3sng5GMktJ7OuikEWG
psapqyTvD2ag3QzIN/OwJFtYoW8bOFCWBoB8m4I7vvssrC/1P2iSRjInPFUg4E3Z
t4vKxH2SXjarvFujrFUtGW8DPt1lBIZFv9rrEvPhyj2RbefOOvhjSW93AV8DWry0
OcT/6J+qepT882KXPKQ2O1PpRFde5BvimfrpEQ3hcc3ZrmmSWRZN4f904+A9+lnY
DQxhafYtM1ZcFHIWKx2P1n6lRqnE5tcr+9ArUZWhEpXQtTRdY/Y2ZjwCUcVW2/ra
k2g6v4j5HXOt0YJRtIanrEsW4BAHG6sdKhUmzo6/GvFmKKuV40s1ouaWcZU4czyj
kKMeVoCdfLCIIueKIsFz41S5Eko9JeWhm5jqsnDtyuf8l9kmmKbNEp4Q8m118cJm
AqHHs8at2rolh4n4vjfaSUa9U4yqdvnM5rxhPhSbTTpK5Afi/kyqS/zeC5b2cjFo
0qJQF9IKFi0Oe3w3YNXXmRpaduCKPywTA1YwGGZMSTB0BEAMseHJsyPD8lxt6P1G
JmICxNG5FEhjWyCeVo3lHXSEMbU510fEmivlGAt/nKDFCn0jJJTeq6ivQfQUKlhv
ePa3Q9JAmW1CbOyhx5uIpfGO3pPwT2tUrvPtWz0BlbAzn95UUZwGM2f2fkk4dlbB
hLBjytvJINJTf3R4t4hgkxHu320WH7y7yA2uWXszmIkdTgIdBSpbV0FESsc+fPW4
VbicuyzaQKPWybm7Kp4RGxj8ix020IYmW/sJz8YbvjIK4FFmX5asLMSjU19Isyv5
BVmGSfec4pGfbu6im9bF9dkeUtA+dkoQzjj9BoaeLOt7CrDvL7FvY88qoGv+20ad
stnZbQ0UjOZy6T0AMpbFruCdjzchlZl8nlWS9Ok1x5eWxXf9efC5kc8iLhrCB/Rm
sYKlDBewsh6C7H9sbWGjcTR5Jg4YwMfC43/PCc9MGMjrFIp5Y+rqWTVEa71/Bfp1
OI8HphTgNRRoB8diD2xmB7xfNnL3Tsxb4boCvqgZ+eJhSCm5fVNrDvLt7tzgKhKd
i5YU2+pHw86v0EWwjnWIkJOXd2l6aafXel0WBx+76Tms2lCjq3ew34JhjuTwLQi3
XeXFzP9/wmNqYCPDKZhBUv+zUd2MDKl0U9roEf0D/vt/0V27YjaQl8DyRTzT0rGL
jzLATWe0xX7Ug7iT2Pe/q8bKZFpfFidrIM+6x8yY0q/Pj60hbCZZWrR9REOKkJzf
YHyJEVajVMRWT7L4AoFcwzYRq5a/I0r679LUWEWl4ADvc5FahgLOTznhn2MEBwQR
U7cxd1kikxz4+igO06JU/Wn2PrRU+Yt4eODcVyZvIRMBrqtXpgd0C6acOjXN/Cr4
BM4MGL1kywLyg1AR7RqbV3TTLtFtY0pY2II1+5m0oXZoElrJy+QQNcQuPSvc04hg
dAUlND3T0+Joz6E0uas+6kIjc6wlRNM2nN8Y7/8+j6XbvCOMQgTYfK06AvyjJU7u
J6hkU3LT1xKYHMV8gT8kvlrqKxFTQ50iLI22685mW5UX7VLwvE6uEgLKwP1u9pdq
RcCujW77q7wN+JKqaKt1anLSBDwB3hiSi+NU2rHMvaT84J9603pu8L6a3Lg/3KCr
FKnipzo8omFpAzasxKbrXX9sLBDOGNxqMtUQIp+yI+z5fVUhYRyptJyFnUktkO5i
L0WHVfKszuxJVOodpoGYjk7LnfmnuG2kQgzsRLwLN1sHZTN7DCrXL93f8r4KJW7v
9qITECKFbFtXZX6K4xt3bNzBIZ6QFZYQ8Ld7+FOh0gHFpv29h8CWoeUcFKE+2BuV
C77EE06udb1M2+qvDbAqYe0yWjQebgyURE+40XkyYCa+bOYLxdIsNiM8tU+cXbE6
zHwZFxUp5xON/cetvorB0hE7iMGwah0BJH4FrFz52OuiPP9pmS3tS9vi+kHBC1m2
47Y98IdVKh7sutXn6jjUt/ZoM56F88nhC3T+iVS3aivKP+eb+zd8Pz3Z7lWGmjE6
gZyjsKIUe0qQnt1D4WOPri9PKSr7EElFzuK94NaDk0dY3PtEjmXWa3yyhB34q5eF
Zv1QAe9SQHugKoU9K7PBzPjYbh1LYMM4R0Ak++QXgp0QgsQ1ld/OhpAslUPUbyDl
9j4kOq48miG2Nw5NqmkEOkRMR+N5ngjEchgBRd6QA2cP9GOxgvbMJQyoQ50iOMVI
cdVmewfwhKs/Ubv3HL3UFlquN95GYaSXPvalBRmutjpZERVNYTZitI7eGz+d552i
pbUmNlKwL9M/JHSb2Kt748K9XAkiE0gNECPZ7MTuh3UROGW6GgneHHcs2Bs/X6Yq
yXELYYOHMJeEn6Jz2pQxShpje+lhHDhxBbFDh6VTGjheoGCb6j9j2gz7UkpTbxGa
EeMuPD/kFpHlmcA6kaEaknKnzltmC6L/shPgBJffck2sM1QenOGba78DshVIdg8K
CHLOXvgp7R1nxle7iGzbewd5u2jPnO/57V9vnHB3yKrH+eKZMfXNbGjIglOugP0k
SqIhQ3mtPDHXFi9D6rOm4Oa5KqnJ768euUK4L5p+nkvQ6KJ0AXUDuipB+buK2Udo
8Eshoj3Dwl2EYU5cQc/3+fbCTD/UY/YrggQ+wJWxkXlCEjD+VS7zpOVs5l+lApXL
t3bWq3Kj4I3VRci4573w731mnnuOJUKJrXocGY5KGQVtOhM0k3IhAlmjPW3JRWXd
twg3+0iLNH+fwoSRCu/0gV6VbqVFvX0LtTMXNxAfCDs8jO+WhgyZNLly0DDTGRZ8
kMhtkvixLZPxIzRKfdzulQupRHVg5HxGyEnvt3c8on99OMeiNlqv8DysS4i3mr/b
Q52LTDiau3wGHOcNnQ1bpDIct/pdUO8FHnNYeq/fCaYXxg5TPU00OISn0JlezQWY
MpUhQoDAB46yJQHE4mgDlsyvfjj4yj6D0JpG8AZvASMZ7ieIvUux2oXsReqTt8JC
jbx3FqCpWI8ZHoPNmgJmd1zVCVyJBqcXL1IgHtztkJGoZDRX143Ls8YyWtwJb+Un
egrdc4EK4pqcrTtstROrO1keMU+1zSp/MWg5qLfeLLEbn2XCfY+pplxwVHOHBG5D
S9eXY+8d6xxzayl+BypQea9OaebyTR0/zYkC6iyU0fX3L9Z8SXeM1yYtab8oOBKG
nlrQJNHmjMFY955J7KN+uN6KweY2U1oVe2bloRkkCVQ5BI8HyGV8fwZDgHeZNusP
eY10HNzN0UxvPbxOd2gWNumu02EveKRt+rnr3FTCiqM4c40GkE539/Dw0jqLQuxq
QPKvpszo8OjSp4q/xcb/AGicCn1hLrcbUGEqqOL8O9ACXm8rjc9GCql56qI4eiHx
Z7O6ZoqbBOMmfsuv3qJaEatAT7H6j6pq0c+yMQKxtDylyo0KhQEhySlapHarCqtC
fZKoe4jn0l4VYkBq71mH2g==
`pragma protect end_protected
