// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:28 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WiwC8zqv47sD+VolxMWpKqdAjbJB+tTwhFy8dfB9pLpiTXDcxPnsZOko8Ylcp1DB
4E8+lQUdHW21DAYyyRk1KsIQJxu38xUn6w+S+E+fC0dknVhouRLbS8tSU4PkK7tX
TnO+H7mUZMrstOmpy9AWT5D9ji4zoJXvS82OqzHMLRU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26032)
IPnmLzvJs52dJK4u+lG+QRgyrOaJns4q4Wps361UX0vi2eoXC0DvZ2nnTMX4StC5
2+1CSDJ9IWorTTlmVpafDbfqjtI0tbholYsCpTPSBgNa4b9HkHxARck0I9Z+Ko8B
BNEJDIXEkzRvIFSOReDInRwGoUJvjf/UnDDllkCmCx0mOvHkKkqfiWDT1l4/4I/V
sTMzaPi7JHzgSRPDYsCXGhtXYU4CVX+Wy6v3SlIgvo14vO/nO6jXi7RmmmOZ5jLI
jql/2VmLwV27jvj+aMIHpu+NNHrvfKPMh0xcZK5uQMSPOGNybD2Y/+3YsdyIsB4S
JtpF0ZOY7MA7qIb/vhg9QWPltgW0aNTG7BpS/TOvjB9CzNUdAD/PRbpiquhSmcpC
pc9w2uBrbDJUY6hNsaccxnNcbfZsQoJAHdUCr80d1Y8L/Oi79brVMJmW+FMVykiX
xzzEk8HQCQVEXjCC8QTdBRtLmrWqQvmmbajYYQUa3K1SciNrq2YpsDMMe4t3cxus
ibxqJh5mJWHKLKd+Y4BcWL8A5ru19ApK2pCP5SYQJ5a4uxDYDlS+GM8+Qk3Bx6Bu
8Xy5sfpU/3m9clSXuTdA0t6Jq4DSkm8TxbZSamf8K9dAJAXDWYGqpNR7kgg+3kYC
41hLYuxkSOUBJmgveBVrVdEI5z+YPOP22Jfks4PGG7jcOYIss5QOLfRA1hQ9AA/F
rx4EohNtIHSEQzR+GDOq//alNqmSA060ShXuK8YuQ/XSIlv5dX/LBEr1Nk5ajxe3
7zc1OwU6axGJ2Sm/MTeF2xTI37+ZRs+bffiUlCZGrrBmSnUl06gAxuq1c2p6o/UI
W6M1Jg4+UYyOr6Cp6vCqFAUO2S1OqNa7CRK6gAuu8U8M+7IFxul5LoZMk0Fg+qY+
RSlYOIXDxROa2FJCom2cnYVI7pmj2lcXGEI/UUHTEd6y2v5fEzhw06Ns+uoWwY1e
essUG414HUA+y5c18X4DrLz1NjjX37LtEcpJK8AY4yLQcuKXSywaoMkbJV5uTuzf
d+F+WOa8oqELgBRZG2fIvDnFPHRwGGtxXEkzOw4IEjJMhN14FM5uVbcbOEK0ghwi
9QAHwIq3/isRUW3EX0OejLmI88wbLwxzVuaohXZGjRjmMp0JCI5Hni1QDxrTE5iw
E3aHWCJkVX0WHz52EgHx/zBOVF980NiKBrRkTP9RnXRbXWA6wzgdwkxmp/rpXYZY
GqBnbHAmLkhDVGuIxULP0KcjFdgNpPCmWGxXlpDNZfzNki4EZ1zsr/SD0tawTTm7
HqAzhbPkYXWt6UrgKzcgR83O9pxUK7ujKPwiDABc2XNwEtSkoU46celft0ou0FAO
Yjlw89L9eGZV5XzK/a9fwJcQmCdpJioUciUjzBWkk8gTHSwH9c+UYwdAGmn3g6RQ
4DUlnluH3HDJG63RvdKHU457ES9xHOwAOKoI6NQSirUrCbgIseEGCPd6bdgCJpXv
uR15W4Pss/i549MPP/QW2mnYS82TWauu4no+6WBuMqF84wLTNLthRyLUF7PaHtB6
dtsmrVpBfi6HJaKO3oyTiyomjq/5CatbhNq9bB0da8vrfct7hevvEhhPfUzpJFft
OmY7YuePs/khOkXj0YnYkzVpYiQzRhF48Db/39iUA318Hg9KEM/kGzxIlIMUDcf1
WUgyq8xUvdPwLVTco3tZQWGZoIPnmeFy0cRrWzVwgJ2FtP2Bhyskd2pzDPGdNO6v
cb/af8QlKdmU/dpFaoeKQSeIGc2rlT1nZKatJJSll4A1Hibpq2US3dsXzoHJUrrQ
KHvD7qWQLgFDgfPIx9krEZOwZax9GjTO01RySjMtQ2FRxHsZWRjzz664PfIv8gnA
iQUeNZx7hAceID6DJrW1yqVMjDER8NJUDBCQjdEnnwUo7WOyyZrU3yefQqCDPCnh
oX5J6z+d+19YhaUh0YLWSWuR9NFQvymaIoVPOni6U4dk22UUbKw4fHBtwQhqxt4i
N+nHXxzNLaNVs9jMRPWiA9iN84Db69V/vYpR/GdxSYG2izouHuu18ZfBZrKcoolW
B4cowBpIeMkKJyIPOCKp/70oqxkccpVGU3GDpOf9bHrtx0Sdk2QNZwWGXJV2uTcO
4kgvcUGb8QItKyBdpR1C50HYg99hsIIreJsCzo27sPgHBLDo34ozmDuiPBHsqvcf
sWsx31DMvWMcUSTEEtBHIhFcC9UsZgl5qip0dUKrmgjWtTQlHLGiYSORshoVyLnY
c2TtCtZZgidyfwEFFND+p2bYM8FqbOPwJH1QMluhpeNMVYXFt5nHhCIHG2+t/J06
tZixIOgTjAo7RtMiaMVgdqj+c2XFZ7pCrnOUO+IPYv4DHm9cYNL/kVrPyUX7b3Uj
vFD54N4kN+iWcg72s7VHTySteglLYpK0NqEQPaavSo7lBc8RS/Pcn9H/GEPkKI1u
gZrVuaMFAt+FZRcWj4e7ur1LG8oLsnN0hjgc0ShhfYSpd7UNidbay8mPcAsKCyJE
U/BzxkMIcgfauDGwHR/BUYtqNujtV9886/MQGUyQk+2MtHKrBC0SGIDJL/HDYbVS
jCNuoidUlpd6IziDDfkzRGy41QCAG/Kw8ShVDI4YkOxjOj2Z5L+DX5mwNvmmOgEQ
ZPDiGIjiRUAfnujhlzm+nOgyj1QX8IXKpFHs7qD1+Ashh7W4/Ng6WkfJs18F/0jZ
mG8BOgMSOWrwiKWffSTQF/d5bQlQ/9nh5/Z+YAa4XHbGVclF4YEUFNd6V61We2Gm
WB1/RV3JJlWimhs8vuxISwPqrgrGPyNAn/wPzxmwOYdAFhpl8cN2//5xcqlBa0D1
eiwO5S/f6BfsSsgfdBtQIWaeZ56W0NKq/ldS/F2RXIHFHWc1XMMd/2/kzxnO/gZg
w6nI3l9X4VdCKggTGKR4UKqI/KP2imKP15doog1XgngwXE5piV/kq36t70NHLtFD
VpKiPvBs/vNvTl9Dys6Q9zF7MBJOXXx/R3YHXJ5o8JcLWUvvSGzKn4eztSFHsQ/l
bGuTUhABml3Jf1PakhiDSwrayeHXDMy4VGU0fHf7F9xRI8tT0le++/qpph0J3xGm
IZqZxJwoVBxL3v5/dcNyaZG9mknNUfyO3BgJsKt4j9iIEiMPBwZqNr7bc3yH3LkU
Cdvz5W1k0Yx6X9gdbAAtpRIZK+yj3ZdLdPH2jgmeKJvyCIlUp9sezgoo4ER/6d2E
qE3hS/Ssv77Xx4tWPErBBCyYjVv7aCgj1uErarm8q7OeoudypIyj9Ri7J+NsShiZ
6e6nZslQnAk76HSXBDxwZxtJ9l7A8vdR+GwNO08ni4cgplbz8CVSksWw++L0FLaN
snlGP5beUM8Hgb4kVkfl1pMGJ/psWwuydbvOc5Z+iSm2RkqeR6Zbs3I8n+Jncok0
O/BXsFVU81BwMVyR/1bdTD+kX2mreuDrn64aBJK35gPh1Rj5LSYSwVzFuDDW5Hl1
IJJ+NSVa1M8FXEIvPlR3BB+bXb87A4rWHzD4r/vcbaJFD26AxpXoaA6s3ry83yPR
qVSRsAU7WVDylgfww5dsTiWXp/pWzQCNtAMIheipU+wwVR0TtVK/ftelNjlJbLBG
T1MtmC4/2uv1A2VWKkoyA+prtTv/p1HKIlVgaf5xiAbyqRW3XHfoiu2XnOdWaq+M
Kz8NnlsVAUBVydV8z77pxTsnt91Ek0pchudZbbyXkz9URpjcRKVQSf6ma6wBOCAL
m8h2xjCV8tr0xkf61CDwM+kxBP/L2g0dc02NSFsF2jXHT25mb6TCQTpGaWHLRziY
Mas8gXlC0rln9tVFbM3J0H2/GJYWYB37bEzJcX5ZJnr9Bc3l0gNCPGsMIPhXLgO+
4/KPHXKPcGnHBFHiPNy9hpJpA1hRNd+xHi6NXcF5DMsfz/e7O8kglI6ozYUk5AMW
rkhPm2MCEpk9QiMZ1AyhnG2tgXkX22dWUcpwTkMIrmnWofQuPapk4KTGRXvAiYQQ
0B8cQ8ohcr2sOqZizbBBOlU7i/4MioDAL9bNrkxypyeDQi9ZJ66dBTQX7Uc0W0Ut
jGdmhyUfGYIeNtiH/IVf5tZeyJJ3JJmes7ggj9oAkhmb0WmLGg9L2qnEKNZO/Q71
PBpPiG9qqy+hbRLjgzyiif+EwBLm1CP5NYfrmuJSwJcl3BX7PclKeT6WDFcggR7W
GsKsffPWLgu5IY2+WzpvCOYj+bzMUJeCTEM8z6VDlIXgxPUAOqKLwQ2JX9FsKzNb
BefWeQ5TiurTzaZEi2PLNrbf30UdE5mlyT1r43/tziNm6K7w5qRAyIiQupw4eVVZ
UYkVzF9dogwSGoLt8mIeRlkCBYkp+TARIXw5r9bgkBegXfm5h8UroUHvaMbiKbnK
+vgO2plpeQAFcRunwOMvLGLRdXvjcdgK/d6Gzoy5+ezFfaAGP8jYT9W2YJOD6zd4
a/rH9AunyGv2SYUdqTCAXpwn6G+B4LRWOK0a/JZuojzyG0zDhp+qgm2sN2ojZSH/
bFFOFgKO4iGyC2BPjZxCurspU7E3VPqaE/Eoc4wX6m5xSw6Dbe1CoTEHSo3cb7ff
xLIzlosbzNjcqj72f80bHpeZqEJTuNwv37Gq6OG9lCFUX06nfnwOHVjhJylvAK3e
2HdxWKpK6dIez3X5QDULG1MN3tq5EkSQtjuIqbnRBw3RLeGJT0KIIsU+C+s6E2My
dDrRldcYNHGbNkjjCb985ZTio48oePus/GUuTsQtKNru+2EnHX7BmIcdx9yXR9Re
0ZZB731zXTmaqxIjlCCBoL+CTr40t8zC6Jp6Mh7hAQnzpQsdhyqTZ6eSy51toBAb
WtXzkKxrXkSwfSp8RL6qj7A25HKdTj02XlMDBS54G9vmqKdrIaZALxryT7UjwwNe
goBCcK5ky0gvYZ9GSrZcdVjlMN5GwvpeoNSBwumwpM8fteH6SVk7khec+IqkIWFK
OtGKxGbgRzO/hF8OdDh4uadG2BY4bHntG7dX3FMCbA02Qx/SgouQo/jsUjV+oEq/
Hrp5XMHGAFhLvt9jwe29nzC0QQmjcKQgwiHu9eT48weNntm+uxF6uM+as/Ov4smd
zWOxTh4KZUZ4nulVjRXqvhu03g4UG0MDXyHluvT81ckgY5YanR22gqNHMcRr3np2
5fmrPc6LUqG6R700zGrWMsUCh/jVuyWSaxMYsh1TkP7P8tkUn70rBSH1WBnG7N4+
imp8P8nR7G/oxBV6LuO70SwQVubfPr9HUCIqpiF16rUImMVgkyt24FCBnBd6Dckn
u6QCtLd5lGzyzr9ZLGMd4m5bpTlrMPz7X5zTmEjwrwDe3y4HTeNBfdCTma9bfIeE
YdlzQe3eElK4ATIV2Wb1kAGSLAiVHNVuTTnqqiadDQEx0ynfvm5BOcJKf2GY4C4S
PG//SxSnnbgaFAx29FwOlaVcarKNAm4ltYX/Z0AHhA2xaA8+ogAnVGGafJdfmcwv
BrP3LKmeO3xhU1fkIAoxBv8TKkpf3SaNPOwSJk9zsdx9XpLgff4sguH+V+Es1wXT
VXVBns8Tjs/QsYciUOEmwt5OU1pbI0NfezrwVrlucsV0rVNIy4O66Tagy+gWgJOh
cesx13Sb4qMXK/sb6i36SaHerDOf7jbCBIqRAg+54fEFVCAFmm6ZLRYlRajb4iIZ
NnwA1NkpOjyuYN/XOR57tlwK19q9X0+dpzFsbIT8IiWOFv5ChXHmAvt3scoXHyiM
7HMxtTXwm9jMubNbGJHNJbCBpPutPhaJ7lP+Ej0X8zwzrp5BmF286e8dKg1dYHAH
Ve0t5iy4f0e8iLu8ilJWQ8/3CI0B1qHirshcUDKmh4lyxGkOLtFqZfmN7fNbTW4z
8Z6272JO3X81LXLR8yeqX60EkFa7F8DR3wnfJLCPtDqkWlYn+lpc6TW7eBCg4VnE
CvpPD86MfGSAnqFvHiP6B+O1WYNadmzVFFKaiOiPUqOoRvthoXWa6gpaXau4CVXF
OIQM8NKpcxh1W+RjW/i85JLcqyWsKH4rYQ5ykLv+dzIATgcafqX9D8z1jGQIJbS1
tmHadahbcT8hTWRgOsXxoevaImxRKW1IOp3Tc1O9C455uY5beIEvCbKKQl6h5/Jk
OHhYq3j3dml0crKxbJRI84lUTPgltZVvmZh3Z3QmQqChpmT3EcyYt9M/iiBdiR6L
YbaVvckvASVUMjWQFYpz/1eO3fC1RaK71lFMmfeCPqQ/4mV/z90XtTbIP0bakZA9
px37JTVkQaIMInIqoxzuchrA8zyxJKILC3T7RHOsoCyqF2jvJOJbbySxT+vqR8S7
AkvBdXdiya8azSPMRoyGdR1aGDnz1T8Hgw2gwvdVCQXVXK/WvLjUplsVL0QHE5tv
cmfqbUmTmKXszhmpmaQX06LL/5gk0uJWJO4QPQaOU/r+PMrX9VFY/NTHFdTh1QtZ
D6gx4jRXiSsExqe1kEkBzueswGs/AKt9MnUqLhQajvw5UDmocqIGsozNNIfsROet
LaCf/78IDV3IQu2pvW0rrWH1z1aX/Ulvir0Hs8DNbidrBGBcfiwulL6NnJ8qs4Ry
5Ggs25kWrrKyTFu7eKfXi3TJBCsgAReB2HXc8JLcoDmfojM9DyDULN0s7cVika8k
Kt7JAKThg+Qj97lXHrnRS/8XoLJfi4UImtFxfdTUs0ylS0kyNAgMCRwcHqJ12O5z
HtMy5duHUeUnLbKOk+e5PjboYwRzhkbe6kWZdJ8ggPpu/A/fGloVwBRfKdVqmdYD
8wdBNOWGW8mXwE0czl31vIehmIh4NJPEidtSjRLCEquXJ1oZRP1pcWFeW6E6ojEv
RG/lhcggEBHGpV6m0pdmxbqEppvnK/s8OB32WxiYKr8DGMj0ygBEsqlFDFl/E1Fg
taPOoMKPQgvIMkHoY3ELwf4elZsjYMKWQivhNgarnyjo/1d1BXNQSuYLeAkdmoOy
BARFKsvBhAVa1vKz/GwuTgYoMIey9TfEJHRWXRypgoUS6Fh2yzcsN6XebgcocDZ7
Laem+cjyPuU3BxmAmov2qbuBM6LyH4IEV7NNGN9qlFT6wpA2IKw/3i5uoFheKOdw
piLMPcXImC9w/FhwYjcyprFc6B1Tbak+viWt3tkJ4q5U4l6V7bQMq1nDVKU53nRO
KZLU6WtYCporoE/c0cJgzUWC69dtoE8I9lvc7o9+RPdXYAfiQNeNrc7lmxPiaY92
bqjThATMPQKk1cyfdI5DzuzBP/bDY2g7CJE0LRdJL1cRo2y+s4Cm6/jfOFPfAIhU
PuT3YfbXZNRQQXKHBXtHy9lOmD2hG5gF8Q2LyEx/5WZ1/qL5uErYEodb4IGPu/eX
3ZxFP0vrFUnSoA4Bm4L7BBo8LEXnYG317Mqp0h6S5d3dCydEBs0vgFZCVaSkUMy+
LFqjefT+13IWntaY+1DKXPeLjlb4EE9DPS9w4CA71Ik/qBVLGV8rvQJbpq4gNGFv
JXYh3uZPcLK9OGSGJTaMOIdta8BKgR44pBF//VJZ11h214oUHM/hOj6EvjBjbvxg
f3gRvhNxSCgJNM7H+T9q+rn/cWB7FmLTaAZW+hELzxVIdIhupI7QqqFStka1dm5J
O/t5+SN0BvkbZCA5w0EOIuP7T1KUJj789OFP8Af+U3OSPFHPbkFFUTluCUcVVLjP
jb45cVtB4hZTKfbnd624cQ3mr6F5KcYlGUYLippz3cV6rgNcqjoMIJJ+zwUTCWuE
+/wdIqDZHOIfNJaIU8YTy/bmq4n0nnifZDPCmB5lUHsAmsPfQlCAHQxCV1jD+NCO
mZgFhKnY7+JCLd2Sxy1Es4T66+qA7L/khDWQg8o3w7W6adPLMKkZXpZv5ibHDUwm
K8sl44LngLaN1oACWYE2gWLzF3q/lUOhdM5wutU3FpCVbcxEmHWKp7n6f/QtDThM
ffwLQ3AFBnV8ldrsR5wZxvtNMzt+xbDKxWSLHteP8FO1c2KbxS/k/P7Ppg0nWyZj
t2OdVqEqye5HB1qmk7h/RD9O9gLRmi9n/a1w4nh1v6vMv8phfDIt9CGKYbpyFokV
8H2pAitoT1GGs9vOQ1WUBl16OfeRzpGEZRFcyb90r8jgcjg0p4Nn8KvaYtZ0RDZd
PsfowneD4U33QEtcehvrkq+XKqnoEzh7jaRutm54IiLNylApf82wyCOQnb8ekYbe
11ER06qIg2xJeEmLLe/D/IdmzGkJiFSlLhG15vEKkc8/iQcbfFwlkkAwTIK8ioDQ
7KZDjRZz4eT/kWhVsUf2mTf2hLwjB3oRsz4uCztvVW7OIQRQwt9Onj5VQYPZ5Kha
kKIUmjFIjV+7TvDeDxcfkoCoh74Mp39MSNWPNS2vY4qrA+UZ+wfry7QWnIGgVxXs
JS9CrQ3fWyNpCQIJxqwjMZ0G7PQiR7xp7SL1xWfD9j8BzrmzH57PrnVmAIH/vl9B
sU9rss1YZuOfAP+TGfommje4D8CD6phllHPaT/G51vVMTho6nUeUKW4SI61nEhZE
omSdWZlh/wKh8p+35ubpEJUqUmH+M1k4kmoSzTwgo3L7hoQ1M60+bpP3t9K2xje+
Fnx1euy9m4lEGpT5WB+r/Lq2ZhFW6tv53etQYbOq661uLMflLOtrJeIEln1bqGwY
95A/o34QSXCK7c/hnkYmIA9iwlrJm0XU6pDiN0uAyaIOaRF9yHou4X7/R5O3yt51
QCCidhtcHwGcLWH4LNp4dgRi7TWzp7osQ26rz/0SatZTelYndQgtl/RFfmqwH8Gy
G2as1eTzId0IY16f1Xv8rZORmGb1LNq3SWNElDq30/8EUEiR6jygtnFYxTWL22M3
zI15Rpwu4+BEabE7eVi0SPrtdRjMyM3zz/juWVfBYSJB0RXsEcaSWJLGb7FRjc5o
IlVtH3nAxBrLQXhWw10JdTLuGM8+dVy03l86NgGkTqgSmfuH17HqTWSqzlwc1npo
q1G6acjeh2IVjDVSxNGfmrYl6zrNJ2TjysdF3Xna/CKWMuUNVkfPGkZ0P4Weu/pl
kqlKxxBNpwKqoHcBRSKVmYctJcsJmpMLISsU/4RFj6S9l7tRUsUgKwV2HzXY7V9B
VnuM1BjGstbg/fAIPxS3C5mzlKWf6GiFvD6ND+q/ydfTy8GcVp9ytCgHZGQZaVhp
FAYfQLKxdrQ7Qm38SVJSLCVx6jI9dZFx1GV6C0TBLPl1SP3tyAA7QMViWedxBddF
TSrh1/Y3ErQd5WOT3SV1+7dA3cZj3mHRhcncu8DhjQ5ql0GpQFHRSPPEybtefCGe
UMqTU6uYS9R1Z9d7j51kaVdy6Cw6KMrJaZQAPrxMFZ3Rp7Ru+P68dLwjyGC+zUb5
DGbKcvAyjJtQ114YAgNq99xO4zwjkguc+IDvx6YlBkok7qiLcLNYUEh7b1MmYkWM
YsRLCZdifBmdDfj+WznN8mLwuBB4CEoIpQo27seOzht8XjzSAkaIC4/zxCT2tXM6
NWCcBOwUqTvF9CrUW2Ul9RkdRMji7KuaUx3UI/9E6Fd8CulyeI3mbCdRLs7PKQNF
UuySflitnEvRG8yAsamYGltv7cf5VapCtkuz0vCZYHd9sUB/T7b/4tC9RrjdfQZu
tl6AhS9j9prqT30O6x16sdHBLWSlO1ntqdZx8GnsQ+ugv4BBKPfHXA+le2Yw/4/o
7MtH9ewecRISikwpv2f21ABWZJoStugfPv62FtNUxmymBP5NV8jplN1w6NH2MxgH
xQ89z6a93gl4vXY+C5BTUW1k4sJm4o0Fo4HCQ8SZ5z9iABtx3YffDz+qe9FAGmu/
nSca1b2a1nuPPap/e0UXANOtjagztYOypQemSXj0obd/EHntCUSCglvjctvQFgh+
pAnzkKW5mi3VebKmLOS4ySmt2vOMCQPRTA/jD0Vom24tFrDc3RW62AnO/n/HtDQp
ZPN+GwI/KvmRHpOJ50oU5OVy4Vp4bxiToPv5jIILV2+a1iUDuEVkFMUNFXu68IeZ
CpCGL6+UnnJzH6F503Uyx8BjECIjkRfY/rcIRI1lwm+fJh1NpkrMdTWI4fZuxP7o
YBXA47JcL3k25UM17hhsfiCIAoM3xsYU/YF3KwWfzfw4ZyQpOREuLOgBQEltvdMB
yG2MwJiJV8BHc8ZcNVV+Bo2v+DVmfHH0VwAS0zzdVQKug3rPaS65Hig5eEE2nzgN
bK4wXe/fMVTg9ghzNC1De27c1uBRET7Jt0dV/FkFAOGfqZgAIBF/2x5xZ+DpTnsf
2Co/NU7JMoJ1NPE92ryM45crqQUvL3cQwycrBAnkCDPertX3ULNy29NpNdClQk94
tXrqTyivCs5wpyJJkPNAMxZxqRiEuwbyR+tzKqC7lobbL7GqOI3bO6t3JyZJLk+1
5TLfbU0cE9OeEWygEqIZy4GQRRgk02hhHP6Ux2xQ2kR9z7eduN4KUdlqUfhJGGOi
VJnncu0wAZpuaSeHtl24+STyGkBN+Dljefr4aWAm19Bc+51BuEdAuIbQsX0lDMBO
+FlEtqSv7l7TphDrc2Sp757FlH0zG7nrHI4Cp8dbdIpvNTorYtBJNK43r1QeUdOn
pzGMQNhlS9KFbn50RpG86/JwomZqFmFa0hsjwIv/D07EWFM5Of5Y5yLOhSAjeJwG
Q/77dnEvESAs59fmvgNaWL+lVDjUBJwTkDUbRm+c07+skIJ/bZvn+r+HXpKMmfz8
RQZbSdArhRZSrFmDdYnA0PpZXBGPFh5oSamaBytOFq9DthTuBmuQ7xRfsaW/PdZQ
zr0sGeihW3jK0i3q3Yj+enyJ6RxXn9cGDNrbMtrXxOiKSV+88+7EpOIifCEgWvXi
xoFA1d+lcBq+wSKweJzlOLsXuojOFRFUrVYfl2MacUlIFJ54NNAjFwu7FLOHfbIt
VIYAkke3UT67QE+vPgM4xpStOLDByWifSVHuK+kuI31ZkviVRV3mU6xna0y6DKK4
fdKe/TTWZTLkH+CNMkt+FH/W5tnJ2sqz9BWhurK8Ts+NZcBmrB60AxEn+wIuKDSC
zAwJK1aX2f8V8UBXc1NQ28uEvWJIM0VOVEsZYAlVEY8XC132/JmnEnDphQwXFFpj
EEWGMtWisqBu6ZqY0qKe9kSaJLUdc4i5rzr1PxOBTmK20RZ0HEbiNwyH63y+KoZ9
a7rmOHaTF2G+ANpn05kjZzonfkhvE0vCYI4uDxFmj9QCkxZy0H3XSTsypOz8Zx3z
qCao2cc3OSYqJiKmuB+wWFwznJ+P9I1Tg+FsRNyg57dKK2AYJ/WcG1l2gc/W1Ufv
rOa/3UC8UkyFo9colQCkLWMcVMaMRCHWrP6xsiOrZfiMb8DgAkx6s6Ca2OcS66od
zj3/BouwluQC3Q1tUgytGFW0zpGF5t30VwSGsfgS02OPSW2Z0cFTfJD7pUw8HLBC
i0YpESEk1tv9qvMlrO1ftN+jfM5LQns47VukoPJACHi6s8p8SZjPX98jQtU3cOHY
4ipgTA3fZX6oEpW6JR0AvR2weX2BrQFDVwExEsmOSIRardIrNaoJnDwEmwUVLdLF
UvwZfajEB/7ikEf7gs+lZDR+apKgZVZ9h1yxcHaCcaXvS8QsreefDz2uNDUheA8a
oV1aVzLiLwOgj4ItGNmqaebVzr4iRU2bKUtao5jki7PlvFGdrV351u6oUB7ac+xp
oewKw0UmQWP9zoEW7iC37r1EzOBfWdtu3xnA30foEQ3fV0MwpLQYaVgXIxv5zWCp
qjsmpl1Miz8ikZmqwArzyEdj94aAyFT+r+LxA1/Be9RySsdHscKiainGO4DdEB+Y
ExTAI11yY231cBl4OoXvNuakBtUrUbNavXmL5FHRQK3nhqpJl2UlT8DjPD0yx8iJ
isIlzehnj7UTPVj2YeY8MzfphAg3aD+LIzh7dqg1fxrT+3/VxXutoi6XKobT9rAb
CX6e9wqDnqmjPs82n2YVS0oX3a/B4UJdTVt/1ZI7e+t/Dn53cw+oZq8TQlTt1HXR
pGsi+0hJJ+Qr/tc379emP9orhEFW9pgbQHWB6mJZoQwVvFD0QK1OMIqHyZOd5Lko
4aJ1bXtBSDUa3fYD94sbDx+O2sukLYmDLzfRPqyoVgL40q1E33arI84SHAixVxFs
ETtqKP/KX22pTfvLMyFe6lRtcwsv58dIMIcEtr6d6HuzKcfW0Xw9DHvd1J5Ids6V
t98CZow5A9ijf86xxTIEOFFF69Hzr68BobogADYJGeF/rM2hgyG4GvAHSGETKqCg
GWRWlvKs94cHOsQq04HIDRBoI9I80QEyfoyDUNDB4vQdGjFNTFReXdyUFGIxeM6t
3oL7eWMzm5mXfd0KPiqMo2be3p6NjCJ3IpggbYKsL4xq7P2mm/qeS8y9ySsdb5T5
TTHn8dXI1/c4o+G/1OUPxPa5wREupO6oOj9DBi9I8sOSRXlzgphEXq9hEivor5MZ
qBLFAPSfC40ngD8cWwfIHolCT27SYoNXs4TwMu3/+tZu9s2UcGAmQuKa5lkNfiiw
E+fVnbJ+peDHoJBt6pPAMJzxSYmYSxmpnUo94ELUV7FnkZUypTsTi64pdQyUale+
871Re5p+WoGCfo1zPevLD/1JNbFAdYXYo2h0Bhqt7WIcXjGcMr9CpcIoCh53fTEj
JWmi1t7jDj6kwdG2QMpi0mnP4dNYej3SlXmAnHRzyOXl/oehzOJ7j72zrbB2388/
6oHA6LzhRw3hRM197pSguYy+VsQTyMGJwxhUrKVQJn5FjqeizsMpYYcv0YKaQTpp
+vFaOYlBsRuzQ7HQHjkGgdP2HVJnL5aaaBSdh/N9sgMfJpcxIsS5Xz3968KQmU3t
bI9xpvINqz6w+G0QXgzEMqzLBnja2bulNzPyXZW0rell6BbIqudP4Xs11TtFGHSP
DL9m6tzvWUTMn0pV/mWqIyDQKjVWYODVDINFEZxmJaX7irRDQdBDl4lpv1GlO49n
b1Vye0p4EqO/YN8PtPSC/gw7uo174yGHLO1CJfWPH/ach82sY84SJ/NpVLeGsr9S
zJRWgOcGLFJDUxAZE4ogRxIa6AA2u/7FOV7Y2b9xoFbrxcUPAAH9H45rAlQ3KVL8
L9sfhX0tgOrj6J0ByQmwJeK6g83XsQKpqS66PiyWMFL9LYv9/9EEZCce3ri05uwK
Jx/ELBy292B7iHe64VBNyYh8xll+5MGbkhiVLFe9LMyR9FavYB3+DI+U8v/9h9GE
MIODqZURgp6Y17LWmK/RPz35cEbjm7Uz3DHoshNcO4UJYXMBiT0WbW6qQKZkUQJk
PpHIrkWYVNzj2SOICqTzb3IL0bKCi2tZ4NQYgKLivqs42bYD59ZVl6MS9LR5CdZV
iwmRduEZP5gloesQlVSYg3ih73CT1YlFDChn85fAZZcVbf6eRuwot584qppCiz4P
SjBuYU0Bl+IMKbJSQo5yOB+evQrMxNN3NU7OEtWrFYDXusBBq8LOn0itPqdkMtlZ
i+ExaBYXvqlko7yugdCMecsS9eHmeUeLfTNuQQH6zLoTdRdYEXOdDaAzthcoUDcG
3TGrfKB9cSuxww91lrfsPEzR3KIKIiCMmqkiRsjvNdwdyRoP6PQuSkegQw/BdmUV
lupmmpcO0j9vJTDQ8vC0LHZnw0sCujhy0IdSm3eFueT/rVqGbp0KIfErkCSs8DSM
vylMVCGVre1JlcbAon9iNG2KmSiJ6vWRuNt88l/zKAvjnUZ26xojbj1TRKJLI1Kr
5TCgoPgu5cTGfSzUYDzSJFsauHKebeS1E4PEbR6/HCZCP3AEdvAOAGH7c+Qgk+43
VLwZh9H31jm0biCsN1VILdq1AwA7XwOn3AUvdDxpYPoQRyZcTA8woIfG/C+ZRMk+
XZXB5BxDvr7RDp7yqVKx8ZMTjCMeR3bTwfEFdy49qoJV3L0BsJ2aTSI/njM5KE5U
irZfuQfq9p6KIcQXRm05rVrfoiq00zxzjojnIYwxE5So3jkUeAL4kybmp2dkhRV1
8koB+ZW9iMeGIyTSbig9T7Ui8SJLriW58h80ootBGFD7QrksJ3fH0NVzTuVxyhkc
2RxedywUzaDc0vKCRjcC1Eoxfdnw8GDORgG2NRWXXGHg7T4JnoflI0ZLGYXpjQW2
+Req0OTBHB+afoODs1u9Ia8iM9lxIzjLCm8OJSb2D33ijtR6jGpLwUmdrD+BTLCD
eAR1L3PpqbU5fzOp6jsSMQlERBH/b6jNxtKrHTQqMIfRBP0IAl9TiX88fIO3krBT
VmSfwyngsfNBOHYU75pgKLyW0ia5mdtb8E2+Z5qI2JIedMmbBquUNjvB96sxX11T
jREXgs+L/QZT03X2qpLjcYx2mT/eyWQSdQcyVGaRwlN6jwmBIPy0Bp7HYs7Z+Y2D
1GlQc8jeiES8wWhW3Td+f6ObGLKaV99KKlMEK09HXEwy3I1TtofB88birXEj8ow9
x+U5MHgGZpuDZdCdJ+f66nUjiSer4BBhF+hZKg5tVJKy/O3Zdd0R0Xa8GOdaApTA
EZ+artuRVslWtgQoUEEmMNyHrQPCXvUpefNtu+XwGjRW9JdNQWraEPQ7SP8ctZQZ
wAgmHn/e13dP1eh2LLRVTyMPrZb/agRtKf4G6c1RqN+0JRoUShJ5DzZ2Yv7/yd0K
cGtqizVSadr21vqh7NI6zhBtBd7JcBwyPFQZdSHBjnNm1ZcNYHAt7lds9twKKsxo
mMQ4jrXuxzChZ1Oi/dz/ED+xglfX2IRgdT4EsNrwNQnMwSmDHZBZXPP6uhYyUeOA
a8AJbfff8oSX4c+LzoFL+s3+0AJp62ZAaf8/NBJUVJFGinf9aoCIy1pWfUPnF/9/
tcG1noGI6Bzm7guHaMJ0GYaGqYI28c7hpwGH/QoEEV6ttyH1iJKSdelrdUR21gW8
9ClNxdHwmJGpMzvm1PEP47LW91xZd8UQCXXO9e0tdHqzYedcLnruaawbTtQjPCoz
c7vGnyIrEPjNE7g9jpEaqhB8j70brol7/A7O+h3tlr0hqYbBRxG7sAWUJhpyxXpk
bQPnMaWqhlX9/iMJpRuaeFOSL3l7uswVWv08oNZb4vkqvGQFWKZDEPtvZhSsXKtW
JPSK7QRsHOBO4iWYyFjuypKozTsGDcKzcfdMSCjbfyEfV40ih8jc6eJtGA5BMr8g
PTjEyMC03s+5UBoTfrNqQJtyrVg1Ne3TI6/J2fw8ellFhqog4rpgdTjo9vUMz4Wx
8JM3e8BAeHGydViUtmM1KnAZwOUYYRjMv/rc0Sco7m+nQ75na1SmFT+1Jv3J4YVH
BKz04dCxDEiTivOMCCCK8lShPD24oH+79ognhU1cQXOI20LI3xXM+nD/ChGEz1W0
0tlqIbAtgh2IJm650Y0zTQoKWUALES1cezW7KLJ0NAb03rG5Wf1R6K/ODmfysO0p
h2WSA7v0iJkCDiD0w/bnLh1yKCAflqAKfxqoTYcQzNUweOwHoy5JRM0c2B9kzMpZ
P43HmaWezVtKUO080r9wKsR9ptGn8ZfWe+0j52J6tw7+RKuSFhYSslgkgTPGc2jH
usDacNroLs2OX6kpboYp2aXFiE3/ECeU+dMaVWQnVthp5qPj+WlYGSd0sK0AN7u6
q7H1fPtHN23x0BhDZSI83H+6vscsD44URc66KRTjPCoPxBL6Pxr5Y4dUeemgifVn
gylm+RCA3u3EUTJfaqXoj6XwSLi401ABSAh8qpGrRCjBTL6QNSOaTlQy+w7zNmw5
Rvwg4ih+Lt8AsYzsUHqp2kwG3/DsfAZmsuPntLBKGzHuzMRHlaGWugVFiEDm7gvD
0iqJKRiKbQgsyfliOntbWOwLsY1BFhDAJThRlOBk/M/IvYTV9IKV9HlBL0/e/52E
RlLzQBt0M24asm3T1xMvqvVORQi4EucmfrYGSWyKQOw68K0fDYF2ghT1zMZEOaam
4SH0hAD5kpOLV21ITC/fyHnbUwzoihI/Ukws3OBo+vHTa15G4mlYTIsWDHxKtzsf
dBkMDyyM3MMUm3pYVfMyc1jZa6reFRPL1sDb8oSR+FQKticlNVdkgUF/4W+vi4iv
tJ+xu3GEmWVzvM6q/+8RoW1BGi84IMjYCGNjJcZeOFrrxsPJC+QjT7avsng9QjLe
U3TglqEv4jI8i2nXJ39d2l+Ye9EY8YTtKvtLtJE6M1Fm/xEO0A+pkL3ufOPiTgtu
ksDQGu5jSpPf2rDZVoDfazF6p6i2HkPOTQNvT2yu270BWrDRDQHfTd/B5FOHqVWN
ddJYRD4nTed7lR0g5R4Nb139Ow7IGGt3mDAgY3k6wxKlW2EfutXT+noA6lwnaag6
oRdQdd3qlrwAAMKBF9tSaVXbTrf78s8QNXN/VTHYOe1ovSrXNSshffq5LPNBlvJS
SudpRX7HnZSBOtLu3nDvNgz0MS3m33306LGbDL5mc9KrfB4hgxzCxVPhNbsu++Vz
eHx7s42kglDXtrVbbTNniCVpDSnPC12+EHW/W8CL9fHmPxChZSxF5/52jlpy72o4
85La73uo6sEmSWhxl36yTY4ZX6/W016De3W+xZ0XDHTDwO+rnKdqCksdC3+ARxe6
Cd9qSj0be8NRH5ulpSo+/bheeHfkG5YJJ2HrzMkGc9uViG+mhOBu27amFEZYnTeJ
7ts+WI8fxil/Vvjcuvd42fGHf/4RVdjTVMLbmSg4XOXYhOSUQhElzgDu2c4j766J
97cUY/+C1C267P7x5nztDAFOkz06N3Bf/IuLXG4ZDedF73xL+HgbGLG58mem0cRR
iqr3wNwkialn8htD0Y1l+pYjOi52A2++803h061aHJ3O8mqAakzF0obHB9TitcnN
ggYLeyEyjhnehoRFT7ncisOG8OF5BVaDJTy1ItIq0sUfD+frbTqmpPpPNDnhN5oa
Jj+MrUgACLu3dM452Ik7ZO7E2/AEIKwDFJVQizzNqJYFy7U8vMbEORMLF6h6/XC8
tmZ3VbQ3jSwK4JGxYE6yWd2IV8K6iHuZcw/NDd2HbX2Qp2hgyYRmarT+PRriViPl
T1Ye0EtCe3xZAZ/ydDXJdTdfjPt7qu6YTDwQQM5jr3fVjYooxFzWBkTTAZTTeDE/
2MeHklhpCfIe3NQddydYHGaTzjrq5EtEKMg+ywRTRQ2/iF6zOhycLw8cI4w6JPGA
FPhEFFRGOvOrXlPwbRHWVurH8uoBj7st6wdqarhHYaQWKPWphtxxg55NKNV9FigB
VAhbeLBWGCOU6osfx+p/GDCuLPQbDgLx9daXS3y2sVAQoD4YmvegTeV3EqmodO2P
qHzIg8uDu2OKi17XMP5M8MGiDSBSKZ1YzOUQGSScloH+TG1A53cwj/TZlmHd8oFU
LUrCBcdi4iAub70ScnIR/6RuIpAXxmcfUNpnmxXx9HtPuJWRpdiP+sEgBAkiedX+
4NsyFwXinB/QMB/xjxMam70zlhfyr2mXgYxdwCsZUPI5dlQrWvjiUha4UfoB4lgZ
WFoziHgi/CMFwofxyjve0MB9pac5xm2p3/tE6Wexb+YOQt2xN3XPwGOP+nN8ATj8
HIeKEGQYRK4iQvjXxh+UWuU+19WsvtkUJ0ohHfuq5ptRg69LegVc73u+iGGzk+sH
9zctRxMWyp0NoVmA7ZLTgvJPCTXgjc9sqpYqeX+fMtDWWEezN+EPN0OJlQDtj/6H
fuqSfQBasz7CJfAaqSahZ+zgeR5ihnTC4rbOU52dv5kQqAMfzgp20+p7sA0EjrHD
uFpq2kC8AsZY8Ijc+oLVk8cA1z4G9ll/kc3kKsh5VCtkUzrv5JSP0myu3yfQqRGk
3qgbq1Z12qbXnnz3UzzxrwufBUYz2M6x3lQWIo5ZMEAu+eaCLZdiCWliFH1sdRm5
jAtN/ZLU2dUhmMn+5HjCbEsySIkFwQXutme0knksZ21V9vOMsreXVISt1M76pJsK
EhpEuQIVHPwySyNGmykRVYcKYBv4VjQcfdLFR0vIz6Nb6B16GCJRs1TO/NGqPGiu
O8ogdTSIcxzN0r+ApArGhgqMJt3Uy4uddQu0kvruJAbj/lwlNp+UA9tyxsMKIOmp
bY6kfshWd+WWjdSHUCg8hTp7GhLMo1Sd5uuIK/kx52TYje7BHbb0feHhxQ4njlry
U7Hf6jDsjnudZcRiYZUmEgO9PosGjYhjXeyHwdLr5wX/+8kbnyHSDwVNrFY90Ck7
OJvExg0fGUv8ydzLWnuOWRHDpyUA0lDn2k9Dip+qQ70NH57h3kTYnBTSsRzjz1aY
p1wrNv1h813RgqH9OcgsG6JUZudtYSxoCHs2AwZVDbIEW0qbHCYcUvNhZ+PB+1Ap
6uKwXYU6HGmlkmfM4bzLTLxIRQ5eURCvWbwtNV/dmAkNa4y26ZHE45/kxHPykYfm
yxUve++wPtR9ovZQ2XDrwy5lmIW9o8EJSM7cz8OCQxpLaRAfTzmxFa9i+CYGbnNo
O4LojXjxSO07GRrkjjJs0X9Q4ZI3kV4TPXN0hYQDcupdiJh0NVVSA2TV6y8RhVoR
Gbrhi2A9/F5md+Z0jO5MrATu3VFYMkGH0ZR8ykdf9g38w0I3Xz9oi3kzhLUpKoP8
GMXs0MAawczRRTyHs7gjDulfORybbun7xZe+RdS10XkGJOj7yPnNMJkTfem5K48r
MGylM6s2SzjanYRITRn07up2KbW94ZN6HHb+sZDhKg13lDKbOpxfVnb59cGC11UK
8kB19T/jKoArND7OgFkRzVKgdyoTIu1Ah5p2tvAjDQV32sDwHk62OTw/3JfanVfU
napfrxlQb05iUAjaUNslJHlBiDChXVxGB4UzWZgSNm9xW3oi9Gyx+2dDKuSZXQHp
Yh2txulsopjfGi36PF1KbSh7jbBmVremDyEs9iTZKXqJPfdvaNNP7ReQav6q4emO
0Zuqee7jk1BA9uBISjQN+4r8oWLkhrgdXsmW3d3HrHHVdUwoPTrFGAINWz35TYxg
xugQammFsv4/uZ/t4E9yp9GJk4Z8j/LtPLiapw8IYhWt3C8ZmYSB47VMsbqSlNkW
c4sws/udOFAmC/ZBP84wH6EDmev8zfFVW6jjIJnBkkStfYzMD16AUTiDPzFJiiUU
rTr7z5g0tZUPcaiIcjjprx1YDFB1Ut/m8H8cshp6w9tNStbpv3xpX25HVgckZuzy
k7JsXqnnOsA/dhl+o+skVDn9/GuZ8NBkqalv60p+hCwu+0F+siCh6jV2nzQWt8g3
PAHi7MJMOq7HJ0V537YTmONduaEhxmYON4bZAanCChOWy/9DxFYJP+Br3dpQaX06
mssrko0Ilb2peoIShwjNzdfDecsLhjcFhn/Pm+AIr+HNdbv0EkOis4IHabkFGEOU
1Z47oPwcAJOTXegDXpy1y9ud1qvKxqWaXcjp0ddU2JRLiRJMmIL3CYkK9GP0l42S
OLq1DBRMOpwECch30mRTiWfyypxGzxnMpx9cB+s81MaCs4sPkY+lDqORN1tZ2z84
JLu93gDerE4b0C4qGGFjNKLBbDxquJN+KeRIBR29KVW+mRwq9EwwNAfPMf7K6UeX
3LCdgsAu9R+k12EChIdqrrRygmLF4PZ7RaGZxdVnAnI8VFBu067RMH13l8vBNqGa
s8+Jn1RH+GSltGQy5hmuqmun4NWZlIHRZCUnzFLzNepnw7X7+3WBD9eLXTs75/Ia
cOdMLeDFKL+2eNH0IMGO+RFn/Bw8jAY+aaGaz+724oIxv4lHZYinILw3EtJ2K3iN
CQyB2lzDUSsUhWk5BMx3T0PbPYQ1jpwQWlocM1I72m+S9wAEpMx0ZvcIAL616efo
o9WkPBlnYGbvz9pSrGxHsRgJkCPtiTl5XCJ94f7V91pyaDSksmSC+dCFrwBpC2A1
tBzbGGSPrMvnjCKF/C+4cZhv9dTsbJH2FVD2dvu9/3QVVPnpKs+9sWv95i3PlkJV
uw08boZy0axTzrJfPZof44g6P3JVwY4OlJavo1fuvPexZvBx6QfrdKP8uAZFg9CI
xTpFnDSi8lFOFncPobTvb2wH75ovrgy3p9HDSnYA5QY56dI/ZmLdIVdYUFRdZn7b
PwK7DibviQqjZEH0Iz2YxjqcGhVGucfsNkY0kZKlqeFqyC8d29cA4hmdD6//g628
gn70qCLs94xqtXIOn1Jls/Lx+FrFRbP9RcWOONg5qVlKQfE7p1y//RVPhIAqVDpq
Vu77kVitjnOL83SRZ6fGAeTH05MqINf6SU/dBxOcOtR5LUC7D8in0xlGDdcJs8rl
x+2nRQvh+9FqnpYIYkEbYUTg0T3RKZPK4uOATdqOOBXCYqqvbhiI94Hs+3507W9+
dA4YDwXQ216BL10t8yv7iuiIE7WlHXgedFb18oxPG6PJHA6mSCbB6D1m8B4JbXCj
2C8ky1q1y0EcV8Ez41NJ2EqOZxS++vH7Gll4AHtpTOVziXt3/RlYU+POOG6BPfXZ
+vIgSnGeyRE35SAZ0TyIodKVk9+4gz15hHZ5Oco+FjHBEDwfoaMb0LNdHAYD/GtL
IrTopVSBjgsKQXpJ92s1pOsGTykMhsLk1Gt/uuTrIEwa/f/0cw4XJbAWjqCX655G
F5h9ApHAiX5Zy04FrNq8HWX4funOlzVdKoaMaZUo3N4EBa0JPqBqgewbQmIh6oVi
GVlALPxM20oAQhBl2IaOs9jw4S29zOhjYOA1XQitl5wlBDhhgElHpcxMvSObeDTH
NSn2hUtGl5fKWF5Vh64hucrbxHwxXevJYCGVt+EEQVEePd4/Z3MxoGMbvbMorF8j
zv8O3OakCklOZL+MMSDrJTUy4MoV8p73FevnDcJGcgQE/7tmZWjT9OzQi5OJ4Wx9
QS8uor5TnPiI9YEhrk8CnhPgMiJm06ZdXIqalEBdhNYk1UBKbEYbCEI4K6lVB5nR
3Lxk+SeJeR32XWwy1nU3g/Mr1FlBktIrtBQw5LqKHihMAvcLVH8O8OSBo5IzRQd0
V3Oklp2gQrDehrXcjTtdK2Ssg54XaJMih7yAYwivN6ze+cg9+qgU1+6edO1sL3xl
Xl/wNYypZlcOlbpcqybMgbz/gqSjUqLe6+0gGJDvY91i0qCH2X+DYgG5K7CNboo6
MVVaXBQExxKRTgCUIcaPZZLHTUTR34Qi5mJlTm8iKA7o832EO9G/JkDIWoTKhoBd
1vcIC0rz8piBsdssvtVGpGGm1z/5cCFKvw3Ev4XZyj98FrlmqAVBvF9/0TDupzrq
Wc8MUTsE7sNfeqJAUdbBiaxhgNqd7aRed7T6bMkFqpghlLUr30/O1rpRmhm42Pfa
XHR1vZn0YsIwleGNpT0k50wmlMaNgrxQhbdeHnwcJJwWB2TuXKD2siTfTsjTNuDR
5GnEm0bqYZeANNyUyny+wd2exVWHDErJRvLX1i5m/uVeivbrdWtQiXSEeMLK/HrK
QrbkjONQYxwZAOuHmzqflY1hQMrCKea/39JQnmvaPsyUzWTzxeN2Nx3GM9A6GaPR
pgDnWVoARyQWEmKFPIKqbTVih9l3V0g6l4BbMp0M1/HQxzNeddHaUv6xlNwLY5Y2
Telbk5Ecodq7BzgXXhMyiuzaylZP9Uri/wDcxUb3JeIW7jzhqoVuFwbn00J5Pws6
fgC3umBPB+z2tKaGwZarOkQiNYzFHGKfUyPH1RL+eDkbkM5JPBjJ4DHMueFdick9
oE+T1yWZR3RgSAoJ7vIyyD5jMk4zC8eyfKnz1hBHI4UH095DTjx49bjDLP1i+ktK
Uc9WOXWydpjfJM77MAL38nmK4BFCBO4jSTnFVy3ct2tk4+B8AReWAITlPi0zGNFo
kRqO7udQYZElzv1dpGY6CDOp5xn0WiLa6Ylaua7s3gt0C5EWcspYyI7AiLlRV0JF
NMHFvptgboqLndD3e8Nc6fwCPdAD82GqFD5LPvIEYszlI88S3KEJ6VAkbzzWbVpl
KNtybn1Zue02CZkULkj0LJfpChWx+fTB9Wcyykkfa3lNw/T3aOUnbX5/2aDCur2x
oAuGYEgbSCF7BWPZbkQHu1i2tQOmdWJH5cop6AWZ/MUMVsxhlM8nyoACG35xLXQI
lfUNklTgDF0w4MWp0Vo2gLotPr/ETxcMvaxXhC2lwrNlxMAxnDpFPP0rS8F4rvFs
1FaKI52ZE3bC/dE9InC4lhONpscpQihNrlUD6i3F2qb2S8gUFpIQFGf1Ofsgt2Rv
ni0JvTpOltvSfibzqZazDnTfFiBTkUpafxkISqohsnrMDcWkRSvTnWmZIf6ISd25
oLPzJslFwZfB3whTeJtUK/T0UKuJzfrvkknlofAF3Ykaw384+wdQfLUAt8QNZwJO
pmb61C+csMN5BHkyWF1NU+0Jq56DyB/nkVcuR5kyqZsC7lU51aKcUjIuDiDr6BAa
ZAeX6aZ0BpP4vourpGIBdfMLmdUozG3+38wY16hBrFbaPDINuLTR69O1IXIPjN8H
7G8tHdjmEKHTxocFjPsr5vz0679n2ffP/85AJvPd5PCek1K8a2dmaTaDpjTZlzqg
720qHVc0m0N7y/q5eQ0GY5Pa4iWsxsLBFIKLQczDk69ktkcOLabefVaAxipbJJM7
R2jrMAvIWdfCPpnUD0nYwaoxZ8IcDCjVhl6tyZqsZAaKcFX7slFUqkRZl+Cxp0qN
jE7BzQ42eyi05Ti0mBltJ7zkXzXejMAl6JJhEqTAq14eEuCoRrtOg2xSo+V17vyh
qD4llzTzUkfLttAGXQmgjkCKi+v1lGNOn58QAL3CziQrDCLPrOb9rit5P7+UmRHl
MzTAtxDbYXaSGbkD2xw8n2Cy6cTd/QAZPC8amsFRd3xtjVlvPsmBbsiBpCBUUust
M7UB45fCOpUV/i28JpYfKnCy726oedBVcSoQHWb0X8aI+rBd6Jo8E0Ift6C1jywS
bMQ5wrRaIy2q6H2Q3s3LDUYdl8uq6FTwH//Fy+NUwlApvmd+azvZAnbRd5ykZjvR
6+FZj9fy3yDyit5kNOun+yuXRI6D/OFxJjwfnoaNmWTtiGBJatEOS/4zQeMUIl7N
AM+RTlLT88GbAgzhUFMqm/G0OjUl3uKCU/evq/Nq7F3VD3MtqBU3zs/I0bv6m4xC
53c2iT/3uFBU87gLQKgyzycOW0SqosElPBFFMFWiLnQ0/iL+aDmtd9l+GinhnR3A
pOcq8Lni7+e9qP7L6Tit1oRpe/4Be7BhjrNzMNdB2FkLO7pxKYcET1mBSTMW4N+4
YmhgBCdGpAWlmfler2z83xHjeSdpeR7/CnKDnBFvtCQ4sXDr1FsCVNsqFVNjbMW6
PwDl0tpQfc1I7Dcw/BCvnDtu7YLae09BgT/nJMaUFEbhTF9xfooXcllYaCgLKgl9
6zkRY60JbxEE1X47cMef5JfPQtyUdCPS/ifZA07PQQr6nRc3tiJHf4vjBWd4QgUZ
njfBlti/5CWCD7+qBjhBBkmcLH/UfxAlIWRlOp4dr0UTLmbh7bdntg8d5epc/tZC
eALVsxdBuqMVS61WSlWPCwfzFfyT3LONw5iUxPIHm+y8abaWYt5J3bEJtGbQTnM3
ld0du7SeTkM6NrFFwsc4foLQw/TNvGT9/WTVP0IBMXas5diCyFlCT9c5w3Gwitj4
vov6m+GGPFbo1xVtFmhDfqmI5ybHksvlsHKTz9yR6+vtLUaVwShPesrVHnyFEGOh
RFSPv6ZCQl/Rd1LfM8XNAKugKY/c1B4Vgu7dTEwJ16ERsDoKInzS0p4QKgvbjLNC
mdlG0kstNSYPoUSh792lhwued/vlCE2UbEGDtZrGynMA9EJXB1+gURQDwNy6bs4Q
Q0pOlfZ6juBcTW5Aw4ZP/LBj0cP2nES+qJgK6JumE/ZJC0X/CWVMwpbBG7oFpS+z
0NecDKc5zfhI69ccsd3mDHf7NTqfxFtx1VDPhLrSWFxn1ggQ6MXf8xJFK3FpRaJy
TI/vf4zsbbfnfb6H4ySbnsoDeDOt47XoVT9mt0jfiMAwu8lbIRM/sCtDV0/8p32K
vyo6CbtokAaiqU/55D61s7CCNBVP1hSo58nynraX90stNwKPhjwlEUdrz6ECMfBw
5HmOMNp3K+elU/GLrM2kzYU3ItBwC2T8culgUAhLl+tq5zEt6fGzfiqAfFiSgowy
rxlx5gZhnqUCC2b2U3+f/Qb0y5xxqVqAEvk7Kz7515f/6ZepA+r+9+QBtJPa7UGJ
f0fpN4OOLVlf+Bquxq9m+xyLBh4Cinwopwu6AxNruS26cf3Ex4yu4/Woi22x5t7W
3Lg4BIpKq2MgAv5P8jCXWaPFwfPhjj1+HBNV723qwrA0yzFwGT8Xr+4ghaxWuzy8
Vq91RNvCsDn5M4lQ3PlwOPNq3I65+D3tzHtnQrI+Kjm6T7hbZUr/iBRsgN67hj1h
+Ol26X1mSctp+q/UgT+FrD+J6AVZ6q+Y2ESbqcctgTkQ8s6Pf5OXfcKyTjz6BA6w
cu4DXYwXeyXUGwQcLWcA2U4vhr1XpJIAp60E3vEaKiWS+eXOOz5wZ47S3XiUkku7
Zk7qVWEGzfl14l9yoQzzay+fEPm8Fg4Q2wNPuiF9+DO7usUrtMqRJkl1HUtQ15aH
BEhZ5aDjWeHCq7o3Yb1S5nohCC9FzMeXvBW62eRy+jTA3JN4kCN/j/4wvMVAE8EZ
1l4ZOLf/wEEqgogduYzV2AsmJXgMPxNDrsIul7aMsu0htnTlxvf/E4njMTDHMYFh
SLzYPCJ7WRpQCiPhsRNULdL6Qb3Cy1IW9Wj5BQAwKK8FC+XQfYSLnV5FxoYw5aOt
lfBx9eXBhvQxVinzV7kZ9qThgRUfZkFUTI0VhUSKHBOfY/+hUMJkoE1Xig40Ia4r
tC/XaKMV+Qy+XB6STDutuzSZGfRA9BPFQ3RH8NLbS1XqZ+cgyaPR7htyL4GZz2e8
GqkrWwBDaRHdswu7f/6uVhBPvjjyeOZr2lofyQ0ep2TortFpr3mb3Z13a6HoS/n/
c62lq55ziGSEFjx7OxI0zGdZb7d2x/SxAT1u/Ze9kNVcWBQt05zTYmkXAnrsnK3N
6L+OMSRFMxrTotFCG53Cl0T/gqhwPDvOS0ETAef8fArG5XnYHKtL3h2qOQbiVWZ9
sHUKvcMVNxEKSo/iDMH8UCclu7jx0tTs/6t+vDkOMa8YmWd2XT/Ny4PGDL5EBZmW
FmItGl+5Cmqvt+0ugNicxyl/FZpTUxDqe/vKz8hDsRynVGuSGfmi15s1z2FiQAea
ZNH9tiO9NqhDaITBUV2KHf2yhlIsRJyMMFqXIGdVwfSthmuoY0rX+gvRYHTl698P
rCK3rxOAke97qOYUUytJ0KxSS5ejZA5FWqG8tb50SSAGN/peaVwSTrc9vg7AkmNI
XK5RflImByiOWbq9cQk9q0F22QQOPRshIFWG+oACeXdFGhrlQYq1GKO2Ua0RyiDy
IwHtVHQnIE53rPadrYpnHaRQiOqYeAn0l6EF0onXNRu3zsd+E7AjioxU+w3aQCoq
3CoROOEDCWafmq0QKQ9CrBaF4GuDBX/cN7xZ0lrtAWq14JNVAj+AVrCy0fdg3tf4
ipCPHvvOEgxU7GzoG1DEtnGdENzV+a9quuzYw/grSpc+DaeRYW4/3zU5K+jyVT3l
JHKLEyPXc+5F2SIFHUWtQR/CsJZva/iTMC5K8XCLg9APs/QowIgDuFBSucQjm2Uo
KNgBZHhck0ZloUZZMQ/xqdh37BMtxpN5n97ZxIPQ0BWjJTVoSYmhOqYD3cnly6yM
4JtZa4PHM11y935ZsXL6bUIxxXUmf4D2Ib9+Rg7NQZtMchNtRBFWZlKcUnbKgl9i
N9Dz68efWifWcse6lcLQRPl6w/qmKy1DCvFvswsy9eKkLB195iZqxGO94aPjsOIG
9ZyxmnXu0baNTnEP0tlfywO/VyLrpp2teSX73NUl9Re6QoKvEolBiqPx0WDkFrKC
ex0ABxEkiOeV0OL7wBrEhwDDY6iSYVXf+HAXScyXGKHNcxSnkZMAJsGPTQCH9FFP
9RBkIoFVDTGO2EhbkSQokrkI1ukEiATrmFNHml72b7YlZpdcBqzWt8hMjKBfdoZ1
CONjrIIcY1zN7WJeq0xyUf/6yNptYzJngMmNpyIEOOJpr7fGc+Sw9TC9P651r4X5
gBKEpy3fHZRfVN4ygiQ7KTb6H3IOTcRpvdpWVCAzcQfd0uUhJ48K8QmfK1ZzZMvW
NhLoT59cbx5GwLwFvwCLSR6zJI8FTxznp+CnFYuh2x786LtQkmcD/NEg6NpF9IqW
QaSg8Hkz7PqOasXZgCE9NzESc1RDJxwHHj/LpkKRHttj8sve6ytF/08pDshLHYam
XkH/ytsyRv9rmxqbooS7l3Sj1t6d+KvCZbgz2x/cQXQRV0AiCFax0hudw7psMcFf
p65nR6mwJH3xvdsFl1Vbvu35CzEpspSHEpVmj+Bd/WpKFQMOMcy2tm7jZ50u8zOU
x9S+BXd99grRnjnuRJ9SQO82GN1fqwOBLhcrfg4xcDGK1T+uRfZUYHFcntyDkpyB
FgaTw1HH2xfa2R48wuHihIa3NBW11jZ1DdYHPmZABxFWhrPvooUbuclUFgt2kv+0
pffmROmy0Ms7iejn5vLbZ+YTylHPcWaxHgntfBg+qL5xF7P1oz7dGiSsQ8rctRF6
iiOyCfHbL6RmUp8nDJoTpOq/La5tDk/sXGAEf4BgxcurClGBfG3W6Y8wCiJqhqHC
VPVRoXevYU3KVIeCYD2cICHKtpmRO0d9gjWv6oX07ya5jHq0DjEY2BBpKrIMgWte
pEK/0dRaK8XLAj1SqzyFoUhkZvnPkiRFCaQZmmtZO0UaYcozbvikbujKUq8KQ14A
nPu3s4TVCDVszmIbOwwpsYA0jakRNXWknuWpWzh+V5VC8gfdWmjoKHy2ZhEidle7
52pd6gs5t3WQ8wBJvQC81EH0Q7z7rK+biwcuMPqtjkyuY1pmoHtM1uoawklwgc5n
Z43pK1PIwuywp68MiJtBsAej99/u3njMkY+mniDiTsJ9deEL4FMIiz1J/oMBQOuN
ADt9kMphbR5iL62IVhZTKzLd9ovlR+/c0Z+CSxosstJ1W+Dqis1k06HqQWlnPQVM
Utq21i+KpNhl5FTe9VZ9jxxZwI2AHXUQ3IZgNvBRonjZ6c2V1pW7s6BaOpSxP72+
V0dHemLUCdt6OEDBZLsRyqmM8HGKkSu/IVtjtENZaqTHljMBBX63Y8lrRGyoGx0u
54gX4icbvKo/PVVkn9oCDwqg9LwkIUWoVpNLxjoXwObjmay25lF/znz9dQRSPgcg
JWfTvrEytuCjK4QAL8qiue9KwdZjIcocvkGDdeO3ORsu6tj5jAn4m738u//Br2Bk
3lwctvB+HYPjiTrK1+8SApaE3iAM0PmQm81CB6u9et7qao8HIObxIOzdlU48Erzz
/OvFOD3e6bvSx5Dk3cG9zc2N/JEyAJfTVEMFZCXEDa0QkPjREplQQTwh8go1tZwg
9lLgaVIFPhgN+7+KmvQ5seIwaJYJT2L9sOKtt5pJ4f4whyfaozoBLJZIdijO1P3l
N9MJIbnjJQyQSKIGJwOJm/ddffrQwicagG0l+F0sjtVuX/w/9TDpgdBE1xPyAFJM
6qXBbtDiqLorANNmmaobWGZD4x7ms5T19PZO+K6yoDod0HyzUFsnBVIwMS3Zjq+S
tXjWxUeB9o+lVHloF1vqpCAnF2q7Sr5EDJteZYsdzGUHEvYTWgPMAVumz16UdBeU
0muuRVgTFgweK5PXQc23DLvoWJ7Ga+3mRdXkXOz9qcHvEZpxBuskWrimSw7xb8JY
wynPxmjvWfNgtyikqJIl6z48C93GXmmwihLqW6nvWNx8VMcPfQmbn8Uf7aoc6d6W
oZTexMSUkXJnKepl7u+45ytBP8l5H7YhZwzQSEiEq1tdHpsBnneG1OyKbX69zolb
+pV4OyhNCBliO7ZZywF8PkZ6ij4hWtU6imqkgf3ghz856cWbTxI1MaDOBvCuFlEl
DDMIkqfl4qhUl+gpiOZcDV0hmBQ5PaZR4XtxTBcFAgac36kqWDanw3q7zd4wZaEA
0csAlj+h9U2PYgqipAvZ1taaMXsBMvAsumkbPt80lWqO17OqqwiG97b48RAmvX8u
9KCXmnOi1uomLU28EbN+4NsZbnrxrYQMWy/xFaygdH+kNl3WtYuOn/yvk8ODVmgH
4dAni+Kt5W7AEY7vwEIXVF+OCdVOV7eBNzQRMdk/V2tfpFW7stxKSSgXyWXCcWLJ
tUL6FvU9TWoHJu1mKBj9Pt3MCZmZPqHyiwdSzUjWjiBXVU197KjwgSUpVcC3FdS0
mrG9ZNew0luNHzPL2EcNlk517A1nLsk/UoVSlQh3nSWSK+qVbuaMilEAQSXVffvV
uTgj8IsWxo2OziR5B7ug5SUdp1tHeH9ci6+9T/1DT8xHYTeiphI7EWx0AnrPaUZ/
8jAzK/WFG7yIXqdDQ4YBUFYYJpvOdXXgWFqvLoVMdLAnz8P4Ot8cGgl8O+Ckoza3
dHRQv+H94Mdo5WjeBKiuHpAR+Y/Q8S+FR/Td6l6wIsGiJQIMbfk9Vb65j2hPdjMx
BtQvsVZ0LPnI56XjMKfNw1vvXMmv46mmAWLN+4+8CU3MT6L/pCZ9/vido+dZuO/C
XunxHfD/4tmLLHN54vo1ed7rGCBR4tCh4WLhf8JEQiqPwCMEP021bwXuOZa5XVrb
+7XCn4DsfYEWKQRXn6sThSwT7asJeqXTrK1bTQvHs0zD3ZeF/Wlflo71sTXz9IlZ
U+nxk+Gf8DOrVw5CjIupjqfo2Jeq/OOM7eaRhixZUiOU3wHKv3cZtQzo8hGNREbF
TSh7/8WU3beJLixMEU+DQSrvxF1eHsnf1AX/EqG+MHskB4AnSASj9cguQMDjwJts
pvp0MuLvEgMRETpXBm08llJK7Pa6PN0fX+/TEhGuK5w+3b7y3Iu4Kp4eKYVW/dIc
kRrTGh5MlkKsjEuXAzQStw07iXRZPm6lFoFHO2eaMNNPzV8Jmy+0Q3Ht0q716k49
BDrsUmjjCo9tGRmb+ueSdRDLHHgUC7MZE+qKAUM3rtzUUWjGGQ/RxabR1N4cO/SY
nZUiNqXm/47tQxloe+LsgNb7l1Zupuz30f5Be/zGrppNtwtozY5l2/n2GQMgktAF
z8FjFWFlTE379l3TUfNzMU5FXMwOwCCsYav0FjgCC173A0royWhBMpXPPcx/T3ht
dutwrtmNFLyjrDRiaFR/8pZ9r4w3CWeug0kVv/MUcBNZQWqnHqf90JuNwO78cr0K
B/hE3Wlbm7IKuXg4b9mbRms62rStTCO5GYtcNWBK3s0HnVJJmYV/fgcy8w+K9VK5
q/X8dXR04UFaKEblP5ytZ2s5Yb1j+ohSatgve/BeN+l+vFYItWTG+6a5R/wHydUK
FuQTm3/ZG1ennJI3Adsz0LNrxULkgeedPTodGLcY8rk1wy9T862eVjuXYnEvKNo7
cblFidKCvurVMj14brjanMzc+7CR+s8FvBJzpKmrwXn/1a/lsdy926YFEEYhbpvw
NVD/lYBFo6C9eJXhNxlneKl8oR1jwqYn2eQLkbFjIB7Ld5iD2oiQyd/R0P4OS0V9
JqA6HKruFROWM3N6XvsdNmFy8i2dO3wn2KX+idq43MXU2VXoQNjMiAb2OlL/W3D8
70bfZTTfwxtNbFakQp+DRFHHPaHT2yBEeasqpEx/ZRzBvOgPkZqKuYCet2YM91t8
ZmnGoPA8BKa9TBmv6ILJm+zpO9o7bVqeQIkEnKJnPrUBRgvy2D89Zi/u4IiWJM8f
wUWRFmAQ0kynPw/te7xopv260Ry6ZCYJWghq6I4ALsoDxokdjJZT8fkKTS4zqaPp
5h0uH3SSrj922vgvb4Usue2DTjtO+iCaP6CVtBgjsvRqs6EUrO24UNd6+6DNSM+t
N3BLuV7I58YHPfDpzgpZEY2GrHYGuXj7ew1RyZ1lZBU76fu8keYZyTxGW6jGgZp2
4+KlQ2RTCu+EAhx7i4mK1z0yh1pFcPckg/hFUJ4fzT47wjueWVytlmJ3/WID6+pK
Cl94RdbPf+1CWJxCFuiWTabB1QJelncGeaa5kVIfhvNUx6nkD2mgqOlHBXPGigmM
DXQwkIhDa6euoorhLVHApATc+sL1PGwmLZwxI6FGNAR+nrKbGzoKor0CQG2DeCXL
FmPDz5CkHAClvtXeyNBsS4kRVS6jsgJnAVNPxdjuJvX5Nx87TtwzicZRqvs+05yC
j3O1F5wxO8kao6szi1BHMBtP4pfeN6HYDa/039j4qQQYDwdwzuMygEDUaMe8fosR
oryouD0D2mg+TNLXvdWdEHwcU63pqjqXddxX687jMt7wbz/K4/KA/w8XKHwc9fXL
pFc6WeRVuGYjL1HJanZessSTPN6fboTxXh/LBTn2URTwjBEqFvRGHvCPYSGlRDQ1
r0Ytpe5ui4G1VvIGOfJ1HYWCP0AsuqDVOYPC9T+5awm+0gbWHpZQoAY3LRMv/Ct+
WnaN0ZPx5O+detpEZs3uo/thiTqqB84r4/TQNk2oyQXvx2z/iZ1Zi2jxZFC1bUA0
aivPvo3x34NHSCIdNjUgLDpBwd2EFGrhhLlkEfzNYXZOB0cpMWVARV7MZaKRdEpu
6esBqp7lwJreF7khDuIGVAsuXAARH68AHRy5fHCZOhm8CV2L4fx8akQxOqoK1RN2
FrIn58NJ+OmSy5cijlmxhFq+0EOLQzUuGasFBay+ctAwYzhRETc67HvUwk4RoYSl
OpDCYUX48p0J77/7tf4PmCzbVFRayrdiTsAxTA5wNuVghKmeSF/e+HT2fy0kZutB
MGsNMv3aWMYP8HDuy5juh2fsVO7hFJoOPxW3sldur/bLfyH6pXnjlN3NoUPDd8ep
vZRmoWW2IEi/Zqxd9s1oOZ1oUT5i3m5j4ZwdaJcVYRVG6XDTUMqvvOjuyFWv4Vn+
CwV6K7LqlCPEqkicNODP0yNtp/tE+ancWFWrwVues9olqXvg3jL7hxZB9NUucACf
Gq6MSg6L37GGonQGn6L6JmJt0WllOAAhmLQ+aN5z7e+XSUtkS1oaecF51+XZVPSX
ehl21CmHCnJISdKCXKCX9il2IMi+EDLVG3pLmG/v4ffBRrWwQ3wQiLPHD0P+/zVV
2DfvXZXIghLd4kWJBp9ckJDJebBw58LA+yWGFFw7bBYfd5jtVLYOJ+nb2+glOn6Z
1a5iCu8PNfUn3lb4eIDhi/zz/GyyEQzBlQtE7VjRA9dhUOD8A8OOPhBqNPVO7adG
ijqvGXGZVEuv64AhHrsQsZ+1SYIyAz0ceWRL59/g9EkXJ7q7VNL37C/43vZwT1Li
JQ1FuVcIBs/6kAULFs9vhNAlEIHqvXBEY/cEpK/tta+VqjXm18dcnbogw/ej9PC6
ROWV/4VoNnwmWMSQIW1GcS9Ugwk7nU7xPgUTjxPj3WWnaL1vsHSC3OMSODfDPVVB
cO6QFmr6WsfL0O8VIZKdB8FF2NwgnG8lzLkcIB/pFFD6thN82fFnPQd1oiVyGTzm
qnqC6pF5rkWWlUzvXXvJBHkoHvczQNdq7dj6FfwzuXTJjeo6VAWsd2LOVSaVni5h
oza9coXH+BckcZ+1a8ckVRDqiogvY2q/5yepCpmTf2zdwSTmZNFi5pcN27il6q4Z
xkcM6DortM+c+yqO0wJkEYzXZaT79ex2D1x/iOxMSH8wfYQXRUCYIJQo0OSt2PFb
PC4h+VSU3NY0nexZLGcJTcyd6ilG5tOPOHBNmOw2PALMPOjQuIOVY5UmUKCFvC66
adOYSDw5s9UbqnS/zcB/bx1INpB1E4B4b8S1SlwzmZ33hhYDkBRHl3d71X/FA4it
8Wmh32+YtK1raO/F9QtCqmpgd0f8Oujx/dvKZraTy+oxZmNUbhxA2WyC5vJ7xzPK
tI2kKpBY16SPDJ8H2FOV6P/FqMM2w3FNFwz35T38o4dy5nnfl9mHlUHfLK/bVrll
c36CIYvbAOO5izEsiXYvurcSVyAZ+bRIN+t0Jyuj33T4Gew1P149N+a9ncxxVATM
6ABixxAhfV4SCZkJhqHGgav7jBqqpf8HlaD5lH2Oisfoi/BaveVt/mg5dYy1/Mps
ZevObByIBTFm0U5ySK0KDmSIXVMfkriJnoD0mvTj6JhAL6CbwXgiNjEPQ7bHTyaL
NC8CgfAkYGy6tnnk5TFLfxQoCX2bPLQrpRGnVbnVzbsFl73VnTImSTNi+A51QzMu
aEdATtzy2QHKv741HiuM0YUIZ+e4+mX+FU7lczeOu4WnlfcJi08b4E/4UHQqXrbI
tTBSLEmlomdayXb25GXf5YPkM0vJ2WAD5hn5jFtvcprdgcVh/+bxI9Q6arEpyDIc
GlPIZKjsC67oOY9O5rUqCdboV1KrUXqYluvqwLlhLZc4x505aE7ABQp3EFg6GIBp
Fky+fVqfXbNTo0fBIQeUbRLnbbXTVd/5toc/XLL7jCno4ncnu+ExE/XaD8rNPoCT
POh0wSBm9NvhuKs5ohPRPthuaIEY66I9QWOuNy9VCId/KTbNrP9QzABYm6ZwTee7
oD+mVlNvPN6yrqPBbXKW4ERVDZflEELcBVb7koDJIdDsPLrmfIT4HGW1aOd94YaR
IZpJ5yZ+e4FLuinj9+VQNPM1+sD1m1bIw/a1iWzWt/dKsSY54BHg7TLGfS7SMZPh
C10QOC3ENnh6mYG365929csxftw+PLpZtzv94artMKVUgvSQdm97aTVp692nwdIW
7F7LIE1tcWl5Vl7b+jxgvsucX91tegl3GOBNSgg1NkfM79+0B7xE6SEExgX+IBkC
RsIZHcp3Dl7uH6W0BnymMwWU+I3dzYftbue5mN32iVi/INKCxM3oqrUPMhl1O0I5
UFHWGfdW8aGWZjicwzt8fk/+SFuoyiQQLwzDGu8jHD6yAcJVLCSbzKnJU3HDppvB
AHLEA8beWMCVvbmZQ16M2JqXJMqKOomA1AqJhl59jk84A5XGaysFvmFkQTxrTmvy
tGDxOQxPubBG7dDGM9KhfhUVxSViHuO+HzfcXCK9TKjuyLpB8EDGp5RSI7YDwRaS
uvk41pbmXFRK9Y7MKOMKNe6wJkuCZdxgNNGIppNgB4brizTrae5ddb4eqXLYKNYR
8oqEzHl+Ni36u9VuNPsJ2xAgZvqoArIEDYPIHe7CZTCMpJVBiUQxf5h5cIQvmY2+
TX4FAAO13Ox1U0pNl2AgGDHbsUBBmvyA2c3TuXwlPJ88R7oL/uyqXSuxGUXf8DeF
Q085YuK+5nTrGX8xtqGyWFf4JR9b6bLLpRs4AEOQ16XN7Q1Bv3FBubbrhfNwPiaG
OsGKVRl1lLyacQF6iiAzNrXZF8h88iN09Uw7xlNgZEvYgob8NjgtUDEUhPDsyq/L
NhXnGirwZpJwkXVqkSHvkzd4+g0ppBx7B4+TZqjA+qzEgABuXlXoHNjm6CA1Joot
qzqkCXEtNkRqhqsiEWwsNDT9zAjT9uYwJxnEiEtPKmO5tw4qXYHmZSZ43zEiXzFt
JKOT7cEonAxBVRH6djRKd6k9EQ2AdGYCB+KOsEyyzT4mk5J+jHd7ef5IoPMCaW6X
v/agBI4h0GMeN6aDXpvjnAFDCeLxoWnOVLvEeOmjhPIZjuhUT3qPeZggmzNrLuY5
cpIZtoHjG9vmwdrfelJ6g8QltdVVPV4oB1GKA9HJaBgpE//lzB5xzty1tWqBeE/m
YeMEk+RAGOuYX/PZ2fum27qAMxlfaICKPEwsUZDw6qEhjJRlr/dxs9kzyYvqXh9P
30P2MRTmHKocD7FOnfq08Iyg4XCRQGxkKw3taMslRBpy65SYELf+r9ua/vxXQMaM
XUItz2oIgjE4faAyT8e4en0tOAbxztVozZpIMTvDUKW4YuMqhUf0sLf/S1RZUGGK
IvurzETyXAtYhIZs3iM6Mt+CfGuchJA/G3/EdWdfTD4kcH6sDQ8M97HW2wcSQQOR
V4kE0+eqrxGm+hVIbTEJ4F6r4L3XgXqFXLr4J4yhTIBIJEhA9K5PAcbHR2Yash1c
2fJ0gFzs0FKLmh6dydr1AeG3CQXYk35C94urjE++IHoJblhFBcFwOxQAPv1oDIEf
VEazdjzfiH0ScapFliQFaKgOUV7V7cQ4XFAkt4u9yUB5Ob7mVdnxxhe5hkrKjFFk
sn3FRoT/0fo6XypD5U2WQoolTzfLozW+pg1ATt5se0EgRViBd0d1ZRDt+fBd78BW
Y4tusJEvtFkBWIiSto5IOrCNv5CYkD0qYp7Sb0R9nXB/t6F2fGf6moRbLlqVKMtD
3xaavNbbqKypEtv5GSNdqnboworj6y1sTla17EFE9af+k+fuLJijvcKNwAT3DfZf
GxCOBIZm9beLmpQJQ2cgzam0vOs9EPQ1u9TNeE7sFLeu3tgg9nXYkkL9ekW+ufCF
uY0D9YAnax/i5Ib04sc72+yS4aWV9j2hsbTOTud/JAnpGf5Pqlhr5J7LnSDpJR84
WVm3aEVNlpWIS0AnNmWQswHJLMBOulkdf6nkOAduUyryoe7e5NKcPL+jjRIvmgbw
1aMe1O4WZU73p5TERSWW8ubrNCPF5N73wCNJL3fovKs8FlLgthub5vZShSm8DOl2
fJNLiIg/j0rQ7Rsq2lFfYvBBRI9Z/uvUMbmSf5vlau2yh4yvlXrlOavj96oltP4C
vOC04DE8i5YPOVu2WRnWkSTS13mul9BNEXu1VnT9lokB+vPQC98d6tvPXvqroDu5
j07tZ/zjCtTx/L11b6ehS2snNXBjEOeKvzW2eld6K/mskYqSMQ5m9eX7SHjKpC4Y
WbUTRaAkY8Uenoszmv/ORcVJYKrdYtFHvhTtJ9lz/oxsGqAn9D5WIk0TB2GFfdFD
DbLDuLp0m0KO8pi6wP1Elr82BQOyMFdqJtyi+7nCR4LrMXCFOMm+c5Dkvkddoh/S
FsNFBUz/j95pY3Fp8mZJIw==
`pragma protect end_protected
