// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:39 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GUtkxkWzEW8wyYFd51+2RX3Bss2ghS0bfSFEzooprsTILj7HtfTDSnQ4RNoN+bF6
hbh5VYVIJfU4PeNndIJINZGmon51EkXyCl8vRxMNgxO3MFcRQuSiaEHZQ3B+7KFh
WVDaKKH2zJ7e7V+zmHYHC7ljtwGJVfze854ssKUMCnk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32800)
o6r5OzYX3ozbkheyoJw0PpzgNK5jBooGnuOAmlgp0boBoP1dXgCJuMcf2bQU/3N6
rdYgLeCrKNhCocJ1reX9Sx/F7od9srKwL94VP9P459UKFB1AEJ4RieEUZEhIXiau
C36IutV1OHlvSPuRBqBdMRGjn132hEt1fEZwBJ7yj+n1Zp8hhLqal6DbLINHOvFT
u4ZtZSQ5UX9bTZ5f2oo4fCiDHXQpkYK6v4ML3mZS+CcxDtM2jcDw0qDqcYDl5ILe
N8su5lmdNKCJ/scCAD/a5RHV572iI++Tk8DXOpvDO0YXY7/sUnc510vJd3eKleJ+
SExmnP8Eu7MxgOYyBhxZ6oLWuq4eQg0oC405uvfdAxLeqSTrQmrYl6TDuZ0XrOAD
orHFyi81v3UI4A3OMjMxFX8PT9zS9Fd0fgJ9qf25BFBAyI7Hjg/MnW06gXuT+zIU
EUk6KibnC7Lm8qgl4oGpGoWYZenzdGnJmJhUc/shc3HicIB/kzwJLk3TJu5AASR2
e0LwfpH5nfQ1srUyHRg15Suq/V55MWa9HS44imppGH0xf3prYLL4RGwVtXjcJ0kv
ufRe3VVk2gRXDXNi0vrpep7zjMl7uixX/MiQDl0l6ZRmkVY5R+qNOl9hrqPCycSR
jebwRt/9DJXbgBqlN3SBUtHCe8S3iLfTgouq1bUtJl6Wzouk6oLhyOmA25W7R4L3
E3imdm1wfFxl3eXNq9YifwDY6a+WIJGN+jAKfJXzNOZCS8LuNR2Ae8XhgHFVaxwQ
5Zyp/iH06ZB5wy+/fC29DBNuDtwLIkCHhpPhXjpADqtm21NW46nDt8424xJTwUFJ
XFNEyO+SrfCqjbWrJAejK9FI/VmKW5GyELegeS0T97Z4DG72GkBrN4YosS+3PaME
bhZLQwTQ8yVbIciGCtlP3kUX7QZ9GvAyYEtEWWpXnx7IA6a0n+FKph9FKxHsboOQ
52G1EUNdl134dPDupk0RkygchrOMGkk61B455jum/L3v/oldBwjI3CzV630RnMEW
Cya1wL+3/JraAIATJPrQ2niK/KaxpELzo912e9+t5JSQ4j0rUk8K2dR4DaQIQb6E
/78VmTa/3H2RnWya+fDxaKYeSRywI3o0l9f0Im60LsH1TbaE4cLO2lUjDhLj/Jt6
bm2Cg0DDGbirctYr8d6Y4K6W6S663H3RRDypp/ci3Cp7wZ889cXthkoFe/elfOzO
cfxdDgRKbKeE0qzcitsyqb1sP3nTeR9xLDlKGc281s4XnDvbA3pueXDy6OlMcDhF
wdwGRFg/+2yw00l6DMb/K9zWXdhGNQbalR9ibMGoYyGTc/7QKLfiPjSU3zT6wLQl
rLUBQHzKdO7c8qgmOu1vh/kIy2DunPYTL+0YuYASUCSXeeVwGWm52PDyI5KJQoJQ
IXEbWZVDLlLCHxSDIyTwM5GqqIAMZrBQFTaBJ4dTaqFRk4cN7SN/WpZRMUuqRgB0
3dDSpJ4kMiRWCVSkL5f+9ILDh05APAK0CUYD7lxcimCJ03AwLQukCX6mDnDYD8BG
u64jLFuwL3m89oiJthy/WyaQC7lym4GuqMtgvy959gyMKfyEkAv8XNclxnCxP2MQ
BU0Y1bYizvWPaWVk3LdR84h5M/kdgdG9MJ9yo/N3KIHsORmmnLpBsLH2Bl7YyVxc
XcJMRI4OWt/B8LyU42L7z6VO0Q2s2LejsUiKBzHG/YnqIQ+eCAYDXl0hj2uVKd1D
rXN4fuOND8ZBwyHRUZP32t6q3dEaC3QP7rVMovv0oe5C8UL4sd0ctTdprb+pEgy7
iu38WWbFVNHj4oi6eBBlDlKkPVw1fCyR/O8s+Er9aa9oFNXpBUFKhOve5QvZIaiH
op3U0WUYhWxxtU9yBZp1Dq7ZO0uiqgwGJ5BtzVX9v8HTGl9t22DN0osNMrnTmPWo
Igy4m6YZ579eYq8Dyeb7C9+Y7RtPd3ntzNL55pRQ+TGGg8+CnZbTcJbVNW/tk2cc
h4eUdulZv0/7H6pV06FarSQBXS8mxgLQVvNJ3QX6k28sxl5Kc5Q3XYjl4+Ujodh9
L0W4Q/qoWn0tg+ay8QTHE1uUvx2QSYkp5Z3Rsw3H4nfXSMCk9qjeGD1cW4oEHm/m
SU8UWPWe9kpyU/FD+P9gpyUefirZc4hDB0pp4H/SSHGUm3B/LZ1yjQByfpaMGT2j
qE9wgHKktl7zISceQyX79tNnoaqxk0O6iwfdwFIGU3nLBMJ4i1XFbMMyanjqOgPG
h7RxMF/n0qQk/nailp2aDfK9F1xqh2LcMFTvdeiBez0tHUZ7mGX+88FR+gi5RF5A
+752JPkcYMq2Fagbh1Uxh4j/TRbsEWZmvNVCzLpgtuzD/PW/+rLMFUTA0qPza0UE
d41hRbrN/ab8Hw/JV2SvIzafKL9HwguNALL800zT7yZgHRNn/wIGax/iSWr+j8F6
prqemZD3whE9liQf9e7X57s613jPnwRIys/GwJiOP05nPmRmLnNsINXvpnZVgai8
wfpvKQDJj99fWU7AGC9kfZRUos5VJP0oY4m07WgSw0EWywKQ9z8HZssA1EuKhQz+
WYdYJkKcEdE7VtrBfrN530j9j4xaoDJJnSdCiu6NDSgj5eAzzUjN8rbWZEqb0/5H
7Vx8gjh/8V+d7ZEatPR3mlodiFDYXxUeHS+X7fnKH0eMzrNBuINrXQcpQ78cI16H
WEhMJyQyUJRlcJonqoEDwORsnGnJmEPPD3PuyhGBr7V0/2YdeNSZQKKZbGGFRbno
eGkpAHP4XJ5zkzaCtTQXwQ/d+K5LVvMJdrsCzjs4XH3eMbDOuvb36AJVGTrS4JSl
HmJPHZFpp1A0H/1l78bHEorq7CDAI9/q6J12uLwqz+bmyNb0EOV0b45ggLMdMedM
xay0gGweZaR0FtS3MrmUq8sbalYvmqgcbjnYtmYbOvXqX3jW5K9bU00a8/DNu1G0
cRZq6QQdHY/ygksLpMX08wBGfw0UwfSbABtsJkLl3FPSxGG/QyJlvpxBCornBTV1
rKiEVpVOy+9p6oua332vqGJXwmhrqY/Vrg2eiDmZEYS50tinI/6kJrovQlFJVI/B
a1m75lucaxgPIfYOqXFiy/jtJFpdE6aXQe9FACOo+IfH2h2XwmNHP0h9aVCUnUWD
p2jI9qEBl4RNifk69hKLv4x/nl9aQefldD1ltdd+gcnonUuZl5o46j9Oty8DEt/G
T8P9yC1pX25q5Mu51K1iRrP7YVeW7GT/+IblDF6AUJUIrFs/nECX7g5uvqJ7XZx7
UJJRfgJY5E9u7GPpYW+TzGBGkpvIHdNfwtF5a7+0aNOXtbhbYTT0ZA9A2oXhLwg7
OsegwZJDq06oM3mBFK+NqQJIcDanowJbEXxuyEZCOLH/hUCga50pUoV0qH+j8LBm
jtgNR62Q/neJx5t6eiNR/S2QOimrNX3BNOIAcdPlMgekNuMoRNvfihRgihu+wu1o
jQ1V24DKmhmIU0Y0RF+GaeAFhccZtMnhz+2fExnu/A6ImiI/XRJl7BdCgJvxcHHa
6/9bFeKo6VH2UocEh1PxLJXt/q3jt6AcB/LPqJmHo1KBiedy2UCSdyu58j8gtQWD
tMDtNBtkR3zwdNzZnT8PMrnVKMKSwgyxqKWBrD84Dhsptqi6y5ZhvXMRoRyjewOq
zUBDfPppZlTG6B1Z53T2/hQHwcNCQAe+GTReMmYD6szZyVYz8pnXXlzkn20vwR7K
AKKQoRaGC7W8dYJLiFg3dZCHz8tLAbo+yk72dOGBW5Uc6gR3V/9PVOCQNUr1CtIN
yeGI+FVJv//rWeDJy0YQpp9E2C09VxVkLH/lQky7AjrErZE2BZKyqDEUTF50ONPC
DdCOgwi56pGirmNtypofR72m2/HfpOUDDn5/sgOfYq360L+iQ7mrtd7BO7C5ofGw
RgdPF1TLeE5fhztZSOdtEejGIb8NRFItG2if9j0t8zGUtVRc/VGzY3h1BLKizfq+
bDDH4wqug/1w3W893nJajLC82sWKwVdaprZTTmISiv3zb71A6fD3EHjqzstmdnKY
CHk3veuRHNQvgZNdX4v/dNplJAA3gOdGK+dv93IPxdHzeN/4bEU2jZ8qCJKmY7wY
j7P6uk3b4nAJpCCOGWuqFrJUQwlLRxfae2obGNfOTLCMj6aC6tgz9Ec+XtQcfgaP
QuI8KO4uwHmY0hFpFRoXvrVSdEcTY9nL1Ez9azsZvM80ZS5F0yMnia3uAFJsSMN+
IzwO6pH9wm/gVG/kMaiARarVw5gBiN0EAGCPJKAHdYQJIXCRFpEJeq6c1rj0Q3s+
3MDsNIfDMPiHzWAPKmtEvjWlnbxmKWGjM975118txCQLtwtOk+RtNpSQHOJ44Mpg
gn9/bzNBep8XB7mapYgIljswh8DmFGxHQCHLr8XPojpg6B6JgWWoTFs8CgBUP2SO
benQDfdwLCXp72TxcOhnHFnleyvq8TtY/uVXUU2epBc9TQzjaNgB2U9wRtIwHrRy
E0ke9N17uhnns6TUrsQ3N0+NlS3lwA+WPUfv8dtwsheaMsbt13o6S0UO9hLSOXbu
63SuL0McVwgZbudXHbHvmjY8xOy92EEVAvEsanL8PPj+DETi/LolddCUKTJvsbNR
AKOB5hK4RMYAkamcd5Lebf/R37mjV9CI1juP49fkRCW2tWUF8FlrSzV19niI4Rzs
k2eZjXCR/A1SY0GMxDwD3T72XcRmsLuNjxRAf2xBmTz5+K7pZk04mkiW8SzngT2l
4yryHA1xCFjNUuXRkFn8Y54Yv/JarW2qkNb/ytpDRZhnYlfYlcoHDoOZct0qB1xb
Vq1BV+hITw3fcsz57/rZT0aaL2+vy88h6Mw0OFwYwyj1rTUhrrB80OS0ZMOrAn7k
cOnChTig+qzRneRZb9uKKEhM8ppb9WZ6l/LnDgU64YvrTfdNl1yePlL+0auOE1V6
4wSqSY0VTI/Q22ae3x9tQ5xnHeU7ToV4EhKCOuq5fz3gpoQ14/06qmxExznAl5PA
8Gp3/j9K6ujVYeDidRkPR8TiX96B/Yzbl7PKZPxQWUKRdjSAlmFji3EzLyKzwV0y
CNMjyXzk/svuGeh5f6pfS9Dic/8GuZnPjJFDv2RALyERKCPBxyMBNnzuT0KUzWGY
oxSmsRpAT/KjTiXIuZkyJit11o50i3x2FjDp2ziX7svzWfxKEXpKUXYJA0FcpEZo
QhEOjUCKK1PLT7MYEfopFqQhfFWhfVVkD+NH83TB8pMdJrkgtvmYE+vzU8tjjECv
Gn1lfIrRKQbLYry6NKrICYbDJK80DBKaiDUHONkB+s6NMqVjGp+fqN77/nSIPC+R
0PDSr2biXH0PevW4L5B+25MDDLKc9+XyJUKwr7l8iiD31QqWh5T7B770Yd3skTdS
iv9mBZrbRU8tzLdwP2pn2UjUpuD5yV5PQpS0UtxWlXfvdZPNimIz1O37Y6/+Lrwd
ZytISLGY6Rc+XKsaF5Xbn8Aj2W4MJEsNy6t8oqt9fYVQoeBm5VTA4EI5tlYOIL7T
X4K34MtCQ9l5uhceic9BQgW1t5I1++SWMpQSK5mcEgxR7B3Klh+tyWGqLhrG+MT3
rvphwVwHgHLR5fI7dtARBKGL14xOmsbSnHZAHMeKuK7Y2qyHIE5P5GV9g3kwpAzP
CHRbFWGpXFuahenGgD5f0+kE9eEx/pDKsq1iJynJUGVZKgN56JGusPuJ/97q8Wly
jSd7X1n4SKeskWNboBHiFSsQgPnAhrsRQGfQCvc6fzMhjP+WLn/EKMM9LFx5RkJc
4IORLLLhS/m4fW4czZfDTWNZZ4a+8I/DaUr80MEl9wRptBfjbTS36nwhZlnQ51kR
LWRIyM6hPkgoHfhGZjl9h6VX+Pk9TdLdbhwdBZh2FsFlacrdKDqkXKXjCzhzltN2
uU6OSSf/lVYe3UT/tQFn3PdJNjccQr5FarqtMrNpdqoTzVajwHwCiJELF15FZyue
ubKFwHM7IbebEx61W8Eb8aMYVU8ZvdnWq5/iUbmGtcinssM/gB/5IPif02stoYVe
qb12QJGK7rxGynCGIjgJU/0bwAl3kN8bNiGxfHQLqtnyD5IHjNRe9iE5L5j+01zw
GI4252aBj7JueaUMqZsdMoPQSZyQQ3bXb3kCoZIn677/1M1C/QfkGRDGWg06HDeb
oJwhGT+Ssqn8a+viWnlq5V97uvadZl2WVCQWQzfIY1MuW52oa1n8jqEEVNSe/o9S
zYABQ97qeZkBf4Z/mAYjcuacRImDCiuI2pyVfPGptBl50MbbScFTYiQernuf5wJv
MYQ62OSSQfDW1VhawVqc+uW85OGEbEFo0eA0xdmQd5fHZBR/kl1/IO3+xaY9VmpT
uR2it14wEjT2jzzHsC/cgo1BgCDCWTzNNc72lDVX7WxeiYyHnkLRBC1DGWYDIgNx
Rl6UtIFCUfQofbPG1AhwYFiwRyw40YPEYqj9pTOJisgEiwgS2TkPb22PCIhJfdUA
vLqHDZ8+47rUEGRgUbxRQlSJ3R90lb36gSsHDwVO0yFR1y27dEbvZ/AqHRZ5woJU
7mXFAZ8VaS/122q+q3KYOSF1DsiknCmlu6/EpCABnRF25W0m4E0fRiXq0/CCA9MU
k9H6yruJmIPys0JmaABRyjAO3mbH1MYmh2Z0Jc3y+wQgeaTf8DT9+u0/MfloZpTZ
b5cyCZNb8KTld1wcrCuQzLmm27+cfm03EKSyu/R/LoiCvvTzaTxWWqLiFxfyj64F
l0I67Qy8mFyOI449HL9JDFj+TJrkImg+wG4tl8CLAfM7WSGBucaIPzjOoO0lJnAI
JdSTfA+lcXX9jHdgo56IkGouHe2iy1JHRpJg2pxmGI9PGGygZGNthxix/qLjH746
Br4XpWhe7H5z6JCA7k8Anf0058LzvrBublFtK3gZsStmulL5IQ40lxL+OS9QVAI7
d5gMtiJzlwSn+xmxLqSnOqBAb198IVtZUNIfPVkYNM1zWzb7UqiKdX3IVoYxjxyF
z0f5GxePZSOTQdsTyqXfoQe5IZRAuoaOsCUUpsYk8PvD9bxxDjNWp0TCjp1KtjX5
572hHTUuMvrQHxmzh79cahNpU/Ozr7yN3/Kl9ObTb5ffNnRa5HN65NMnwRyYTMo2
Dltv9YtQoLwlQG7L+QEw3QyCgLjf3Ny12o6uEWJyh+WIomar/WcZuRJuMOy7i8Zr
hJk3Wb8jfKL2bvFRc6XDfoYmDISE0HzOxPROwSxMnf2LiN77lnsDuRrFOOVqbzVu
jbtEzQIBRyXNmiDHXFcHX8WXhY1s6dZuyCsprTAigzl4szKr1Kfrv0qfg8h3GZgE
hRwGZCMhhGRqx+3hiY44hLvrdQzf5TzmecaTdJQWYe9RTG+WcMzSDAT2MRjurMqB
Psc6Nc/cwTbkmG0jd3yCzNUpt26OyyV/xTSuJU2NGCPO35br5v9uqQfJPP7p3P2q
CXqfM/URY5sTbb3/HsvCqcb/v52hMtIAmB+oJf6Hxs791r0QyDLqR/50Ruo87JRg
t7HZU78iEgHH+oTsDDjlbyyH+DENst8VsGWhzqRX6l9s5GIY08AG/LBY/oL7C1MX
R0hDbIPYLAkTr1kX56kNmdfLOYP8JwYFxif1luvN3cGW9/JpvmPZ0BgkWUTrwb5P
WCgTwa3SBtJg34WinsES1reWHBpkvmDeH35/Jb7Gxlpq3D8pXMr2RJteTuxssmpl
SH5RQDKjDrNBejN+8aupTNrqUrAX3Gf75J8hs9VrIpDpWGXjhz9/9TYd9fny0Pwr
7Hzro/BC6VjaFeS3xI3KsyZcCedzpMO1qAyzM2tF76MmWAoeDyyo3j7uUHmB+vUo
+ykFLYJmAY3kKR5yiQ5KRx0X8hR15b7T9e7KDJJgHzKWpGWSrxp1uFIH9EZSccbz
tnctgcyiWcPZ2irMFkmvZB5bZaawdSO7hLc7j1OqY2ySN1/fexWZR5ygUElc6KfC
FN2Uhp9iThuoSl+Kpvl1ZbMZrvKIU70h+KGGl4KXM3NojiQJ/OxJjz3xHq3figbT
lUsDTX+TCjtiZGxGJRzB/PCinPMa1L0OAXDEkJVDpPFoxbmE6avMA1vc7uRtZeTC
L9EnwmusV/GoYgxAfck/VlgqDk8jVrHL1lr25u5D1dTEZvGXYc8f1MDdbcEud9Uk
9vbXwi6UWt2qmM2gIeLMUT4ucimCrjos2cRH/1qNHw9g0zhmXyoq1ubZQx/5jtwQ
rUE7JleqqknXFsRu/wmVwFH/cnshOGYw6kfnlvIk9tI6OIOYhDRAMZ7dZGCEuT/Q
ZgKeYMQT01rF5GuC6zi6+c5JLnp7y0Lvrcpe2O15xAxx2bO4Am5JiALdJBjlAYZT
0jzPf8u3f+1pgG5FYlzYbzGBFjHgk5W+93N+n4H1U/g8CoFhC1q0MgrohzIeUt5F
pMQF2IBZ3IjpyeqxE23BcYKqDzf8DOuDdrbc+ZMt4Kvg6PpwkPjYAyJkD3X3NtW2
SBMdLwIxU4JgCJHGYB93PHE+0K+OpFQAVtCmU6b2b4C0uyk+IDVhv3WXj2G4LJeY
EeBEEIy3LHNaeu/r33zjWNQHPz+tlzEuq8dU6JWPEg2UrrB3/vshCxghhimwcz7Z
w+zrrYdpjMC3j17iFE135FzHMB6RwcSmDS+cqU+Zu0dMNPgIAwixOJtCqC/v472J
ZAEabc9/G4VqiZfyh5Pv4kLxQDk7eMP4yXIF/uUMRehlleUtoo8W/GU96JUyym+9
Bqdt2aMeO/IL62ksaFla7VNhOxsvl3a7BOtr8rqV/dtgSkA+A7wieeI8ZCObjSlc
O9NE9PR71YYY+bjOVqfPoh/dOYqGybhbiK9mzgsXdGC/hm+uCEhRk0kbiu3N+A9m
cpYZvytaY8x5v+QRuBxxYy+GO+bGozu4bfBxL4wtiJu5gjRPLL2fnBFZ/CBG2N6P
lt8ifOcNxVVkvPtR4ty+IRE/HN5jEx2rXJRsUX5YCzRex4aDgic+vxhn2EaNs7tL
MdfsfTrEpnETiKGAAI8X5+BDeXzY5qrvKW8dMRznBRJ2tn2+Py4nfg8NEruLtOp2
Y3lu66D2t/UU7iG0kH7PAFWjd2/t8xJyOjdTwtm+Mu39Qewf/oNYWT6uk2vGq68i
hbR3R6NHJemGv00kS5XFEbm+2Y/nlQjKDbBCSMIXrXPrO8I556uucqV2GB8j4Rxy
usFjHLSbnJGgLUrVZ0JDCY/oNUtjfaj5ryl3/p7X+dTVJaKMBGFsapIwgWMFQK45
/3WmyeVEqCV2PWJysMA7xnkSLOBgQds/j+2zbCjp24rcs0LAG00jxucG2IIuq4xM
Cc0pGoOCLqBwipWlcXxsjgFtbRP8vS77AFhM2mFugOA8gvZRTrtkl8h6aUKAGIQy
HbjzavyHiMv5AMWS9gbKXDvGBeeNau0ly35/lW+QJ5Z/AKuRXRdqTH+/5zjcrHKX
4bApik99p0EeY6pv5w7WdhiteoAHyWhG1sdkbCfH3mtmehL+Rvw91eOToeEVo2sz
nPeUYyBwv7sfTNI5a8pT/QbyFhynoYaGg17ukFV+2d3CFW55NIOgSX7uENd626wO
66nk3yFZDsi+xpsAxel36gZ5S68fOe3z+DUzKc/klyO5CXADZIt34dUNWExiLwTR
xv6+SFr6VzCY2I6vz07IwoY4sJ83xTJPbxysD1eYUkG/m2KeczIHHC4EQ3KvMual
waXsRNKmIs1WzT+lcm3gi2POOjA7+HcikVHFovZkJdxZtQDLfKnm/NTNym7gBVMZ
9YEu0Mve2wx49u339Z9y8m+iuOnnTO79/4p3xoRSLM9YJKL7TJdNr9nZvAwiSJeJ
8YodBXmLB0KtncoOhXBORY8TZZm0G9+44olKkjF+bJJfm61gV/hmGXHH2C5LDcrF
shys0iHT4lYL8w1p074ujaRZdOJ07DRB2LceMTsLBjEMEbwIJpNNmFIc1tiESDKA
+P5HyQ7WteBCubPgBi+GxxIkhnuvyLrwl9YsBEuc8Iy71c1zUtkU0I3BtQyaQcHt
w/GXVtdeK0z1K7hcrM2TKXYmDi1hTTeeKKgRCmfVXhBKjt/ZdBRa5T+tV0cWigf3
t93d7FEV1CKWS0mXjZU9ugYQovkRsaJa3S0W28d2lR1S2YT2ki2GSACKeux+1DCs
r7kX0VtlQTxHKreH9k+z3ne8baekptVsSe9Mzi4QmHMdMMcVflAlEPUkkG+QYiGJ
BFs7NR1MlY//1zuQNCxjwNQP2JAvSR5+o22YjEcj/loNrkLMoeGcjbzG86J7utEg
28LBALnaHIGc+tcSXcZN/fi1KCbi17Lj3VlhJ24Zw1fw+b3RnYNT9e/Ftnv1CsvL
ql8+4NeTkzh/YKqD5OTKYWKnEYwCcxdscUD//Ue2qPsatWr8kA4EQvPO8a9nipvr
MCmd2iJCS/IqamcxB/UTPlvfp76wthzwiPnVeY2C2h6w2t9/1MLsJG5F1grr6rhr
zdri7453tnWfbW+//Nv9a7Dq6p6gbPcfOhMqXDzA+ZMNIbEgu6XyXh25EWhxR56U
Lam3iGv3Ox9qJFgKl2v0h4G0BZ/v7w9flU9ZUIf2N5oeI+Wef1iICVXyRC8Biimq
Lev4PGMgBV0gChsvSAeKLB9G7Tw/CdoPdBo6fuDDWS9ACX0gq49ggA9O3wuL8OAA
+t9B9wjMYnFdAlXywbBriryo+cU2L5jxsfZXshREyLYp7g4JuXHNOueyHCaIL/Ox
no0DR6eJsj0ZfGtVlmcknOAaADJ37nk+MkBQl8eIwSEMn9IHIOKWDpaFWoZBE6j1
HyF2yVnqLHaNRsdjHhdox6Z81pihrPaLiysVHgEnuC3sVjysMZ/iQKl4dpVQblu0
jcqT8EBFW0yPLjw42Or65/iQU2BFdpl/hcshUo6MwQdRhNZUzoJl0F7klS4qAZjR
WXqlH/t/XQCb6lw3oxHm+68X49ifnfNEuk2Mb1CykP2JcZv7tyCxbtkU4iKHhoHZ
G09dHXTk27pSWoe7D/FFE/5kO5pKIvEm7J3Wg6oBslHmzGR3pqmU0mg2J2QCoIYF
TWsPzlmzzJfllVARiEfE1YTf/3GOOGkjr7RlspH4wupCnrjIYGoyJipxCAIMjA+J
dpCBtHD9f+5yz74XZnMkLw1+VGxDCWfJOwKQxjVMzXgiETx1bk6Li02f0NQDcxtV
Z0W54rlykCyqlUZQwWnh9E1S7i7QIUXPh90ruUSli0N4jvmeMEoSyn9u1OQ4AzUJ
RGGqOoc+sqXnmZ1g1Or/I6QuB7wnz2sityfrKbjoEjJoYNXd+iMERAcnmzhxxU+4
FiUHCqRJiEHgErOfwoXy2iKJA3JIHwi8y5sCyQr6AZTtkUHLBEjcTc3ehWrlFSvu
3rdrmtZvVxzdMNg6PrA5z7cb4fvt5/tsMs3raqvTDHD6qjY8n3zqWvv3CvUPSeT7
Owy5d8OIhZ2RxRBQwQ8+p6/JRohRb00ZAl0twURGft4Tx6xmhwaTD/bruDQWbP1r
7BqFOvJ25WPxXgjo7t1IX8DIqbFploixExRfVoBObRtx0iHrzXFgwIfu9KaM6Ar7
/bjFvbWFLZVk1GrQNQHp7sfvSsyxvNuV5Mv4iAgG5kQG6ntt3fuM62YgOJB3WZTj
+CfCZvkbHzf8vHXx0C4SCzj6VEFXAtdu+IualCIvPd7+aQ7dTkaLJol+REwpsR02
+2HGct4oZgQkwzTxlCx1EvKkJrfm8BiXsEowTeL03TXnHYEaqrNpCbVA8D5QK/cw
FYTwg4iyUdZifcnUISA4y20L4CdsvRxhVoQLQZfu/D1PxFOmU0CXqQQ46jjlf85o
jrk/X6ZEHp/k8I/6ULwoG3TUDh6Tw22B+Aa+8Kv5i+voM4EvvXSJUSIg1I6qeV08
FFnaeB1KAkqAlkDtaqfv1sKvUC7kw/2RT19QDgYxzipESgtAllXU3P8CAJTUuOze
TlYlwKN6IkR+/9rz4QNMH3LR8Em8Wwe519ZhCvntEUu5TP3sgSkPGMbXve7N+MEQ
y6mUQr7l6wcUB9RrEgV7u6FD7WnqJHq92KTFzdarjmbaziO8XMUeUoh8V1ZBVWp7
Vd4dQrgjnphjbwj0WA3M/Ib3G0q0FRvsM256dNjfVIPlN524TQ/2kv6+OjMrmTxA
lSaqI3uajUom6JZ9KPUJM/USmG4QgSNx/E8qxVSdesH19L6Gl+EZiDnj7MRPq+mF
p3h9UJMQD9xQiS92Fzj5jXRT8VUl6LRyvZpmRtxGO7K8z21q0/uQhJS2MrBOKl70
mOLWhWP09jS7Zs0gmqxG8QmqQCG5ckQG97s6YL9+nBdbjerauD1or8aDUgAI0FcN
NsrED0RhK+KtWgVRd2o3D5XOgx9lp2Q0sFg/egEEifNLGRdAyCQs9K2E23ZYcv3z
E51hjgjzKPDlzJGYZoum7/iCQrNlefxGPm7JW4Wr12s3hAIA/jALwbXB3bQ5u4ig
QEFa7zTLS0ZCq0rlm74iqGSKyW0HNrwgAOPRy9Ln77N0Kyb64fQlUZscFAM6MYWx
DCG++lWb9W5y/O+FmCpGPbng1+7hA7Xmt5pGw1e6wEhTckFJ5ge4zHfI2/RweYoD
ZPpVsfaddJW5GGHSBYZxkZ1xTxqUaDJH7rb6OuUa4lOzPmM48em9uNp78Ivgg6KO
HwGsGTtRnXWX2R1L6SVkrTU8TjWRyYpaqKtsR/uaYI2k4sh07W5+y3Zuodb5JVjq
gdQviQtX+tnP6J4U0YAuTDaypAmgT0j1d4PV4zqEC4E9lQZ5Yne4ua3vj+g0jshP
X5/ryBUmahbw4lNm6Rv0ZdN8VnawrlhQ6TCNOz18DJzNj7aEMdhnmuV8IFQlQAxh
a22KhhaKoekYldfmQlQHXyBDRthvVdWaASGkUr1rHzx0MtcYU6EfsFepwpAc+33b
il6YtrmwJ1Dt0zjrdYmkmJk99zSLi5Mzd0QiTFlj2x7ldfQDgQvNT/fY4P+oSJl6
zsRj6BA/qZLrjG0gzgxImK/OKWbr8ON1HnkuIxSRuzX6w3NQH8p166wm1ZlWZcr1
iziBxImpfS3d1sVIlfqR/IMFZDAIWTjMy5bRw9sSmbYGPN3cNER1wll9B3WueE8l
Kua3yMI+QVMPYXC3kYfnvQSvFiDTN7DsQWcG2iN91SHfK0wZL1ac7/AWJ5yXz/iI
owKJaMRLcBIZR6Ru+pAM9IaCEJknSfh+Le+M5aVTelmHwJhFgJiCWYd/1bgt9zK4
Dor5APu3jAgbn/hCKsLcqVoIhWxJfiRUf/EdUBM6WVVcFL30/JOxtSWT7VdmmoJi
keivaQypa6bupzjsP/IDexnozbbGVbjK/4bAiCMOynHnPPWQOGYLWnmBUxav7Z3Y
gWcppk9TF2dubndlhNs02zo4nyG/qxh3MQHxqoL5EUPPtOzN6EWay31t9O9FPqXR
mFQx+6WlO5Fx02/fJzo3RgfuOoavQqwiRYp4u1N0NgT7NX/4RcWe1RAq+xNeUX9L
5sHaJpHNDLc12hw8toMaW8O1AwmFSG3g6yd6a3s67cO3h9eKNs8+/IL/pTHif1z+
X0P0rD5aVQw/ajRa1bxu42WB8NnmsBbCiKirgkiBO5V8XWm4T+jeS9QDj9mrinF5
mgqOXaeavmsliyaK0F49SRD2+LzZr25lXiBYsG/e8a3SVI7r39vveAdZMjI9hGRT
fO8MgKS9R+x03ily9X6j2EVoFM9MYFe7/TCmiULe2bXamDO4y1cF+3Bf8A8DZgVp
FcJ07dULIAaufi4tcoDxj1qEF8Uso7vNSbNrsOOD3V9/GbRa/GqlihTEYtZ16Jl9
yRXI0opdn9MxdJ4vxovu1Pv6LcDkPngksI69LwcN1fWuhVw5mBakZzjjW8/7ww5R
flplehj3tNNjpb4s3X0wVAcyGtsWQ97dZPbD0V15f7dc+S+NzJHL8fuMYfGVFVDe
D0GP6lOkILj9J8GRfwuHp/vJRnlr/mk6m1Q2eyHk1ePw1ip0gb/ReL9MDaGvhbi3
0kSI3dRMnMFI8Fc4l3QrbXVZe+4rLknEkLGgis4dCUjzvt1ESOgzdgW+CvlXkwNe
jNgNvL8s6ayDbMfEN+uWOkZb729hd8ecTONgVWryuewXUBYw/O+y0MSeXAhq1GG5
jzIe/P/Vd7N/1fLoB6loe6PiRo4qe5dc2qPXmPwONg4ET9DKnBsEMGQd6G9EeaOZ
eX7QcXnBW2CrsrRMna4LgOwBCg2NAzyPHh93aQWi1RjZHOTOmjH238M2s541mUYk
XnbtfG1K6ImrC/cENNvDlEcmy+8Sbmu0Oouhewj85ypBGL9mgxhZc8R8SpFGHSoE
reS8ENlB2Neoq20kjGp21cCva4WZ2oABSQ8Cjbd74wdm2rWrMclGYyWUoRiZg/O4
1jmF1PtGRab1r5UaGTgR/OdKCoklP/2+P2Uwd+iUyxjq0lncv9cgK3NVsEuaNH/X
+Kwm4kN8i/tnHuZp8IPx0N8iGvuE8gANHJ5bOWSBiqR0j7nu2UeQDG0TJRhhKvoT
ydwE+A3qk3qQmgCjazBcRRhwTBaBAk2YrMWOx8OzmcZNk91oWIieYHjC6JRiaAmg
e2/6CS7hLdzGBulf1MMja9xM10APTvOwAo7FKqOFTLIftpi11tV9r8fkGuqkgq4F
aeol/TeRPA/FYtUASs280irkZY53wyyJ4qDv+1S9rlDE+xOxVAp9GjnRLGo6DnEX
hWiKzQCl6CKPsI+VgfTfIpenbiH8hNx8Z5tmgRG8MhuutMJ2fgT2zOcGc3XS+v/t
IqC3cqYDtzHuXvBuSUzpyiW3pWJHgc+QksuaxWhlyOUQQnxF4kgOdzPhH/U2lrIQ
7pkmFGCdn8YAAyyJ9Q8UHcJXqkazud6NEOBfHf5tk3FQvGM4ceeaeG9eP0A1ZLXh
+BM+qrEzdbOErs52D9wE6sy+PJ5q1JNeHkBehkCY4OTrzkrE0yPGz4W1n4PmYmka
lxO49OJYmkdPXZFalRv60FnI4S7mbZx3fVAR7mowjKwB8POFogiKq/AV7EkH3tWf
wxHSgfqm0hfGljZPpk291eWvs0O/JUwv6wSPXhtywyc1BK8h5b3Z6hDk4IxcdiEX
NCFAig1Z3YJBmliyDqQbFi8QMJG4xGML5vK+9kDtDS3lPIH4w8G641bwhxMhlYvI
xOAfJjfjZsGwrEjD3BiTn/ca8Xx9A9y7xSF2PjTkAjbARTTQC89y5St0zRC2W54q
mt5lsHJmR8f1wbL7mac6NEbpmOtcs+yzvG7A1ScuBSf7m0Es42Y7oPIDYNtiVmy9
achiL7v8SIfW4aN+LpnwcDJeLD+xy/oVpJHqB28KyZnHpVDiqhyPTAJly5z5q4Jy
wBnX2wXmWcKaxop0gEPhm7nPxgJ7EZZx4Vo4KT3UR0D0Kx4u37q1I9oN/k66cvFm
HU1xpn3pJobNCvsGiCJPeUTzgg2q1gNoIWxm6xGNHWQ9ld7WGlehLN3DGB5qp5KY
Z0070Kam2oKDuUK/DzK/1MakBs4fvKjraIBPawn+HsLfheY3Ck/xxKK+IXLhsraz
Qt1Mmm0STjNdjysaTOBX/RmsEzMLY8jGiPwpBk4OVYVoJL353Cxj/M1OBr2icFZy
xDkYbp98m3sbkSsB4tOfRtiUlrLBk3P6fMPyz81/qrGAyg5x2TZS3YU0YprwA9ca
dlnWn04zrLUmEtb84h//KERRJcA6qQOWu5C7wT1aDT7amtcsc6gDovJUWtaTEbWN
jqQCmihD/kFlWFNCAPSm4QUY7hTmaRGIxtJ6pgos5iYSNWaKJXy5v2DYfjGx69eD
PQt5beq00/8EnCZmU/ME+ReaQxdqCQ6cIo9jUpyiEaTKcpNtT6iZOYiasKe1NxyA
Z6QMsJ+0yt61vdIKu06q4olHa2uu+oziemQD369RldxUZhYw0FOeVwf74R2nusTu
a3WFIQtli7MUE/qLtSJyvtlg9YAJTc9ZDcQrpUfC1GhwqXTPbHUJoQ9ValYqreg/
rOx5Y2vrARCkc6wghfUEZ8xA9bTlNXIfTz09uj35wQbtFMUUYIcMCiw2VC9YlhIC
aMYgQM+s4sP6hZV/wM6dIuZQcxW9M0V+JDLI7JnB25OiSDXJFWO1Z1yOuTuUVbbY
M8if7vK8lbbIoT+GIT/QcQXpDxZrf4sS/u+AEAKIwVzSHu0Xa/8KkqiukhmnOeie
RjvPFgiegDi5yietI9GQmBtzimWI2mrr/6TwKyi+G2jf/9ZbHDJOS4XKllqhZfIq
FiD4crJgQT3oOzd9rfKf5niP7Zuhj3UWNzqe98aYCL71Hwx6+wc1+JxC9AJm1Pbi
GjpfxtksH0qoS3RhtltS5GdxlWTOEQk0qofcnLaOy7uwSgYQQW//22kHJfqujO24
1TQXZMWf5nkIa5wodH64XhoUlDkrcD9ClZyqb8P06Ej+5hk2b6TGteVejk11cA+u
Bed0IZPDfFo9En+2eflYylcErIhrUoV13oAMhyUHlwRmXwS6IfP3oA19sVYQg3n6
lnyDHpao9MMWrWNgcPXksBsD1hL8DsCBqimmllSn6/cx6xy5ZyWeZ1QUciyid+RR
WU5gysgKqrvToMz4J/ZL8Rh4QOKn8diMPqGY+i3312WO0RWUoBNqXhOg5KB8WypI
LsKq7qxnaXEqjr0bnOIb1VYpB+IITC9twVbhOy5I94oajZpwOKlknkgdUQUlCtmG
jDKMARBPvb0WeKsG4SSxbpoH/daRwGBJ94ZO+450XqKJCTcaDyqOu8PG16rA8CXz
gp/rXriXhINwhEQwLhX6allKX7rBtl5p+QaLL63uLXwqrKeE7eusrRV3xxgVI5i/
ug6vC0QZ0m8M/WKNEmJDLVK5w4NdOUsHmgz8p/d6qlL9deQfPwXpFg9XKn3Dvi+/
U0u0LGy1XLPzovzfZv9xZGxr5ZZLFXXHw+x1L7B38lnmN9Au0AAHpZWWCMmcHSxb
+/8HKWCl2wvbITS6Ofsois+4W+W1DuVuGTtxMDUJh/BLGUtRWUZNhe3/hwfQB9gq
oz4NHMBf3y3aPFEKaVJOyemyLVIPZFfkW1uX8AvPFIKyhnTLK/GiQq2YXJFrl3uv
Pw3nmbEfqijqRHHeEJIO8D1xdFPhBljS+R6bZprrzNCUPtLk3b0hST/nyZSi8BFu
FhCEoFcLnENKXBJynqIP7uwI8pBy/YNKEVDCZYWZ5mSVMK4IJq8CiSOyv7aSHZVr
Q8uvssoZI6qs3qq/O2ZB3y6gM7sVpS6nZGQ0/ld4Rw4G5Znt8Xc8yQmvAzdgL2im
ncRfDH8N0V+4bRiCKmTU6LL+JgvcGf0rCltE4VtuDIgF9umWVENXvdE0Yc94hBjZ
UPHlIjSKogTucl3o2LsXF/pSORaUsu2qnNoXGlMIbWYx58HVQgQEdKOEyZk/1KXq
X4ijaqmuec16NXnChlKcs1My0uVmNS4OusR53sIMiDja6HcpXTYPss4WwYCtY6gG
mKrsB3bHGm1kV8fsPa5Ak+z5dfdv6iUKO+LOiZQmFWOVgpbBZIBpio5H909xjImo
ShideDrNfMVTIXXz9btY61kn0jqwAbjzF31Fv6OUiaOKr4wlnk+/Fce62b+eVNSC
sqsDyE/BbgCI1gP8rdediamekjDDA0zfOOEd9cqb1/o0r2blWIXLEm+xRMuWXEHs
WugyiX2Hbic2wBF7Ks5tb+GVWZvHq0zBBECXjdogiR3wU/c69Hsi4//hCnVke7qz
t4FAl71JYSGpq/gx23VRCsSKq61j6fR8M8F8vhbNeZy5H3WPRo1S/q5U9w1UPVbG
2My3WGq3IEZWFkObG4U4jQLcJVMTl7mxTcDog4D7Mg4Om3z5weZG4ZYS/eSzL9IC
Traddqfwe+qYGqNdmiasdNskBTQ5pGBNp0pb4uCVq+N/SNfHqS3KhxFCbhgb0Xfv
Ysed+/RvDxonpvcwH/g5QI+YeIpuqbj/ap1nJOZlBfRJ6ieHtjAhbILl0J0O3ewB
VLJBv08fVccPuZZTl4g6I1VGBQc40iqv2xz0xYft//54U+tQkuV3UvABHzteM2cx
WYig2xrzExfvQEwwJ2HQtjBgadM8g/24H1EY9plSLX5zURIZLglK0khuDIM5KPgd
KHA9/gCVjCtFNGhDtC+FRe7u1mDv/IzFUNI0A9OIy+ciZCoRTT8Qlz5O22Y/Zw8/
TtPt0yb5XG5I17zHy5HKVjYCVAJEew2Z1huGGvCT/xQy2ofmhiHQrN76enpKHNwv
oSWV9DxkJbbfon9J37c3QPUuLtHgpi1mY4o+k27owyqEmOx07kEKM2HnN8SqxxHl
nCO1AzFiBxPlemf10VzPvihQXe7DTDZOU1wa6eQqzKac172O+/fArlgCGE3J8KJt
aLnahWGYdXssZ/MC+zBzRIq8U90SUqvmdrbMa/4qzeoR8i09OilRiyXcbG2E+tp9
2Otpml7wATOYuQ9V+yR3ubBZRTuHTDFshMnYwq9MkaX1a82QwKCZzRVebWvzo0Li
BEXa3VxfKkAVp4TMJC9ne3kwKcB8tWaLzFPky/7zcC5VQIFSTur8T71HZe97/JyR
/0O2qPwLirn+jALEDGCDFzODzkyLm3iMo1wpc4qopEDvXFr8DpmA8qqtyo2GRTfJ
gsZyuJxaHJYPt6GlDt6YgydcRLB7mUNH++1lCaVn9r7oBwjqWDgcH96kHifW5Z9s
8XhgASRA5kF8YsY7jHNfP3X4hbdTk9EdmDCm8Fqy8c/0UsUgJ3gaNJHZhbD9htlV
WSdUpV6pdV+1B6OhWcT4mWi8lDMwfK2gRIWc+BUf2stGwS2PIuP/LZdRz9rpph0j
PQtpwKW4YknVkYONJtLkKoNzXKfj0GZhrnsB2Bdd/x/zDdN6oE8k8SAgNdq71rHo
+5tf39MxjC5U1syoqCKmwgMAQe7+bvJskgIXhw7XV2/sQiMShGcb5hLxQOatWiW9
Dcuag0mL4ezpzLlm78AiwCo/WZUA4Vpra3qhaKyiO5kvnaOz/Z02xx79dyjf/R/w
j5FzLSatCliqOGRjvNxsD0Bag0Z9MhAde+N277LaucXC6wQ4CW4P67cR4aV/uTxE
JrPnDLI9PGFsmOEvZ4wFX06QDqMCyz91T5Rv9WwPTobyuZRZArLaPCMRG2ctgCno
E5UjP97njzli1Jj+MIaqMAMNETe1rNpHZ5drInqi0fQQsptD9NGCh6s907svGpNh
gzClH1JvRW4cXlxc2IJ0lbEFKbq2PTPd7Geg8+yMzMJ97ITfBMg0r1FY4mF6o+GD
VfBerIoAEdtOPoLL8PM1bl5zqbQmGtQmR9GzIjdwP1lQHLlhp6ePrxOOfmtDVl8q
Erf5fDl2Ue+WdyaAn+KizxozxXYGPQLKxXcQ3yFVSs5d4Uho3MWWSOb7/kvU9I+D
DyjdUJkEsm6fUEP1c3dFto4AWURol3VtvT8XSNixeaD8pVWmTjBdFcUbffHQI0pb
kBjXkhT7/yOTIFchrDxPFj+Y736XbxqBToStacNrAD3OP04/7eZDaw/0goJVY81U
pym0l0MBx371yu+aM5nyM65vsvxjHSReOPx22ResuSTrv6iMYPSLk0Cqa+Cjqv4Q
A2JjcMHKU4aVGgKMUa1COWlaoa3k+nDV+TI1vgdnhMrr50jNRBJ6ncl7pdBnxzEr
TchTuM3dnW6ijfbOjUZbe8dovXePjkh91LFISAPw+RVJgO0rbp3l4MDBp8j4NVqA
N0YIQDKPQ188xDQnsA5TDRxTBVyzDAjLk6ljQXjtsRawz3LB+bMNXreXqx0+LpVQ
+6SDNg7pcJlZBzF1WqK1+QzD5+eyT3IxM0O5tv4xut3xkOndPb3L3JaDs+qFXfmq
7jSXpyvLxKmCo1cZQzJaL34of7P+a5CIdj3cvGd0vw0Uy0ktCRrWWqu0H79Ygsjj
mrtf/ioGEucxMB/Q9SqQo7Frz+fzQpAxrX+QgbGpWTEHyRyLj3O+/xQx7wN0XiMh
JQB79Ys64HG6dEaKeDDOBaCMrhKo5UrFpj96ClMbT1cl5MxFr6+V+ef8/taAbzd8
vdn2kWcYM1h3/AX8TWu89Tl1zjoo0dvJuUQbwn9OC71Tou8z8Vaxv4wV+fU5ax6O
9M2rNtiAvKDVuGoLAr7bm10WlWvR/FOUaskUDZ2saYDpk52sDcP3gTVtvqiJGi4r
llndfLzLuxpHXtQyt3hQZqJxha6zHvzhWHwm2vRVFuzFcs4WJhdnpqtU1A/Qzm5u
UndqynLUeVBr9f0MeaUlOO7uxGgtLQN59ypwyut0B6bsH7opPBJNlffjx0goFztn
6eoemFU49wN5i3Uz3wj9e12nv6S0363oRwV84ar2saJP7LMA/u3MyZFxL5Vj9JYG
23uXK8vGdgXlfNScbIX6GgH4atEHUHncJkqh/V6VWXI0qa3rlb0vyQjeze7TVD9t
RAiHR/KU//DXJSE0KEBegcMdfRvHZCyYxLjNl6XfC9mGjPN4a3AaGNS+R/izFkEt
vtVbLHoJ+RyR8q/Ofc5rDBUoZcBG6iQka/eTrcJ4XXeNXE+qeV8wlvW3R/pgSP+M
6qCufKvtTLDmtmgZ14DpeOwG0h5BTqIpN+YR8nkZzFqjckHPyBJ6jK466HBzBc7D
Y/xpZ+FmfR837kGGBFqM3C29IyiX+3umGeNqhMuNY7tvloOga0GVNzLzH0rMAnY8
jvYBhnGHYBOOrsudOTdGq0ZoRlbA66upeEyyyNVHf919ozzLSm7ZPzGzjQoj7lyh
tWXyq3XbqAXd1fDdsDW4/XKlz05gD1NdXzxeFcki4n0XbSKP7RBnWuGITl7RG/hO
T5p9Jm36n2fMMBXMIhVS/EqEehloZMkt59X1ZpKNFwjBNb5sYfe8jIWH6yG8Aiee
a6M6IeXOiyIIoDKUqNx3iQjH4w750oRy4U0XXCMzBt1VuBbWjLR0q9SIsZJVb1W1
Vni6W8gm179M3dsO+65ZDzUl4/PBIKHNZAQkumb0QFcUfoEApnZDW2/ou7DNxZod
+lWxscfUCpI2jRHro7QdQnuElc7JgGK7DhtvrXEumoEnq1hzKujBKGMfEUlSRbbj
NLu6+eU3v57G4+c1qAwfayW6r0zr3l8sdKZqsdzolq2mHFMJtXGoo9YvEpqGYbTt
Ia97iUDiGA6JHh/aP4sFpsOklmNg4jqAg2FKodU7/RYQeuhJ9/ITv4LsnnzsJSPn
pxDxA7DZNyl62pKR8QkAkcGhbO2Zf7ioVQ7khNGv3+9Dh6+8NClIjD7T9C2Nu0yY
LA+CIfj4QTb2R7rZ+sR/NzEEcVIk8saKVlQKXRIZn0/y6CrDVJBMdxF6yd+Bepce
AQWO2BYvh17EV55GyhNjIflrTCZeWVf9iTD3mQ1zMPN39DwsAgWHYYBeTkuMF5Zn
Z8831YiVyntFmONMeYspG2310KoZ8AAksRY1r0qPY3vq6WdlYZAgaR6h9jTsR7ku
kM0fdnEZpsNlv7+6s7nYFNuYOn4EJ9wuWSdTGhAs8gFsmBjlO7RbHznATvEzFfuM
vjCMbYAb+vYeIJsXCWZqvysDQUo45mlJWjLXujNP1gZnJ2WkxG6RpyIqQsFE1fDN
wAWG4xI3nC/SZnTVsjMUEbhpQL3m0a68oRpxWDysdMeXB9aAzPUFIEmrgyM/z+bh
ytXODZZPketz4jY4xcFu/wtb+pr26ri5HJZsfKoRp73cIOV1Ypk5oLmOwSnqoNbC
Dli0JBgw0/nFvOZtb2NYbBbr/rt/IjHwbBFBFzAKSxoqiX6427gRVMNpKFfS8yI6
TA7FeyxAbLga0Y8yd616byQGnINY34Qtb+yQYnaQUAgWrUmIH+1twIdQD1Tk+Eh2
ZWXyfWpnsMk7GZuxKv3g64+UwwCQad3xO3xZScezG4BracP2pJnmWrRaXMi1hM+4
iWKEKbNRoLHhV8F35FTBZo79OuufDQqdPH5BhSbB1ES0q+rwJW+UtgYkngeO+WTg
HZVuwow+9BtIn1ZiVMcEbx6y3LlIfMz9A3XkYNCrTgMhZZ0rC6U+Pi7SDsnpeh8B
BI+XxnB2cxQLBoM/akD+8fUgOiOal3IML8DjiF7rhZoNSdnO8SKzI57mVlRJAX/3
Ipi3zVrK8tdfpmsnYsm8POvHCKtFsq8X2YPAh7IAcb9kcx57riWklkICv80arKte
SPJkGxZO0XDgOi3lfb5r4p5L6uLL9izkoTtqHR3lcbeTvKDRuppdv78LCdHjnWG0
VBpteI7HFdfuJ8FcRiT0ulaKFrtwPkFe7QlNzepGUvNxy1WPnkX0rfWyGRDBPd1y
Qr5J4Bxs23+2iP6j2L4YYN3Cbg49/Drvbfi3kz8eZ1SN8H6gY8IzEKSuL8JSy6nZ
ro7RPUCvKqYxGlZyILll3CBoDwWhcZd4KRzqTpODXz/KLuPwCLgPpseN0PRQiTyz
D5bcMdY8GQ3PmYo+kFARIUAWwT2/XHmcnb5HZtuQQHV0C30dlDF8t3zaqviWA9Zo
aNYQMKG4C3/96uiClZEpeH2cjhejvHACoH0kxMmPr9TQJZp+kPfRkw9MUGlY0Fen
u3xgsDeiHOzXybSVRyjDiJMYmCTvuPYokDbzRw+WkjIhf/oYtZ5YFV8dMREgc+2b
zFfevcQi7DV2p3CHwCHpuNC8uEih9qCKoU60W0H4WHHKrKzeJc1BHDbRj2F/OFyT
XPzT8UzuFYwOMdD1R0+JVMi+/Ab+WbRR6QnhqlMVlmMynFu9ybSevybS9IAo/EQO
bWDCu5TplboJkJiUuqbI7K1fw3jluXruvIs/3YaKQwr7duOxTpfyPWz+aDXk8KDm
YoDKvAWBYkMLy3M8laYKdVETljKWwGSlFCwEJ0K0paOVS0Ju4DCRay/fikVyLhSp
HmRhDhr25TQlujPeMAOb9xYmRFwd5LX1qNSBrhgkMqE3isHsj+cyWlC6JaxyuYbO
ydVCXelyoQX3GtgeR9n3oW0md2UKvmccRti71tAfdAcZQy+BxpNPPhGVyY6BZZ3o
ei1IQrnUaqsb8xAGLFMdOC4Cohas0lAf3NUH63EBCaseTPDK684d0+nlsIafwHN9
f13lEtl2Uyxud96UKUyzErLMwEJu4UaxY6ldEuBCITdvXIT7sWmIxS9AXsy7r93u
4eMU9x+ejDNYlS8FQ9tn7HRHEbS0F8oGiDzzbF6dX8UrdZ1fwZakRRZ3PrUaTvy2
0Uin9CYLE/1OOVCu+hCpttgOl1uF4+PfVCPc4S+GJMG6byfKTVc7Ur0T6aU01Fx3
NEGbrdzCww0ou2K4VVRNbf/9dtigZOB90iYukDaUZCQrx1Z9Mv4f9hopmt9KH+ni
qLw+4iLuoCZPALbP+LQtUnF8DJ12FZGd2aDle/e6yAmJ2Z8G+3yGjH/1kG0dkyfM
q9MOiCXM4PVemJENilun/8Rj9aksqpOxx3sQcjzuk+lCsYS9u2VktXLVtG9XFEVg
WR4nbeGE3Xfo5GvRZcA+WGswqy2MS7xBBwDG3up803dpit30I2HaYELCsun4IysA
nY0SMrLfh1giK6k9Ph+9L3kKYQE5Oeljje3hPxqMDv3a/RnzcxD+ubyBD/9RofMb
7zrFbmOjPE+4VStQoomxjDx2uM/hUZ5uIV+hOUTyRt40LqJMaWkpL/YSvOdJ94j0
uoTfCMJ07Wdw7vW5xBJQcWB3ZeTSweWxvQB8wpBaw+QnvKOG2sNOLklAapN4FOuN
hDlnxVVzMBDgZBBYN/oi0sWH4R49StqC7toDvJLs+QU3oDttmURx5GBHMDFnH7nG
kOKcgJ2en5I/hb0jKFc9Y49xo2wI1HvsqN253QglIPpEPcHKV5EoXTPJLsBZG2rL
Yj2hnmv+nib4Rh72jm2lpkJSx/wmzhhId4mKTjxAU9VPvllf7J0ND1Q5fentpuLx
Aw1gIidjXkbHiIxWgGvgOb55T5aPLJgld9W5ji+qxT1SWFFpBOTav45gHe5lxsIw
m0+xJwUanl/X7UcHnphEPV433eu1fM7DuvHxMOdwXOoWbf0rqVseijwhxmM54LIm
AYsqDwDUs3VNpoEDUQn5AH+5VBFZY0TVIP2zus1RqDs42M0S00jF1mrkEy4qzUdG
+USNzhOMbLeoGXUu7Dlpna+2gl2/idwQiBkxYw14Tii1tGD5RjVwGKmW3p6obnZW
Acj4KtEgi1UJL7Av4xmTOMKBmDAKI50mFurDWVfj3zBp06oL0c+evbk0Cs6rlTWb
T2t6sSW2nK+orutWOK7o/RUp/L0u/Wpil0YUEBaPA4kvLgpPo0dbwohT5eyZTXa9
my8mZAPuSPXGbzq7GmxBR5L0nZZCI4M3OmcVmprqoJue+gHQ1VTWCVPiLCoSjRE0
xWlNpdGG56qY7phadWyEo3NeXa0HgLqbXwj6f3YnbAMNkE1XlqSwfZr0ppUuuE9h
hWbhDIheWIEVkarLgh3bu8yaCFwd7C2Nxih9cPKVBh1lIaPXfD/rNm+IWD0110gf
RB44bPu1k7NI5fZ2D9gfFU6ognylRmV+xDnpFRzlg7jkjyX94ZXh7hvq0KDZEp0z
/GeGG3Bp7xmywNpK5jfbiG7qXfIdDzck5TvgfPlX811A2wb1Jza4XsI371tPTF4n
xlQT6BqjDn6g5xlgzD1079on+VUpIXGKT6GzAO0GVLZBTsUb1hbHbk1e3fbycVOu
PGzX52swB+n0KSvGEen/dVlFtnYXEcai132uNViNUyTHmMOVq+FrgPduatGmFj5o
AZMR4siNThoyU9Yu/jhfHhgrLrgo4QuffqUjwqdQ+9F/irofxMgWLx+IWMt6jpmT
Y9iT27v539Rg6uht/nKULt2+xSY4VSfkNAjMY1Nxg6zKCq2cSc6pzMEPDoV3T0I3
NdeZts12Raghgq6Dnq0wpZSqutBRKP8/vNDhPqzTLk6uwqfgcqcIxT2BpZDcjmXg
XTNrWBe8elFbU3mt67Yte5ETe0Umf7Y0cESWdDAi0EpBjO7DQcvOgurqO7zwB8pU
FtgvSB90uNkK91FVyRgR1txoXmRhujLpz2d01id82I3XneMEBMj71f4edOH1uwDS
i0FEHvYMT86m4lwQ/rMRc9Aw2rPn1YXKWURlyLk9BIkwEqYQX3OaMYAR97fuq79P
76sxnoOP7YrLL+toCRPgAvm1N65k+OO3WTTcWT/8ZCr8/0wU+Uryvv2K9wij97IT
7ZV5AtgA9d7RXjCje6tLl85WbWRtMi2w3THwpjpXjqtRXOmbUejtG1qsrnCLHFoU
RKrInDeBYBR2/wRBv1dlo4MI3uewUZT3jz6sAqAZ0DVT2gjZUtyuoBgI9HZhi2fO
WU4XxiFNGDqoiMKyWTKS9Esyz2sRDNiILS5aiq/6vykwbm6+F3+7P1Uk5SfZTtlY
/Qc9zHAOp0vXxTcmIGISyhkjJqsiB9XRj1JC2QO7kREogkFbrcyyFrMOpgxNHU6w
yDObNBfoxwnZbynShRqcvQHyU1tGtfZe9gKNtEp/WXXpE+dqkJjNYlQtfUMAEg50
PdlAyAjJqVEC6MTUrGycgwHJVj+IuDnpptAfY9m5YxT4AKc9mV2dcMW3r8Lwo/72
pfSR9FkWVzll7j/VVaPlmxqz6mkHmfOF8uAQRQfNjGNcpA1Ovov5UsBXgKcPLb2S
u2PDlbukMejfzOibTH10KfeQaueykqDPzsHfegeAWRc+L4g7Oy1eZrdet+XPt5ok
4mp5g87XQFKyEr3NE7+Cj3E4r7RtvUNoHubK/CclqgewPcPkp+2RwKM3fNKD4xSa
9cYJBsZlI6kO3fRxTh/WWbZD0Smv/W6FHB3WgMfDZUchovaDZ5FrMKT64n10oCYv
wATkujJlnePmRVxLPVRkyL6c2JtxwOuXyLaCTj8oCjxXQzYRNn/PtlzEUj50gHX1
GCPrGMNgwlx7x0BIcNmT6ioH/8zDTofO6WjfJolw+Gjk9aZEVoHsZmG2BTaNCncV
dM5DWmaAckqbSzuHEfiEItRVigAKOk7aTM2n4CCD2VFvnZT9OWlubIARTtl/vQQv
gNiujTMDEv/S4fGxX7oUwDE7I/mBKGCmuvISfSyc4a21Nz+ulgN1hE+dh4yoqlyt
UD0ueqQTeqTZPtLHmIaZA35i001w2vCNoFWI6ZvaPpo2fre/13ImqtXSTkfYSvQ7
RtoQJ5TQp9eL6GsjkkOfta2/a9IAXq2EFitw4tHalxwmUIWIaxQXv5tx4z/nMwp1
vRS1Iq505YhGrIkonkIN/tln058QMQgbJqv7is7W+9k7ZtcFrmP69wIFeHPf51sW
ecJw3iaVOOvTwg3VvMfw7YqNDhI5bKSaY3SzLeBDPtd6Z1IMJafN6QCct4O2L4+V
66b0Fh6yJbL4RJbMT6A6tLbJztxHyzJmupYa5UKWwHY/L+g4e17clfuFQVWkf95P
V621zV/zdzmWUUiJLtxc/jBlybIBA0bx47qpLbjKjypuHH9uEKysQ/azcaFCSju2
eqVe5KAXH66WuKDVheOd6PosqJlsSUdmyvtBKY9nW0CbcVvzdQNuqal9D69WQ709
VlYXlb3BVnW9oZjsOj2hhCUi4zXoB5t+StSb/0fd67GP30e2W5XXJDFaZvnrU0MU
aHOmGNUWBKN0ur/DVd0Hq2q/ReQtgRhEC40DQWwTFTfc3uvBHrg+Up495aQsTP9/
VgITcHw6epVZAHq4YnnH9EObRDlGiRU8CmdwAYZ0V3XGw28IaTwx7/9S8tXJ13sG
ctsrBQcHW50mgCc2vckklfyhRK1e2FoHKQMzy21qzKjm2hZWAKB7IKwcJ0um+3w7
ZURDHMF8cLCjtg3O0+qB8xLZAiyA407/tI5hCghkGmTW22frcx/NWxEDSo+4SKCw
n2M3+eIliwbybZz51Qs+KvwaMdKr4TeNJNzH6RIkCD7N1KgCXaQPwvfRkSnjrvis
UPaiYUl9QHrhaQ6vateLyVbebkoatKqhMy/Vcm8fVGqRUWprp/uDcW2Nnlz9GTLM
V65eYxdcGUMFWF1WG9E6aWfXQ0HCs8T+8tQcdDe0BOFifts1fwU3oDHuXm2SyNrg
MLtQQIMGmXdADC0FV7mcdBYylIrkZbLiSpiXN9d9kczY8JQGUDpl3/UZoJhBKUVh
vsyytJW9hp1A6lDMQWWmNNje8H4AX7+H61ILrRdLXKG7ir4AeOifJKj9gTvUnqeD
WRqXzeiZN4wMoSNbhlTFaUgJ0eV23Upzv8Xepghu7hbnmuCHRaZ6Kdg048nq2cPT
RQ4s1m8Z7GN44vL280VSimZegkTViYQqLlA3JnsAHZvLGgMuNXb4MdP8q2YXKeWW
1iLPX2JRGR37ZPXHxT4f23A/ITEzC1kOHINo2SP4As58LUMm+E54MtGS0pH0eLjO
jhIrZhfj5gr2Tw6wekK2D8A0/vjFNAUHPJ1/jAPXfcDuscV3Ml3bh4/dNmj5+KEJ
8Zrw2xaDTN5jySHyQGRVSyQyewfKvMgCNLjidiG3S4zih6/junaeawmCT6YxWWT+
oSHDZWr/fpvlk7Y6M7eQwPd0AIsw6h2UNvsNjBma5ZYOfTLvc2t8IlrnGKPl1RAK
bqtQ0efzpTt82dLDkuUHGylK1cGriTEfkvQAzznP+VCBtVG5SUlS6gzxEYjDyN87
5aTTqswj7BcAE4o8qKY02rus2POxmCps9x1tk+G+rpX7xd6SlZ9WTtT6fZnzOtgD
Tf2FWmAoTsyuCUAhkOFjuGKBqN1tNYqeEJEnOFLF8P1GU1GbESOsNs3PcbcTcHnR
0XO7agcpbztSM5lRGwOOslMN0sDJ00CMvVJpszQaXAddlVxwz9ptWsuh+E6mNPf7
csTScKIk63CevcsQe5a2onXdhNsYfunnSwzlYt9cVS9F9Im6lXJFkoOF8lf1nZzI
GtziaQGvpw4hXO8Uelgk9OQpjogUycz+UBcuI22TLTJfL142s+uI7724i7OTbvGH
wJ8CjC3Cluba3v6J+7rwoUfdBlkMQTY1nCzRIm0PKV+FBJtockJ4wVkK4opakscA
J1XuRCJGJhhOdzKlB+srdZpmINLj/snxz8d//5TczncIfms12rSP4PUlQ9IZLthE
jrI+SnbZTRzypp6MRGFvEBmfle1eBB1BbFsawFvhRG7o+3iUkgJzC0vClcOZlNw0
OMOsO7uu5sX00OIxJpt2vXUmPYXuBa776uwIUmfGTjztRQ1QXivHteUASPTPHRp2
o/E7BxQoUhkXs0DHGswoxkxSC6mPDbys/ttKSZ3kLKsX4+sIeHfKKizBcYpdW22J
keShjT4J8lW1hPtzlyPZ6IJ6MEdG/sje8MEnmuSUgyuUXDWYd7a7Yl3upkqevGJX
dyvn4WOXcuHqGVfqSLZyB6rwG7ueN827RjS/FN91ksCJKnn7pF1noMnKvXW/h9fc
3m3xvlDjusFF57zVHUHHCdUb4lim6xJTWs/jJdwbaY+s1IjjjGzVRaT6ZRVFw49M
vuE5nUr8tXc92uGJ1QQJzbUxKTnZsi379loEZnppyKKLOex59R/uy/kO5gF+Sx2U
VFN4hmjgQBm+QLQG7sGxAwHJ7zTZSVGmFOW+4u/2E1CMR/sIFKY1YJXd+m/DccaK
V9pV8mvJHPq1JsmWm+dR+VdDRd1oM2SoKqn6QuSx5kQiZx9hpM1tzdxrm2CczNQP
ts+1jU1nRyhgiSeILLFLk/SCJigSChIR3th/pMDi6apLNm5WhOYYg8khA7/TxJKl
ux8/8Ugltyxt4+rWXVq+f09yZk/4rrBWiO+H+t1P00R5n+wh9IidokwefF41+i0N
MUXjKHhw5frUkUZk1ixgFcbilv9SCSRpIt3rt0/jI3nND/kL5dxVv4NfYI+Kil9e
jG+BYIoPge55qz1lfh0wxJ/UCpef7/txxTiuyLTQsZHZeHicEE3ZPn3ruTye4Udf
Um0V9aXtMql7vt2TgjMddKo8ELqQZ81XV9c1/7mYKwkPqi6BrfOV53l7eUcMBUVw
fZLmyWmHF5pN/qh4ZKB+StOKXXTbZL0AtqSGnNRNu/vCOtNVT4hIsfz3/7wlojm8
GFkg04xLupvoNwxHvPSwGLT+prERE1B1YQnGTHwif3aDI5z8iGjGmrS76kWovIwY
oiRxQJ3E649v5S3qn/qX+0LjUxXayOe+0fBVtuYA5UeePWXUiGWA3fclz50esZEL
uORvRhQ/9DUQCPh8CsbwcOMYveYHgn7RQw2n9S8zG9vc9JbioXC512jAk2enMtsO
fG99HuOn7E8Aqv0pNeM1yfAZE2Wfj0ffwlrP4ko2HsOhPfB6QVUD1QnD9nzZqlFD
J02YfTVV+A9yAXsi/WP/9AzxQDVIHIHxy+jlXT1dZ+9S7L76H3ZKNGsI+sDHfRhJ
+m6zFM3VieVNbNRHFXr9dEaYp4aMlPXnOCBUL4UjGf+OfGDmXqSEm9QwsU1PhcSP
6hWFBCxmZYEBZzLQ/zJW4GdQvCvrGY35T9nC6n0CxL1vV8MSe6XZunQZn9Qq+1JL
BQJ2f99vatnLQX6brK7vArVfFGSDwMqYSKkhvfEm3G62qOycDSADDdExn/GFf6fh
nDfXKxF00GV1qggiPEEzDpyVn6lcdiM0ZF/49gsyJqxeBehs+9Kk4xLkKXrYM7e6
5V+MFj4OFdNTIzUfE+I21pKRm0y42mh0DoiU2aQUko400JCWihg1ohnXetAX6+cL
tAX6CheqwAtBpDyL2prB14HY2C0qvN9OZq8E+Oihxl1OqfFG+vuBS9b9k81WlKlg
OO2GEY7IpwyG6MrCZ4pVwSwLi8DtZTDd0zaSb8eVa0yuwo8jbqKpVoSkrfDoDx3H
OU5PrncqtA2L/cjhrIyN+gI7dI/kgDJwXWku17xqt0XbAwckzJ1lyRkTTcpfzBf5
U/qAf7A5TaLY7C+Q0kcnb5wMkBw3+g6iBN7IdPgaEK68L8j2JeDDI+8T9kfOdsVJ
//PapYfnobvl5s8bBGWzO19vMXbZiiOQSLLF4LCD6ukE9qj8bwmrWYfGa1hbZYIc
YlprVxELxomvcRmcCoFEHjen54z4dKq41gVRGLjYhpqUpgd70bimwFoUA6Qr4UhF
XK7N+mB2+iejT/rtfsr0ens2YiqhC3TnHK4kw3JIHzY2kXDHcNqArwZ3iFVntg0e
tVoTp/7ph/rbrivjrBgL5jnYqSpi35Tn3fhVGzDv49xfisB2xX34DPpjNiemDHWv
2ywmAoFrfXQ6shdXzOyNmItMstjXYhkpxBgk2K0O1FBDyRqXfdsVktX1XcSo9CKY
6Pk1iUXVxvLQ8JcTPcDy+nb+u/ESf1kKdqa/D7VJGYaBH+lZYbhqY8PMQYdMJrPR
G5oZ4DpxXy2kH2+TlsnK0uobwhCcBDkg9C3GB2L2KldfnqTwWxMXtGak/jJDkYpg
/LXX26tYqIAb5uFpnD6exX8nQMZfEY7Rwr7vMAJwq+MyRtHBS01xUlvrgOR/2CnG
rU8V4TlUJt6HnaiG9ubcy/Svp/WxjZ+17YM0T7asuhwAqGQdWsh0rm946cQBWqkx
uJCO/rKsVXIC59hK73Zx7/n/BVd4PPsBXe08IGDv0EQlfnaHLfGmRUvj3EaXb7PW
WIYSjmFDn12IpKrhqGePy82vYPVIemd8vAz6BPWJ6rewMxOYXhNSHnQXMhl8Y0HA
5z8DAiFtzPbZRnSTsVWshNqAO32uDfg5s9mhrYImsrrhpxdeLJjsTSkB1DtdwAw2
qDINRO1tA51CN8lADpzBKHw616rlANqLB5P6bHPNJ9KMtPasai9v0qv9zPxGFnl8
5qjGxoSe8xIAU1i9OEbM91cgOFC3uMwGpGaeQYjbfxkt+xeY0JSeW3lWwFdI0kh5
pmJYexB9SjnDDoMgoVOtD/WH1e12Ssq9oT6EaTLadG+cu1H4iUp0QKF3ezkKR+KO
A/PIPg/8zVWSBBnqaMVVIAVlZJ3TsbMZa+q2WAlD8Ohg5e8MHdB7PRw1Y6T3wX0X
jXO9wMgXNbIxX4QZHXrMQIYtPaxIXHDGbLB1hp1sZsETXQAcprG4syPsNGQNGCJo
4gWbQbeSf5k203379z7S67HVvHG1uTeZmz6mVvQsaQvKlNySu/5vx+42dqVTG7pe
ZV47I6GihZAL95c8b0PnGjguSNyanRPkThO2bgPLNp4G12/LIwkIGNmNue5nqa/J
qdPovOmnH6956NPTvegfqo5CEA0Nzr+5lWotG2vdLg4vWMoDDskcWbOLbgvv6tEP
NbG+4rNyAxo6VxROPrIJIYknjpGNc6Fqoksjo/CFfdL1t5YYTzsYGrEPW/jgX0ee
K2B/2vep1epTZGdBKgEdKv3Exf6/O6LihuCsiPY/DgjQj9vDT58zFU7W02KYjeA6
nsBkdpBh93ej7xSLZsM/05IQ4rvVQ5zKK9+h4AxeunjX+kVWjexSiNPWTImpf51n
dxWSGIQWQPyIiZ0Uxx4wcva9kfniktOCxWLtqyrWk5M153sMHCqhE7W3+LgEuIqR
w+ZKGQYT7saYh/ei8ozIQsHmmmXbq293GcOsWpS1JOgPkVXUCoBL4U+hLF+KSGyd
rOinHXEW4WPyJwbwnjuxFmDLp+RN62aXeW+HvTUbCSXsyimB8M29y4C5PnwqGGYO
Mqzjnu9mOMQ6LlFkz3ddsF0aURKH6k3Bod+YnUOduXwNAwCIwrzgcH8rc2hPYnDE
yCmrEmR7EuGqUmwwFN0KgrFssJ4FDOzVdhkNX4MBldy3piDnrQoroBNAQzOqWNPH
zkfb8xLrsM7Z+GaFFWcuP/+cXwtpqiJRm0ckJGJGHoYdJVpCBgK7t1fmvXog9AWz
yMo+cn1Z0ks4XZE4HuNvKPs25YNQOcfJssNXx6hzcC/KHBOGk8UwI9X/0B0CkaMN
KJm7ETpjuldAl08D2JYAdkHVklj/i6zVV8Iytr5d+eLYSzl6bTirWIw8AcwTLjSb
kcThAwfzJgwd/72/vsuTtZQEVXibPoLPMlLIRdYhjV4r1YsrENmO+p+sJqv+5odZ
NQZ/eX8wjQcxNBoHBKCot4HjmducpK9PsmRArXUZWwH6PIH/aBIaPg2ia/K83Ue7
GZHfri5jUjfCQHb192kdeUfj5893j44rOZkRx5c0NEcVLDgvS8rqrn8LorUqj2FE
/HS8Cejnuj2FOeOB1id2A+zIFrjN79Dv16r5aKHH20KMOwVlOKLqzpBfF8oge4m5
8PZ7S0BaBBAsj/FC/Fh7w7EVKNXoL12A85MLh1hzP9+/qSjv9yuFJhj+JeLygn/V
2mPvDgrQdtJd7+kAwYUGv19+yMiXg359vtyXxzdSx9jjXmLLgEqhNrXd+HG6o/jf
z1NvFGZLfqtLZoIvZpuSDTulv8xcVXriK5q9f0olPTuv9J7rc0ztHNBpXXtIy1Pg
Us2n6G/PpHNcVKDvrSsF7x7fkQsVtteFOJpcvEuS8B6JwwWoDuUWP117qIGR5BXO
gr1G7VsA2tTtM6WMPvtBx2qVltU2hgO/BXsWWS3pnqv1/yACralqoiAkTeEfCTyw
y9lgH+xjQHe87I0cefaSGGii9GqxU83aFLg9L/6HrvXk+/QukCIR8OuGJ3Cx188A
C8AdOPMsyUP1KDb/rf8reDCQkUmhCbVp7XsMTYtLa6zb6wQPkL7QBLuuTgV/tUg3
6hCI5T+YZxHkIT7d99cHPWSfRztiZu1xR7dccmrCSnad4sS8fbM3LuhrQ/jjWLiC
3HdO7tDa3lxyYX7jcR4iCbQbYrBDWMzHFNDnSlKgUE6F7e3GCcLPgMIDFeJ6Kdhe
ZCyouk7/LRYRTqzDNBuk6QhNC+yAzZ0zr2TjtqvPNRr7g8PqaJQM3YG60L1VOmyv
vXKEenKgjGP7qo8qPbXINUNwrqmLAtmyOhJPNLcbfBG5eIedLBeWkF/yB05WPR3u
NBaFpm7HpGIstt7ZxHImUruHhkb9212Z58V++FW3z9lyCoMg86zJnqnfufkxD1Tj
TbmwI8WKQ0F4sbmVSMLjudGPX7g6FzyyW508u4azwB1FLrtVTpD7jSBhH3sezpm/
yGto2gkHqhelRmW18ocRpjgTlDI+ETbfJWDNyzhCg+Iy2VtctNhzcKKhLIsVsPl4
eZi1iVpbMIB5h7BlPjQnCOZTdmafjgU1EwsOJ0AglRn3oiBDt3J9xU42ng4JL9++
m6jMsGrECA1muiKwaaXJHBKo03968mPfMU2baOQ49hdnmOMBNj+QaOjNE7k5QVG9
NpduCglFLc2UuXBc+9H60tXfQV/ciQPa7KA1yhx0fjtr+VHLPPoFuoJrnn16UMP8
hmFwB1TIz6uQfVIeZ5xD+jIBa2ue8TgarVnNe1Zv0XPZY4TcNxgC1Kpnl6Lux2Tc
l1BwhJPrrt1XApTQvl764dRq3z2dNWQZGKlFlIFaof7EqS3YgmieHO04r4mmq8kZ
tTybBScADLGr3JcBr0Q8IPIMRw/kIjR6fKfqGIAW3DCEbqCzYxWOTO3Di5mMA9yI
0qdLFJYXfXZ+YFgoZy/pIUSRQSr46Rx7Ryen6gGVL83QcWPMyVIEmU9JDCF0Yryr
ZlS726FGk8gtc1palHiNp0xZ0RcGcwi4Y5pgnJAH+agA8DjzjA2ftAnuZzpoAJLY
qZ+5X5MA5old9ca/vMuctb/BG9gDUUClcSgSx0FON73W/qDuawZ02bgbWoVA6aZY
WQ8PW5gNxVRqBh1ChtNo0A507qbH3HYdNEAsixBnX23jRM2TvkoI6QQVhCh7J215
3IiTUtspNZtUTZpF0YKGByTNeaOPXU2TlKjtX8eyKUTg8Iv6k23241hzKb0tuaaa
DThEIaGogQRww1CPypdTWkqbUbEUSdzK6isV6ztLbCKRXNyhiVPCdKSXAP6BcYz5
CMCH9ZXBJwdidmgsVNlrTPci/1NOnV4/BqC5dVQJzl/OTbMuMj1wy1b9CVLNJM6D
RIMrfN7YVH8XWCBX/XdyDNIDotYxM0BpPEOg2ybo3fpCW9CW7J28W55dKMTAvwG/
bGLVanmIPOinaRumgWxzACg1zQUg/TtbjQ5I6cVjsjpAt8g5Us+zh9pG632ZR8MD
0wMPZ0yX5WBH6pC5cDmVfUjHwDURuQLemk/8M9QhA18T1pItVquiKUx+crjouUuM
DOjT0hg/QE7GNxx2g5qwZ4+pSGYL8cu1CKObYssIlJMEF94CmJB4bcdgl/tXZmM4
pTWNh8EE/WPmqR5UKHW0dUxmMex9n+LZcTbzPyPGNjNy3foQISFnHP7cYxMgACm+
KK7HpCguJd/TfoZf3tzmK+C52lXiouZIFnCF2yoQRuMoowASaxWa76xrIs/4We/J
tAz+V+simKId87MXdXvLSd2wpyyNCUZytMBC5tJmg+OIjaJUtzzzjEue5RHHvmq8
Rk4Si5ADRzx0OIPVqezOZGPWvpjTEj9By3+3ga9ZOYa26sc5DzCNpmY6gj1piLUG
1faz2AUbUmF06F4YFF7uDxmQancCz79j3k0nibvzIDH6jx8kxyp3fsvlGJC/5XbT
WHDFT4INBWJUMM08N1SwYbAhkdlrtG+2OruqAMXSdZ5ek26EQtT2CPnMKM8XGzrZ
jFpljii5YWEb4K6S6ESNp+atnbqu9bu+kGPnVJPOzRTPi5PnbVgPqSONcdCv0sJ8
nWCxmO70lA6mjN9veFpjaUH2ei1dUJWKZAcHcvxrfyepv5Pacv9v2yTOPOUdE0hW
Vwdggt6G36OhdBNF1PYYbv+Q1lEjofV30tTcSm/RlS9GQtnokYHN8nOax2SlzsGk
7MJwqJ1ps63T5KHTFUKXIUYkDTkdWZw08h8+RxXsitD4M99UXQjPPVTtmj9Rg5/s
ZVAsXOaZe2QI3X0mno9yxPhkbc0YZty951nXOZ1BtS+8ifxmnpwz9i8SHxOMQnYd
JDJmDNBNPaUHkYIa+axR8icT0Hg/tBWhQm9iFNe+A+WJ5Kk41r+c3OxZXT8MNnwX
3h4suoyGukSoMGS6VcpiwBoQv4ZePBIAsULPWTzgSD7KnykMoqpZi6M7rUiqBXyj
yO1UCji2MNplLbuQq+iXWCGzpSFFJNdvfzlPkn2+tvrpFfsgFmTZFZl2xOINJj8k
obdd4+1RiaydslP9v333UsKlK9DIhFBykPXeLZOBBmIUdwe7ErzONJ+HK+9+Of8A
Z7OuzeS4pqMqLTMnZZtDXi1UZ8XUi3sGLW5RvOlRPpfbBFSkz3ZSfnG8+oJ+XxBp
zf+w4NPh6Z5pIfzYRqQyk8pk17m/9kMFSkCcsW2VQCJ+1y2a0l0HPU0c+7JHxHQ0
V+xViBdJSkxHUSp3SW7zZst5ln/jfVOmnp1v/mz7MkkR/rTRhrEavaRBWxh/+Rrr
Avhar3H89p4UdqcG8TNrLTdi3qeF49wHN8v4U72k75KWx/xeXc0O8BzPmqc/GCyC
FzOScoCwtFfBmSY4yTwRxei/sxxqZKuyQKUl8WFt6lKfb48KP27GwGJRWI4+1olE
5IJgq9t7h5qRwZknNXVtbP0J/grFgsB2m5RJMpWB3EzKp9hBKrm7qAN2PB8x5Se3
jItR27H65tVvPjJ1LZFkOyUFRJ2o/BkE9OfP6LyNgXmmn2Apx1ciZWeYVP9iHcBs
y0eaUjxAJEnbRRHkIEnJBHfv80pYacsgcutR+bPtr2OjMEpp1cJyxuEOdaU+caDu
skxT5f4GF4F2aQFFiapL82A4vKDRIuzKUdwEFPcA0Dnlsi+PigFca8IvCkTvKc9N
h3Yv0y21bOCv4Vo2CmoMUqVhk7HJNK/jtOiuPwMJeQEhFIJCSVaOo2wo3ZRPoovX
CDuV3jU6CpOMCQT9CQqs0CRkMxs0fgSPlhoH20F7pSU4FsBGbWDDQPAHdZmG3p9Q
VA0aWhthA3miYKRafdkZ+zNEImpE/L4YNZX2agQqmrbSVtMYBF95vKSrShsMX3aT
JRukNhkRkIPvuv5syTfzPVyIutpR7yc1GQv+HPCb6M0oUFbmZI0Fqq6ZkBsoDVCe
gneWeIUa5IyO1n5pTdwyrMDXaWF1g0wC1NYwY94w+Ye/OEtxUbQk13VzzZxXTCfO
6Xp/Vds148v6qV+hCHC2ygT78xMAHJyjJ3+6BpKGzb0Hnvj5g7GTKD4JFQQ2bEiR
nbGxpzp+S9Ygdbq5WrpmrRr8lK1FWHYWQccYOHXnQzehL8SBFKFH5zziXbpEKJZF
RjwvYbSpSfFfBwL0DZZMRidl7KD4Vdl4FA+7IQuTCCoqwAPCLu7HEdGSucnpn2ON
3sdo8TUDOnn+pEAzrJ7+uaKMBklKk4T4uXQZeXcPnh/0BBgL9xtjGPiwzbHVFW/b
qn61HknjHcWBs6BjyX2C4h3MX3y7ufYUInyfCOHWwlWTY+AntI4ZT+n0r+4lwiIO
VY781oN5Buayp6H1cXdexIrgXXncmylD4gd7GzBiHZusgCtzG1Sp+0P87xvY5+BE
rXjq8NkQQhdD5jvqP7TMuQtQzIqLrE81DHtdeek3Sw/1FrFA3mGu6Tq4n086LR+8
HgdubMgYnBZhLZVyaTVhc3rCl3V7aHbKxNG1+2YT2xhYjmdpRXcJ1wTsE+95db20
ojSb66/tAT6P7Jwr/MjS6Si62h9khDaoY3YmO1BLAFDtHfaqgwKaF2IhArSkV8L8
69hm0M974TbMHpl4fxUmtyD+L8GahlEwNyc3Skxlctloga6cHLZnl5lld2Z+XYk6
+F1Mo9ueVNCAjNh+OJT8VKYe7FLDl1zwxMs1IjJsGqcUv8lwGUkBUfh0ehe4WeuM
dqe4jdMbaLNZ8FlX9VyqguYoHy79QI7uSzioXEPL7PI6HjUwlavw8UWDg52Q8hSs
AidKdjios52OMUFRdSkgVohtFYjCs8Cq8bl0Ae0HYJo1D1o1xMDXZt7KTsE/C9X5
2pdxF3IYCfPigLRgQz76GlxDbrobve+jaLDodXvP9A2QnS9SbJpfwaVdK80UZ/EC
yQ08Ty7X94MrgMCTdES/vPtmGVt0yLPECcw+AHNkdpM0WtZfYPeO+ADO68yHQmkP
RZuxRbGmBYOt06dh/+q8Re6vyl3EGUHD1ciUS3mJkSrRmV1TrCQBiBAj3XdkuCm3
/qKbe9ONm6yrnMsHpF2J4Z7DEHb9FXDe43CEfjBBvQnsLYnaG7QBnDifOyokdCPY
GthIcM9ZuEEDKKKBx1R50zNT+eIBy1E8i5bMMVbn3/23QxdQYniwORqFl6GzHTF5
mdiOOGYOqzEHirlEWFxEMTHyqWd1bsflsdqCzWrvZ3AZU0uy3W6E6Cj2d+aHHcrZ
1k2oMwx7btiD63Dmj/cZJW8m+n/en+uWrYYl2KNZutnuTYXyDhCehnoynn+NJc/8
HwRwRSxQaZ64pbeZdHPwqyF1c0wfI0ouSlYeu7MCqY+3fP6IHbpu0T8fSp/+FgNh
csgVuwFBTltDO78z2JLlIYAd/F3B6KwyybzZgcD3DaT/CzTTEV7RlbW9p1/RgsIJ
m+YAPDQCHySpQv9TFQFlX7oREZSzgIVzEjLe8Y0jLXvo2UXAb5P1Er8/onSp/539
6HJwqWAxYOfB08nZBathX8VSj5RKKXfzJYsOYnF83emiqAtVfDxl4+vR/xnWM8l2
oZhD59mIIP/a5CetitErIbSlrRZrxkYS30AIvA4WC76DW+szrpphh47rC2N7MkmY
Q2x/OlPVT1P5cG7i3tqW1+52vmbrG/ZhutpW4WQ437yqmGY2Luqna/bUcnwkaX8q
WlPMzMB4Bp2ecWrfi8ePd+egzy1b6+kmp/c+wWncC/yqESrV8ujS3hGmXWt/BXpo
xk2j6QGemrDfJe/C8d7AWyOpX+8V1jfz/iCNH0f9SYOI0n49kUDB3i9DVfUuYC0d
iY9HBQpZutGww9hnIMt6OkjijsmW1L+nFJRgNeLiakpByf5vBOSgP6vA3NO/HN4t
NE5QJEvmGu1J8SPfHSg9UjWprEt/q/5qaOMApFqCzNbW8AacfMm7DnovvQwfOS/G
mmmTN7S80o0Y6BRkeH9PS7ttHAHSEJisRAQabcCS2Q7lBJUaz7AUzIldiAHvsj3A
WcLh6fJ2FebQ5PWMCmMMFsU1XEs8YOzE6gotormLeKRVwYI1YVnf3QqAgobWaImZ
l8RTSxHfDP7yjKv376mdHeKJQW6RsPAQEFBd5nubB6LnKJy2IYVFoEtXyRDwCFrc
d4pMi+yUNfhsd3imeY5v7O2JpJ3rXrH+6jSVpj3RLsX3SWVlJYyBQBpFCvoHENeT
phttDc/1xjtt0JUNo3zyzIlBqBNUwQF+l3NOM6/OTFol4/jbKjjzh1nHVjfMosNY
owzBSM2o6yO62NpFBtHZvSpKlwWNK/fUb0WnY+fuTMXsSAFC93TjKO966YvbJ9h/
7fZXvyUcy0BTutFGZfMZb/ojagSaLhOXToHAhEXz+hdl2t7EYb4jsh8rWcKiq10y
uSUhRjSi61cV3y/PptInEh3g91n63aDbUIc4lJVkrXZty8r03RahRvrCs8JOzWsK
cdDUVMfqRwaLu2iPLuUMDQ2TMcf1gTTS0EBkOHXYcAsxD2M6RcrS8Xq80n5+nMRl
TpUYNiuWg9XDQr5W1l3OaiSo5e62sPrVUENmedLxid8wIVY0eQMFtkjVfj7lcFO5
P7C+TJkf4UiUo2LeD2drVM3okvo7/UzbLNjP6VscfONOfkUwPpwWGbrsW4VrtHz8
tEKQOwo8GEqtgMfFCuEXUyV25oo8kOzQ7EhGrXUERelN1ipW5kSL2t9eg20YSQJ+
KUfIF8CxKNzwZ5nVZBSWbRLrpENU1fjsXfDj9A++8BTZTJ1Hu6C77wSIlFhWp6hy
vu3V2LxA1i4CRZWLfg683UpGAYNPTZ5T3uKq3AC2mbKQoX/ZeP+1F3PGiRVN15Nr
tXof/mVW5UvpqsexwTeZboFQ506L+zrSPHI7pt3h1qi3pRYKq/UtWlLwXN0Q1mmb
+U18KC3ljA07k4XpM4zKvpK5J5Wl9/STfwsE4lbN/FmpDIL0i1642XFu8fepBA2p
X/kzjni03R6fjFWNFzr+RFtxoYwZrJtkKRMdGSGxD0CQjYB6tIcAaCwHMCWLWZes
O7B/A0t0udNc06RXuWgPkCDuuV9lHAxcBXAk/ojaJQQUTLufkmWQEde2/dVYKGHr
VUf0jfhbvT8eGrhalvjV0yetmHpEALe8hlJslsRvSQAE/PS0BjlOzgrkzNKgmBPb
HcWZ3O1m/MJpBMSFEOirwpQJS+NED0yHJmXtePXoYJR2PCy4FRYREg0FRe5KpzxF
fRzZugIjqnobkthlfikKZZr4caMTX0NKAsgGXKYUkdgkA0m+4u5HLUYvNxLYj8Nh
yYLwz+hMRlr5spBUJpuX/a/Na3Ww862OIjdKYcYpamPadeWoHZuYiQMgu9qMiNfm
Sve9g/OkbaNEn67Wtun0walARDR+1Okj7lRgmN62oxCZwKpmC1mUP1iLH0F1dhBs
dvUAnnZSs+4qwligT+4mB90pboj7CkLQ4C0WYrYltWT6CW2oYzc4RxHhD4QKBvgD
xCLNbEYSn/G+4GhiHy9SA9bG5ViN/gBqvErG9tFaXPjHGx3mImGiFFd3OBs8A4XU
53TCB9XKX6+aUuq4wy35qOWEhkLsdYtIbF4bCG7L7OtyqaARXHBwOQEx2AnxciBo
1KwCnCTQYqc01zyqGdD0seKipOtrM1yHavkaS1223XV9C1rQw3e1iOkV+pSMLi+0
RUFbWO4gezH9mvxowTwmDDiJwnldSoq7/JTFVeVfnJQ4yC+uK7VrZnPatyjjYsZ1
yTiNgBfvK14Fl0HC5AYoDrcVMEBUfUIbSeCScaYPwYFrkQF9fDMrF2+HK3FHQjNc
7qVL8dK1TMzvpBB/+VGZaCcg+4OTC2v4GhuNVUhbHH8qbgJmDOJUg0rZx9VTX+cR
YOK53JA9TfBi6h3gIXP24m7O2zBGTl4/LP/knHWd9kcp/6wRKjw8kAeZcpY83Akr
QyKRgoLUaLUIwRJF7EMJnsO4FrWUzPAYLdwP4rGHaQLZiv2RhwLJEyO3yGTO3DVR
gf08soFQqV1WEEEVkdEXe55q+Q3EimOGL3erfwcLtvwImVj1gYmUViZH1EQOf1cQ
S4XWajzvfp/BqKTBw7Vlep+3/nEfrYrlb90EZbGWwC78CBQyVxuCOSLAPFIpYr8v
MiBPrwJWukjcoNm+H9cEnTW/2KwqKS+1f3OgEnH40ZChqojFZ5TO++pEYkJgPWbh
fSim7HYNfkpV6Ps31zdE+J9etcu4pB2zsBLDTRgSow/RQ/7vxia4Gaw/5ujk8q9d
DXCXa4KvgG4rNLwsa+2OpWQ3d6ian0bZObKdQW0O5WQmaa3xl1f45ZWouxI9QOWx
W3xWo4RRLwETVeKbOuim/zr5URswda1SMxpBRi9JJxFLktpX4MaGOp5ltY/cgT+T
Jxu7F/2QF0r7Bl6NkbAfFiiUcy2rVU6DFpDj/7Z+gkzxzbQUN3AhSMqIyEIoiSQK
Kn5OZ5YEAC5bILAyfqL1qsuBxIDuIdrvuxCRW+OB+0rvhGFzWMlsl/pxz3dgE89+
LsnBaTIquWWUR1nbCp4uofDjzXvaRpZkT0499sFx825z2cza58DwaVNmeLJXRIoh
JV2A5okqYT8Whc/HPO3GhCooK701PqfWMUn30oxIISnA8jj7Jdmy+EkB4hJw6Ffx
ASKRZULkflbz6PTjTnMh6pwCO+kcI0ZDEcgJhTn+RwHcl3qVeNJtn2K64XnIDFxe
rFrk8p1gRKA3aW89l4K6COXLkocpvCJ17jRCrWurvl9V4kh71tjku/Qkp6XOzDGR
hf/u5GwG0Opmlt2MGm9u3KPnxbRMZHi1k60yHoVgz4r9KY0OyDhUy40osi3srddS
UNyTTxzHn/F1Ae3pAY5JriUvY2v2DVavwuV4tF3LGgKZXZAycVFfXkwr0+bvOziQ
88YIMJEmSns9sQBH4xwr1ZhXOcSp3bUpcBinJVMCpC1pIWvmjePPckbx5pLWXq9M
5UH5QdL4KcMrADAbjtM8s9Bce/EwnujfT7Mnm3Qcw+0I53lPfkkUFvkgBR2wOIps
3tkuLPqwHU/DFQDU/0VpOk1QPHLm7ramaXnaAS0BunZhaXP4BzGdjwGlaSxr/F7/
hgPCUYCwOeDbGlU4ecausjfzYQ72/7gjukIB2Dce5i8VgTvBdjexLnM/l24KSsLq
fz1+FdHDC6bGI1OTJp+z+pYt8SFBViqjbak5g0K2MxNRetfPGWlzw0p/peqH6ixg
zfLLqn+QuxfhndD122PEv+5sSYsX2M1u4Hcxhz65b+zjk2dZS7Zn85Uw6ugdZpBs
Qpfvsk2fydpjVK14n0nTr/U9pgkoWTZOXB/yCrKAo1sOlQSV3amGJtuSFjefeCpH
ldZcZX1VQ8fST+LUWE1QvUKANqMiYAoe2zkddbMaPaBRGUUBM6DmUUVG3n4MihbA
lJe5JVy5LFtPY1qFl7RCH2rOW+esZAHvxqRxr+gFiHhm2xuXNyDlD70m6J+/DAyh
RNRJkZQyrJur4m/Fh0/BpXNMY8NdtTEgVMEAcUCnSKgRQqewhV2q6kCtIwl77cfs
WCBIFW2mbZVHePVnC849/C7qpXa37FCCc7YxmwFZ9rneBUbKKrlMzPxO2bLT2k3D
qxuDjcnYVPukXk1s/wC7/21pXn/toO3jWxuO7hTRx+kygxbAMCH1zUrQhXvEcG/i
VsB5j68ONrZsyCcYGGBNBF8mEnCEJFow7FonQcNxk5jlKryznUbNL0T7VlL+Sg1d
CweCqP0Gpml+nDWJ2SALZzKD8VLZ2Oc3wfkM6cv78RWTQC+J7UkjyI5ylzcbonP/
756pq+UHCio3v7PB9TZne3R1Mo3Qdv6Yb9elAkgYkAIBGgUbS+8vcfX5MAze+mwZ
puth+nXupr0UG19z3n7N9v232h7MZFs9RRsdtBUuVlOuEaAv+/Aj3X19j5qcR2eF
NU7kva1MBoYYKLmWs2g5OaWW4RBTLVsl5axatpdeArmF4je+vZ2qW4+dswrjkh/N
Mq37sr+nM1+3Ukzo4PffssMsL+hL8dEQ53kWwPe7c28a80aA07i4H7wakt2JWuKj
ncM6/t2VH0iii1AzV+PLahL+OSI+CHcy9au+NEH9YzO3r/T3qdXndB1JDasZAjZN
Arqw8PyrchtE72kcwqKKVUO6zs2YaZD9fPt78tm8pAwNvt9xvtVmM7/wy1TKm/6U
dcNEXeffXa4vq2nZNTlE4E+9R/2zpLbxTmxynLvDaVukE/8opYTKasjqba1UHeAu
rm/4uO2kImlfFI75Q7JFuFth8iOgE9eEgDsBMGvP4iLnxFaV9PXESQ1UODW4UHnG
iYM7rKFL8wGWKvrFEHtpyWFeNKdaX/oTXZP7kKkm9GX4JM2dcC/4w38NtyQL3pUL
V8JC33pvdT3At963nTVfzw61rndZGRSXVQw0GOKonVkC0D019zC3wHUsnwqYgEHb
cGnBeWXCxpAwqCA6MokbEpHZd9W/cOto/SjeDkXoGThqliqXmgNVT1DSqfldmiSY
Z+H09XiflMrJ8u93+GS21Y8ALX2Byr7FWOVtMMxuB4NfHNcTcax3gxHVOH3vp5MY
ojrK08TwY37AeMWL+6AE0lJiRdS62GLdJOkAXEqTIETt1dGqJhX5E4HZjiD7SscT
2I7l5iUS78my0BHT7//hbyi86h/9vYAPfuT4IYDb+4ZmglkzqX6pxzeQHcrBBiF3
fbNVXUoaovRJaHILnHQ9cS8zxykCFCCEgrrzEPerAv9gNVSwAWEb0r2IsZRvX9lo
dpdYLSDO/tIZWwPGQWuLZ/pQ1/RVzs2jLR7iWPDkc078uG+iwA3u8rL4gR2g2mIc
70o00DKHEIbfjG4ySFVXaLQREn/DuDIKwH6WiFtAnsCrSMFKuYmEUN30OA4KjbKC
EaD92hKb6dlo4CZZ6iEClQ14+nULoS9seRzNbTHfAhlSxn2U4aWuEoabXdnGnX0R
anZmMOvawXQajGOYsEovSvIjkVxD23qm/AmnoSqtxRbCueowxVTMDjgyu6gO7RQ6
rdNYCY5lXiOlraHScm57AlQUqqihrpePpbKmxrj+g5lxltvaw/IYwHOyG2VhvLWR
d179XTBBndwfIf0r4OC/v99Zgebh4wv+24fcF4r/rO4JDjDdk2gN2SCy0o9enneW
4LQyCQh77eIGoygCePHhj645V8I+8Ey6+mvrUw/PBQycgDyepjolDPCtKuUDmRVB
BExt44+1Qm9BaTVQmZuDFU+CFO5zc8T+2uJWVdYdkTGGmiAe8QU3ul7WhpXz4Kow
3AXh2lce8wNOjNmylIQCJk4PzWhMwJnugSEk7ioOTvFYtcYnX6orumx17MaJiBcI
JRMqAhHkg28GI82rfNmdsdwZCekODo9QEAgYfG2aZfQR61Z34B8W0kTO2KJJsiTd
ASqSL84lwREZAK5954KCc/513E/xYhpjX7/NLvNUFOu78VgCJcwbhWDlR2A0nY6i
K1MwMUMe/sOMXw6fTRMjGMEdkRnviGf9zigO7nXva78bW9+fcvCtvsLsgN3u7JFR
qU5K92RU+J7dSIL4kgJ7A5I1a7YaDTZPgVpG35I+LA28C1mSV5VIID2jhJt/VG7b
Qb8jZh1hTgva9DWAD9m5GndJeeyLUaBVHCWhCpyfqctgDgU+aEwoiD7+YifSN5IA
YTJr6yjUPHVgdYdkgxAwGtrwpYwo3aYX5mtA952EeM5GTPWHmsnAdNEYQwj5nhhc
rteZ/NtnWweUbeOkwoMtT66qRIWoEm8RoWLCwrEIVvSp23WPVXNP7K5BuVRJaeN2
2MOMVOVdZ1BFVrluvW3SLGtxYfbfupO4H8m4t2Bk4kpbhBn3QX9EnmOwZEDzRVo6
JOsu5fUdD/lKmi6pEjrMiQ==
`pragma protect end_protected
