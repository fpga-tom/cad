// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:30 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ww8g4lLiuMyTPev5n1YhHKwsuSz1Jk49jyxbGvEYSoD/2MHX4LHTer+m6OfXy18p
hIkd5Pd1ybCXy0B0ez93QRAPm+zB/Pe4wXREyI0lA3V69mC4aDaDsYiNkLf0WlLl
AiII7WW+CRU8oWy2UwyIa7PmrHXu/RV0Nea9MFTBy2o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3328)
pppbfc5LDici6Mi5kvUhnnSwi1A7W7/ufmjKb/wW/BLkVZpkLrDHF6ydPNS5bTF8
h1H6V+/h8qPJ2uhK6rcagVK7a7fR/bhF6gLuqgGni39TekRvH2s1/2oPl/i/vEYz
sXsBZmh5idKTZAr5NZERnkmczdKdv/YdORcyfypK8X0MLdteVZus0gTyIVgFQ/n3
Rvt+jeLalNa6mADs2CGdRTOlDH372800/UUmztRhg/RFpQe7F76Dos7xSEjoQLQc
S6bwWt3zoMxxL2OlpJkzY+jVqvGfJta45WYWtX7cN1vRItLzsElVy6fAo/k8X+1A
p6aiEAiSLn7HAfTndNWOdWjaiUpsckb8c8cxDfPuQACLJxsDUUmlt+eqsO9pg7+b
8piem0xpMk6/IFcSyzIvgUvyhpIC+Y5B+OHJu70xBxpZGFwWSGJFme1uAJnlqrN9
F1Ed/U6OCh9SxTn+HVEFxh33XRmiPi12N6x3odd2dYQIyszfqhnIxpIYxjbdhOsT
taQKrYrWKzWA+4TdmQFSYpECnzovZlPsDZd1cJRUpI1TIqPAKLJkDJ+dgtyG98PW
4J2PdbjnIlB5ucc8Nv6N+TPkCprfxXAAcc1CiGUQyWgekvdzeVeLmcCcVNtUFOsE
HML9dwsMZKvOrm3a4gbedQ/sdru06Zurlt5LrwcXqGUWk6DcCdWnB1762ZzLKcDU
giejB4DabfAwW7KWUGPhfrskLZxFbw4ZyyiPyI5bqvy7w/v7uodgE3A3HzZ5gix4
1gXeK4EnvLU/RIH8mErivSkOqiHxu+QCnjugpUW8l4YIMqVKZSLzLDMBMyovi1AF
DStfYTsblK0dciyNwllz9vEd/txpyMrYsQal9cUZ9SrAkNhqWx/00SuBHFuVq3Lo
osQ5IlS/zKL5B2xf4p1a1KcHJnv2HPDx9gNXx5fg6oHiFBAQLlLZfLNmJHxvvV7W
X2JkIkljXVnnAxqa064S+Hwm4pSTk6bXQfR8dfGJStEWCAsW6Tg8gWEAxT7J3bnO
xKWu88Djm4Ui+2uHjil/lu1gGUAwptf0rMKjSngftXgo4F7hkR5FnUYGWl5R87bG
42D7xHlBbPD5mB41OQhMJiUlorWaAwbMPHd8euJKSLmuqAAm8HTM3eGTN8a+1pnQ
LiOHFDcvFBsCszbB8/FiEG9pyaJ0GGLgTvxWI0zMoYwOxuIZ97TNTgcix183Z0tq
rSbSGbLyS03OKrRGK33LZauuB3k0KG9csIbmZpdtkirhKJJrHTAUdOFzdMMC0PLu
5Gdl9oRIqbryggcVse2KzkNeKk24PQVV+rPlCDPmQDGH64B/4WrOsxnYRoG/rSJF
G68NAWCcYKIlRWZRUhzGreScy9abtw4mnZB8GNQxloYxz5dwzkAP1Xf2I77j0mdT
KlIJglY+rEIDXhiOFKJyu2BDCTR59iSOnp3DuP4J7UVhuP3CvhkjdWb8CT1E9nTt
WwyjUpuPtJfiPPlqg7H9wS63/MEz5JlETxfbPneY0yUjoo8nwaOKQFfQPrVelJAI
lRTTnXmTbgtuAdukQosnOQkWFdAmaEkzAGVj2A8tHA7Qsj1RRJsYx+JTmaXjyCor
c1XtBc8eW+4ykKpaejIMuy3msYzG5wvs86uHEtjLo5+4WQk0uXyJ/Tqjhv5/thhy
oBG9dkLblBLvbinU7tm01Svawsqv37vMst2g+5TB6vrBIIDNDyVrQhy1DtZRRKfM
E0iGlSTwndHqukqh2RJJmjwH8v/6qKbuuqCSObOY3qj+eFiPuTFku9EHoN/Y3iZl
9FtAvkSUd4zu8M4FuJYNPfQi8AhlGH76DaHZtLm/48/kfiMNz4+GE/KMuwP+UhFa
zPqTxqj55UQ/z5g66IAGeZawTLNKqTcgip+hy8UsPKqUSu0iZ2hO/gYsu9436dU8
Dt/cm8T55p1/lmk+WuKP4ikYypLRRyWeXS257bDnEzR6butE1SRTgdFG1T5PL7ed
HdcqkKdKn2beaLL+aaz2IzGxF3gI/7H4h0x4SMij2lSj20x/jXoLB3WLKiRkPkxU
fYrgiLNfPXZDRYQCstulD7gOiYCxgoswQYpqwHMojszKHYhttMNhJKPFvjgoYO9Z
E7gUxTVC9WwBdr33eHiB3v58yyGBmv9yPK4ZYqxuPcBO/13X8PI/vKqjDuu8/pIE
WO6jBMOKJxzednBuavtIrXKkIBdhOiFOHZ9rOSauCv4w7SoIywdaEXMbGrbvr0XN
yXbvJDehKD4PwkLusXax179gS856UyRBh+OK+Zu8xpPL6hdwD9RdEl1OHSYQJLmx
MeJTRVMsDeLQNw1RgZG4do3JNq2z/4iZLtI5evh/Xr+VuIjYHVYA3J7oDs95jQoq
i0VHKrU3S2j6fAGB6aTepNtFNGghqmcgx1tjfnzU6yPUBf5AlsVkt8k5W0P56lof
Fayl/nles5Q11GZ4Uag8nzMUZgA2sF2UoXZ3aPXhzh6RKz6J3ujRg8ZL9I1AlOE4
QY1FO1W9lOc303cBN6al6gO4ugMIqyHcwyVc3UF5SuV9vdaQ4gu+pcRwTq5QC4KR
EHsiu89OKoZS3CNZIDzHfaZJ5AQxVioFZvTNmIARhmb9ELYFXv4BAC+wMmlqvEUJ
DUjFGUlJ2STSjigXPMJaX6PH2kBHFot6paRZpGPFo2qLuDS2cstPCORjbgAUjddb
eWEIUo/inFN3lbJWiQj9cjD5sGvQzWreNnwskw1yvN060Vzt0Wdmn2oWYDIVN5+G
1XRqu+5g/PGXsfrcf9B0xPVpgwiWYKmB0NdW3o967nqsWKvUVTFTSTaSxXN9YUgV
Dnm8JXEA41db6i3Z/AqP7Y3YgQC/URZZb9sjDPkmn5E3Nn3FS2ZCaaojFvD5OHPJ
wC2/A2lgbZPSZ0LVOLTrS2bfV+/1acmthq4nYm8/5q6obLTfXdTzTfOqlBwGCkqv
yTbFTkPq2VFLDW9fU+C9veSOGMahW0h481xtdbX8YjG9AjF0K3U7QoLbuDJ7hReM
45Q308Zg0eOuy1xlSjUIpV1LZmiVimxDaGleD7LkpwpLdg2r0q42sGSyuBIRrDPL
yytSByagUeHLaqA/SP00HQle72TvarpwVLxzVRb5exRcbGozk3QbawO67qSQYEqU
iZO5NveN0lJTjSH2N5rTKy2yE9kdmcKUeju9ux/wcz8zIiQW6pb9B3mi6kDTBgGK
NMVWuVm9kqPW5RQmLQXpeDVbgUO6GqF0bvwK1effgB69rH7GMd+zzPnsZlOi2oC9
AhRtFxpLENU0kBsSQOInjdtyvI+1HLrlsxmFCoO8cD9eVIk9SFir5mzeqMqtgC/O
cMK0AimwuPJpX9ccsUxStZ5ncu0blwtKAWDQzj8l8vdwU4W5Vcx4tcGFOdvpwy8W
GTonywcoPfmdJk2ar7FYu95nJgAlAFSAUCnX4uYDNKzSCbZWDVFyYq3UKNW33jwE
wUy4dW6OSgT29P+hfvfqjsWFjbjcUFfRor9kaNhXHOGo/xV1oknb1pPhKlBcUaJX
z68AmxWBUbsA47ujC+DLwZ6HWp1dQmmLIvukAFhUoBKqcvt4759ZJ1b/N60UBKeT
oOLe+8kmxHLse2EhIQnJl6EZnZ4CupY+7EVuBq3DtxWu97nJL4bUBTghWpoUmU0m
3Eba/XD4peSJnSCyfdNBTBWAHgOWUP4/+E16RJ6kLHkwCjasYSye4WTOfv7AlPDI
V7s3Hoo0l62LmwgzhwTut+/rEByhNMAtbMCA+YTPMH5nPEljQ3cRKBzzL6LXtE+d
9b9+DdQSsUtPZRuj2UL8LKsbTNJpsSu+e2vNR1naC6WCkPPoexHk8FvGZc174mIA
P9RyVed9kLG9YVZW+E0GPlR7ACI/US5QfcxMogLk4F6LonwgCWOz3rfiRri1CWlI
QbeSaxJkiq9fjZp5BpHs0Ht6fJxrdqUN7VxgfNVTawbNson0I4rwl4v8KGBCUPVZ
PIGvc5z6OKoa9WufWexCc4oWtQ+vZWPvAtVENuwkxAIHPjH0JHv6qosghKsIDrOe
gwUQsK1KT6nd0LuqGoqetvHwLB0zrn2f73NpagOMHLMVPgHSMp8LRaG5LhMft96x
p9IphBSO5hf08Bzz7sS3JT2o+neU2APNLuTLYLRyOQE3XQtSUHjkgQzynoPjekPd
FGdBeKli/4cqH5eOdo6hBv/z0j5tnqR51rT2kqtz/Wxor1/QKYiiPJObkYp1Mwsa
zfZGVxH5h14zv95KOa6VveVda8N2cFH++ss3h7xLqQLe6BOAeA6Rxbf/KSCBnr9G
KH3hoI8fPnVdwB6AkW/fuf25XtdpJn4QBQfZQb+0do4Pftu4ot5x7+yCdfyiBPDv
p4J1ZnkZR899LIvHTLMQLgqeAN27QIzHHALGV+gNORd5lsndAkodtIr0cL+oflae
e8lkF7ousbD5sjModvjjFg==
`pragma protect end_protected
