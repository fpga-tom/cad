// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BMsvOBcKfki4C1ouAfmyeOmddwtGrTSmfMYSyG7N2G2NUwvopyylMU4V2W4Vip9Y
Rdels1vt3Dp541Q56wmioyW3AvSGBkeQmm49oT/97ILZ0PdLMcKQXhpi+KVyGN3i
qWrJ6itOjyU+jpFypWa9e/XEDW7FuciW40EtP7zutMA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27696)
GkxIhnoa3nVE5supu+S5jlAEsPfIO8DUIv1f18os+3oiL+GhRnBJXQgj/BdH26ii
82XATneyVUTJvbwL6iwNooMnnth0CiODje+HzIhOs7fsMUR1qTSF4FNVi5RnYn1Y
W6AiI/kYzYfSETE5zuOwtQqcJhIAs9DN07iXcasW9D2M3Zw4k+F/HKmUEmQwlzL8
+dKtZtBmnIAa/M/GJJ3+VwSH9SIrOwbDZYLUei1tiCtavz86ROw0NKglymCroLuz
/OxoxIezn1+wfdSMx90t44dAl5TTeWPMxBM4IQ1nkJxUgHfNqWAKSbS/4AXsS0Jr
/FYHU30gDemVWmwYxrrE3QddX9J3aVA8Ezek4yCUmD9/crm0poMVxibuh+Pq7ttw
Z3cBI4Al/x2q9mGyfoKYVn4pfxzScI7iiw6AhlEjAu3IcoTF56zsoiQvPg4eaJlN
XSKlOkAwWRG2zk64k9oiaeZ/bMGCrzM4lXFcQHNCIWiPJptLqrCimS+jnVKwr/e4
jsZ4PdxuqNuJ5ODuyhUoTrrDj9wisQNxKgbSHgjTNPH5XY1xrTu25evZA9Z48YR3
CGBAHcA1sOhc220hcvLDCXJtrCYODyfMX70GTWjHGAsD80wYG34jL+IVx7dety6q
ln+Y2Le+SZIwSo+atPD0eZhfB0PEJOgRZK1nS7C2vKExUxfdOmKB+bq0pmBMM4dX
ASzpOVrjkDEvQx+ZmwNR0kSErCqqIU1aFTsAGYBppCKZqh7d9PtlrGfO3jHsdWLV
FkbQY1Sw/v/zJBuSxj3xMrZqm7pxNYAt/MZHjrgdqekzbEpkN9fCrBjVNnB7eLAj
JMtoJpp2tym7FFpAVte8jjQodXaD0edYSEoBmz2I9mYGJeB8o/zZvltL4IQK1jw3
+6MvZysMiPU4hWIjRg3l09G+rvAqmzu8M4Sz7UH2U9zvaY0aZxgEh/arrL54Gh1I
U+HuBhjzHM/iVYWTPf+3k53/6vgNCl3Zv7xEzkYEElhOfrPX9yWoyx/2GIhg8WZU
/5AV1Vh3AlhgYAgpSKGgCLTUY5Se/uNIjv0tFN51hn2g8v7TXC6RHzOHhD76ty5X
uadCl8PazNaSvAgI0REIIbnNvcBgbjz0DTSzZ4JJ8z966LbDghUyJBM2J+mrpGUp
Q/TRVULNK98NvnSoOJlAzKOXLOA47qcwUMwaj0GbyOQ3Q7UEZfFymy7lWTCI++T4
ETMhMK+9EqYjyZkq/Z14eDxua5pGF/9/URyapgvh4J8Z7cMlSWs+VgXHdlKD73nI
i0psO+OdIsD9j/AHwiJe4MfdiC3VVl3eQ6xrRJzbYbyO71NG1o6FE4zyPERGvLF0
JyF11mwp/hQl2Z3P+rkuVZZs9cLL+Hck2QH6O6YlpWG0MvLT1sDY975mp5CJ6Ror
wPhMOLwM0EUlBoXYwLaZkVetizD4YE3ifYx/c3acXyyzn+1L+F9rUQv68+3PISvB
8D19acY63QuO7Nv9n5OzX3SLA3nmAkg3q26XvyF8qlFtGNLx9D/AZZi9KnLHwzyi
TUYMGmU5sjxBSrt3vfalCLSqXIbmR+YEDKUhDaH5UVbb2+QiVjdQMJ4/5XgGyTUC
BfKLTRG0rhAXHCYhj6Uein+P68t9162KH2aI5oAE/xLvSd+QSsV8feXbmUtXegoI
Ngn8cNzIH2JxGi9ifag02JHkGvXaLm6p4rMGNlSM2sRrY+DIwvK3qkcp3AatQ1Z9
ybgddhNzlaiycxSVIK25b2wpVatimpJhytXwqVn0qD9/CeI7k4QJZZ0aQyVQdCtU
htn3DxIvBRwf0sX0SrK++VbegNvslO4Vdc0GcGrLzJq/Nl/lJvscAIgJkxKEpdKY
VcQbUcsiP1lOa/MlWsbMcDWzwBoypfk9nskFrv5LZpmJsVQWKwAf6cfpnFsV+Gbp
TFhINHAxrF/UfsQCdub8JImIv8huVaUjyZb/86pVqWXEiQ6qwxVTvvxJz0sjeErR
2AQGCkWwM2zATTWDQGf7Y7lXRCfe/KwqpIdJo0WGsj0BJ6OErXDcB6ecg5CdMRGP
Gk/6q4/2y0SFEwMpUYkazWlDT8Gb2+3M+mJUtuVb7HzPBxlx1OqST0eUP/G8+U3E
pAKYJ4zxvdSAYPeP10qzoNj+vMxYGtwIYtjlxkhTBUQRDokVWSO1F0G02/06olPS
fhxoLNmY+qrKPE5fDApkGglrqzNbylbO7oxgJ4X4MjJLAMmFB/7J9+UufoqH0U6Y
vRq0wADXKBkoh/KNmEVYbf5sSD++IUbav5j5DeznN1iuUUhdqPchZu+JphZAYnGR
PbI+SO/cn7xWE0yRBcEeKdLfglh1ni1MCodad+JFD3XpH5PDw511bQX5P7pVaghF
lnRMlvfkIi2Bd5KWPK6nrv+K+ZXteae0rHekhJcKuBdP23EsNWXu25Gau0LjNvlM
I/rCIWn0mV1cjDIi4rRTK2YqtIL0KYCJCYfiEiKAOL14tRUpI6iDvMpDQ4OCdYxI
Jz9gixlD9aqvdQD8xNyc50tz8BjUvaUqCKNt/OTVfrdWgHvY0kBnt9T5uNmHfemc
GYbUWgx98drkMKP7BDCQlT4w/ainhy3P7zzeO3x2scIwV/USyu0fImcvEuKRlzdT
Gbghoajo2D5jS0afjyLC1QdTpLW4+yhUK9n4Wee0SrOAYLL/1dl4xc8uVgClwHip
T06YOjiSDx8DWRTcFQ4qoLs2X9nYY0M1EbhxcOTIUNGI7LkrRFPNjc2lxdgn/VXK
V6MjsBM0yt6dziU0GBN3l/G4AS7Hpmf2FhzrZ7ZTedUT2xo/xIdNC6aC7gLchzqq
WWoVLkpsdhcgvYxBhQu4UF7Dol+i+q6WRifkGiqMF+20YzUn6hKqLE2lNiqKLSVs
4i6IcuUYnoFZdE6HiDET6aoJUasnP6ukmwpC1tTgAMKW1H3hZ46YFKRyeYaHPLxy
QIfAAt2xNpybjExUngWUOMZ0QSMERWqCGns9K8ImYieqyNktvmkCmYco9fua95iV
O03Um6/HFR5PhH8r+SKorilHTxDJ1iwrP/p6iBzbKTnVel6rcaqF9BUh6smv3VEx
douL5w1+TAa5uqyto8LKbXzIq3UcS1EX0ITAmPJ/W0bi74IxbNLfJooD1WXunoxg
kpePojwdhmUoXbEJeKMXtps3G9cBIEib/Y3tW5esOa6KcXNwXNb1uj+TddLQnvHD
etOMsSnHgp4Xlr0upG6JOFA3r9POrixSEt81NxZmh9EKUb+hv/dCwYKdg17YY+h9
z6ZZU4ETNHmvX234sX8Yxb+qaRum+oXfEbAMkVbqHt1GhjG+wrYCHHodVPBi3yE2
QYFyffJ7QpMUSfSuH1qbNU8XB6NjWHb1vNcrP4z9uBDNKTJIl3oSsnk57NxTn3C7
tlN22VWc4pUQAShmcjVOopiq1x508RDtfqxqIu7d07OMDEsc4qvgvUgtaNfvh3+m
k8shPAjPKjxCxQK0+qKL2Pe9+rxdG3e4MkJX/uLr3aqAidF1tBGklmURYyQYNmMJ
OIHPGjBhNngv/GI//LwwdtNtnr8DXg3gD1sDuqx3qD0doKZ7VolbWZd1g84ohRqJ
RlTAlP6Mq1ujmRPLTrX77AXutZSRtOc22kA2K8VrLjqamE9S/OAntgmld4UUuUnz
hz5cNOpuYPA9nZJUGFLR5xRNSCTdKpB6ctXbLmwq/6ziJz/zwSdH83c4wbcS1Lm9
Lm6tP7PxzzW+rJH7y8PbAND5viX+1UCpV3gq/kWZHOEfQQp6dR4uE5ZY54esGBTW
ACcrM2eNIdjh3YwdfJFeh054aCXRD+wlIfpdrMImiDg9Wm4XProYKEups4cI9F9L
C+aFH0Uh0fGu9D+P2cbdQqeUXvN7MdMV8Su+5roE2Xia7VYqYQWxFroV7FzPes8G
9Be/rdLnA3ePF2E6ZVLWmuAL1T1voN0YtVhykesdv5GlPcQr/fgBy8RL/HXuDRcj
slbwYhQe7FUWn8AFVplo5smuICXRJz0XDLEXJ3dI/JgfXb9UxjComYsh2Yw7rgE7
G1BWXaVcJnPaV+iPCKyPwlDvpyRD1Ypy8ZGpt7IaJQ7aBnhayzi/mwXfFbMrZQmE
TcilCVPlIEQTeeUpGsc0VtuMV9pnGOUppltel3iHHbWEaaO56rduI+mJfupsuA39
hsgSOL42ryFNk8+iGdh0Cuv4nbJBqi/CaF2b46ynF3vdEdRUd4aD2pvmmCPUMiyn
3Obl5ytrLpnIO26HzrzK1pBHhqk6WeVVZzb74X8KgjtjfmTXgyzKVzTtf5hef4WT
b+hWa9tcDvuENSI7AfuWZPR+cLK/ikL8DX9PQkOEGktWMVmgANKkHIvYE/L/sHrD
rnBfkDRAdgHfUCAFzDMLGIPHkplF9u3NhOK68NEJMjOIHAmtd9xjn7z+LB+0MCc/
Lc0+MYgDNGi7n+1XzdG8jnS1BK7bOc/ewMoO20fUa4wCwIcvxxFRewXIkVmzEaWN
Z68y4ffxfYnYX7OSBW35Rm90MWmOT0jsxqK4G/1xIqrGNZC6wGC9rrNT/ESc2700
6nneghpvTivRDyxeVE6abenB4DWukX+wqE77Lo1obvL8uxe4SmrwI5WNN5Y4nYmC
nx1bXQaSAsXv/e0U2azDR4ofnmWjUbGYG8vHPCFapomRMP4urP0gXDOCfyrBMBxR
NhDN9mwSEgpI1r3bkca1eEO8PwFoIewCjCWrcpBrJYL8h2IC6KwdioyD0BpUexGr
lDW1T2QWmwGVFblR/eTfbOff1LE9QMlaFdEUkVgOD7XcXmxeUvJV0GCXGDfVBVFb
fx4P9Pq8aTqqv7KMJHSYpBj5TN1TlaM/MFQpuHkyNv8Fr+wCmGMK4D/J+uKTk4O8
rkBLawLn526qIhjV7q9GHWHdkOWoVfSV1X7lSgGuVc6CXSgtNWFT3htijU1OBo0L
UJibb5oi7q7x8K8uporUCPXMbey9ZzvntB+Pu3ZXVqWPzKYiX2RLwORpDRCop8oN
t7U0a2/fLoKJTTzfvRQOUcgxYBXvP8N34o7P03y4AH5RgphfLLCAdkx7AVLykkVv
GXapJ36fMXd3Ag3dC+xD+jx8CJO5yV87ntN9P9udoI2m0ZMDERwyBnPBjupAD3kQ
341Ax1lGWgBgsFNBHLxdItxB1Zhu5B6054LpzZUbQ4YOgJbPP6blV1HNi/oh5TtA
KFFl5HYvztpIgdoKu6gd7hIyhrA9MyEc3DuOJdhXmNARTxx0Z43VNsNN5r1kJu73
bmlRDIrIthZYZ//lcGqsQndwRxXIYQIn5gOmqeFTftL8v/aUqSjq5d5JIvwfV0Us
ru6NQYB60IldOQUBtexiB6QkOI5Ypymg7/fEfyXY5T/rhIvl7yKK/JnMnCv+AB9E
aGINBb7F42e5L66s36wxSGjMtGfcpN7Gmj4CbggbYYh7VkAi9jvAxk0E03x1hWBN
DIpenGU/it4IYWZrb3ZDMCVfs7FcHWa0MWn3t/DOaxIhxXqHhXnmsUnEJVZTSsX7
N1/YH6mKKb946QL0/ryoyfKn5gcCtJD+IkDAetZueOdzK3R9D27N41UYdE8MQOrm
BK7Hn2kwdIYTw4WvLsxGSQKZ9z3CIYd4XUkwRUSb/4dxWK8L5E9pQdLOk0hRQ+ot
QXhJGRdTcpl5KvMzrNngVhLAW1c/DI2qAq9Dok1UDtWL9M19KK3+wYlIlBJsP+1z
jEwHR68h8m8js2bl44MpEPBzqqnbQIctI9YmxxRJUYAGubcqspTfjK+EVg4dTRJG
iFRO9k9ojo2D3RDUzIedyMrFej+KPO5ux9sJhR4QABxYRIgv3LZ1/Wb77ZV7FK79
6LnjU+D28NU1zq/5HqgYRRQsUeRUhUdTGzBg5BhJm66++liAjhH+fJacpl/5Xrfh
Crx3Xmbt8EQbXjrAaz/LL3MvtDiB7kpm7K9Nq58EucmFPCkV3y8agsStxQjWlJsw
nGa+NDC/pkGGM/sr+KkfmMlla4h69TCRCQwKLy9lcleLEP4H0M+WJKUNIqvYvFJK
CkkWat0u9NNXbcgwSoHOAKUKP0kbxvBibDMOdUVP/JtfFbC2kBW8hGI0scTM+oeb
TyQEU2yJ2dcNg21rA/pFRg938+3bb7FwLOiRcG/QNKL03/o6DhBXewxjstv+983x
BA2PDGoX+OwYb9e92Wh9ODKNJsiGiO3yFOtJAPWHIGHA4wOF8h3HKFxQL8f2zSYO
FJeCLVGpHVezeknXxjIo6O+Fbq8DoxzG7d98Urc2wvcAVkXQpes0JovE5qD3mkp+
TQ/vGdxgBRQcNORVcPA2cvgPV5hC5KuclxAsc1uJ4038THJjrFrjwdPqMXQIrQT6
Ypqm3nn45jgVmfHee9T959OrZUMW0ricWkYgpGJZGBUjQINMb1khAXUp89AM8NZO
pty3RWy9aFEf8INF9KSoQn4kA+0PvMpr4JGQfHiv2GFkPFHgotIeKowbMmAIT7eA
Q2FZs7+0u1+6CG8w8BLUT7KbXQgm5oKIO3P/sc7FAEw0l0fSasgVpRM462p6JpTf
WMeXoHYlq2gUFkQkbFc9zrgWMIYYHOi+HjFqNR9M6kyPaZL5TPBGJucUJ5mJlRr/
w9h9PFmmvRIjpkEIfBMtsHjV8slDUB/JjCTDHSYxS+gn7Aon1OMStBNn5lW68Y13
ACnTpIA99NrqHJm9HSozl66rC1whYkRjlaHnyLZsh797WzmM0SRlaQnqbZc9FCPw
oMbknhPaYV5h14TD2GQT5oUc4dQm/osh4s/ybowBUfArrJkE7b86tH3BBwqRN2Hi
8pa0XQKYv+lRixii0y7dXDqGR4/orKLpasW2C12ZHjprTiBMIRAChEqddWaz9mOF
A9Z27mVH8KF0X5z8uPpMycx+O5ob9rk6rofqW9fPSqybLVfns8xR07Koe1zbuSq9
ixi+psWaZcK6QpTnu3vfdH0hmlZQ+Esb3FmFgqzLXoa8T69BRsCQh3aYn5TSev46
pfR14aTY3dOqq5jkEDrgqkQXbHt6tyl9CNQiRTB5ojt7sQ5XVKmvfxcp6VawlRnN
XDQq58u5eRoJnx4t86fwJrm//aaRqjKK9spJ+YVeCW7D1qdpHV526EcILhRhESzU
kBe0Crtz94hB2VI9BDlF6VgeUhByp+MCwnNpi6CMp+5cZpo5cUMWMq7j+J2IdOfF
cZ5R0wlTktpf7nCsR2JC/ctoFmCTc5kNUv/gufJsiWK4SDcTfQ0zipBF4r5fCi1D
PnCZdnkrgYPoCucIz+Tzcpngd5J2SN8ptENbvJ09FDH3sHvMl+Re6URzGpElCIts
uYT62R9J36vpPtpVfP6BxWCd2SDWo1E+oTD2Fkl50NX6UIFc1kNHu1+bF+VwNmG0
gbszGeCyYr+QWs1NHlpEMcPffmbXmrvi2IxcV0HJiT0rZnpQblP3HAH8qPLMSWHm
aHymgs/GnN0TuMrUm/Sv5iV2B4fWqcU69uyiRLcYOyi5lk1UrY4/1GunlH7uQ+yn
EIhigjg51ylnsEknCurRqAvOz67VnL7lMQxXUwrMGFLTOWcDqTeuJMODF0aWwWBj
zfZBZxi9Iw9p9Hh/QkFFC1n1VYMhU+gHWpD27dPF60QRO4adQdGiKL9Az3y8J+Dk
kV7mDph91n6T0FXmTR/NPCCHGsUYItFtW+6lYQDrG84XqPbW2GjH6s/C1P+93u1l
rBEUrKpuC6Sc5RWgaLMlxGMUIvvysFsJf22H1q/emK2IoUs3BQKVTp+Vdqf3ITE5
tkkQXnnWapNrM6qugPX5eAUSfLCpzKy1dIuyLwdwxoDnmPRPuxzAqtYPyKB2zBIl
cXjrigKfElOFzlAHl2XsnPcY+PAdiTu6bOAB4A8vwQ7ElvxKUotyTZjp009yhlv5
pObOVEQuzPFgn6qZyk1k43biLSvq3UezE1rSzOqsu7ildZEwHqF8oxUolQucE5L1
vX1P0te6yjp99U30rrsizmvUvzvBqsWVJ+Z1nHD3mJ6Tk7cMKv5MsPwBs50taYrg
YkvFt1t5RYzFkzNQxpVnkK4lStQKO9fI5v59P6KSP1dCP1RktzPw0q+u/HGtAhS9
mVModbAYHRTrSmAi+mlfI1fC0octZ4+PVVRhegR5bSUmJyN8c9X0vhb90KKSUcjd
nNTV8pKqgVup7zGnJSQs/4eSvjRiojvsUrkAzALU2jzhJotWczvVnY+4vsrgBD6L
U93GBv065KnNTuxXJfxXRxK1jNEMgH16KacdbGD45TGKJcf4zhWgx2rDh1GfCQ5/
N2BPfPf2R2Qb5rOOc+WNwljeibVGbOuM1fTCG1l0AGqk0YCFCNvrzRHsUKjzRL/3
MzkSfTLwonqG2ZmUPJK+5LLbb4mZBHgpY/HeDDf+bzuIKFSANLhCU6oloLkeMDtO
e2+BKydb5qpWeh+SbghyqOBHb7TRHBffcyFGIUvIQeU7OFG+5mlvmXUcVYqoS6sy
am8pcOrfliedEI4eCwQM4muhfIcf2P/QIgJKg7zl+cJ6IZI62Xmz1X107hTOLn5Z
+W0Y53awJg5QU6Dl2YyjaKgpsKAW+JI091VfSOVBsR56Gp+ekZE8fEvEaQ2rHCTK
FiXt6jrQOf7z+OX5Zpr403ySjblV73mI8sgqIHP/a5SDtSFvg5Io+Mw/FAeqWMdy
rLUZHqiO16FbTXiVKt8btov3i4QNQfRwKdQ8LeG/84lIxeB8xM6+zBaDl8uk8MZo
JO9QUpCFIbuctgsls7SThMaDKGPbHQ9Ucibe63arAVp9rUA4c58fOly6DEhICmGT
PaoxRPNinl+WJ/59UM1Zdg2w1zLGBuhkua1B19MGd1wXbaH2zpq7Byhpp29/DWj4
pf//gMOpIUSbpqxRh9cdgSQUAxWeS2eh3b+CPa7pdx33KvgTscHHzgDCrHpmtk/M
+J7ligVQIpfslEVAKP+YnNkYyLoZbSKbvMmpFhuekqwo2vhpMQaAqeCyZO62kynu
I8O0jiB7bIBL8qf6ZltiGQ6BposqwhRKgw1qgnSDSGm0UsgFZs+0m5YV1WxQG8ir
ZfBEi/YLPINZcej5BWNxGuZ9u+wbC5prgBOsqebCauJK7M4YVz2sO7fyhqO0R/VM
ibvnZzbXoF5XWJsX5gIviQb02NNqG3OgsywpI1ptpfckt+IPhNratWmQjiozDcNn
eJbdWkgzBCQwLDZLRWoNsZCp1E8a9uWlxiAYcxTq997KWsHcRdI/er6eaDdO9hgw
FD5elRkInr5aic5SW4//Q4hgT0tyM/EFgWCg7bTuMjIMgipTFf6eio4pGPZ+dlIT
rkwnjsQmehrKrguDohOARhkMEtf/lIAKvBtQCVR/s1N8rJ8OpB0AOCEv3WvMd5B5
LA9i58OC+9KidO92NfgfEMkeXU0UK6GfidFdcBIhilJUb+vKvW5UmkwIeoHLIK/6
1TctqxT9qoMfvkODf9Cuek5QZh1ZGejAl26tnXNRmrSaZ2x7ay51/OXjPJdRVJZ6
d1STtJXEzyegcQG04nhm+70dzoHFI1uH0pD6FWsPdi9vmRCsSZJvUx26lpXZwboq
E5UQ1OGqs5DNn/mFoPN4FFKY5L00uxqvG+ev/7/in5eOFJacCvytb+AEah1OHto4
svaSc5yZRInTxwFiaB3RSoJ2hkcYVaj24tejwQUL8CbW+NYwaumGHm7kkDGKKE8d
bcSZ7WJQ2uHMfQFMYmdT0/8ijjZ4Q23ExdSqaZF0reuaZhgiccS+Stslwd9BCZKP
wFtn2ZCM7ygFLMn3wbAkNn70mQWjhj0bYfFY5GOU3l/l62VfW4TY0UqJMOnLzhuf
usRpMxqiyWYZYmUV44ZooFq5GlEVegPH2+2pQ/rQ0FLEzuI/EvP2p0uKh5JFn+bJ
sqqt9H3G7FjY2ShomXKgUBF/+jubzqZTbWxVO5O227XbsCIf+aG6PyJ12uU0Daj2
xopDo0EKx3U8ZeeBOFrMs6RHo+Jq/KqbZ+U9B7jTEiR4Yjk/Z9Oe4xB4KYNNmALN
adx3Xy+Wvz9FOhfa4ymiQGnQoU0irTxUjZ2QIB+dMK7sAU57h0l6g8NzfOsl5FXc
fNKok32K5y7tsyDvUSb5kEhl9sMy0W+gyHGjz2zq/eYCvKgAM+9hqLsa/PSp1jVM
uhdmUuajJaKFs42WauQ77g3oil5PqgTLhOJebuEfbTKM9m/DP9QqGzJuNwiDVDD4
txZjvwHvI/6NrBqhv0Ug14k8io2c4m9TDA8kCXoyrV83Zlqsy40FpHggpt/rB7Mo
WgGWESUqrU85OEjwPhgOhbWwl6cexOrxBZzuPkXAdV71xACaFG5SVJmndG7nRKas
4x+p3LtE/pnMH4WJgIzwgdrNdFYmTmF6y5DK/wk+iiHPbhpwesK162HRwx1h3sKF
CSRkMNBFkLmJF8qWOdSyhplSWInY2WUnQEKkUj9sKBVitVa7VQtP1YgJEPw7r4F+
pDkoP2wjZ1oYd7hJ8mw0MfGVGdC16wRml2PG3urZQnYOkK5WvEkzOnksg+HLGBgQ
V+bGnee9wxApEN66c08E1KuSPfJnrXhS0NBdJ36b9NaVWel8DSktOtHHRdtE6TT4
b1+g0ZWP2QFi5y1Pe1d08GQZjz5iA7asJWUFJNuJcjGdXe+TKL5/Rvxc2uTveP3Z
j6vBNzYW6m632b721XnqtDBSj+XoeTRd9Ex9o+UIax+kTD4YdWZ3kKKooGteSv6f
6gFTA0Bo4hWKksr1NaBzXD4K8DWBEU/QNY2+5l7ZxQ50YkkCWIlZ6N3T7wB9ExkN
TT0E4Qjxq5YbWvvcWYtNP+1ywaNne+QCsQ3nWPuHWu9RZYdp0TbJUiMc018ussqw
iryXg6j/h2TaRaeB8gGs2EhLoeUVkZY1TWR3EvBPN4dVJyDd0QBixfqm+FH7PvSw
xTP5sboqxe4kWz6HUuy5ZBXsAVWE31u+JCvpp7C8Hj0j0G6w5lq0dDFMWkxQ4q8n
zJkG+EH3Ry7YEcYCzLzZK2RNBREKFVg1mp3Mlg3dHBHbFertYGhllcJlBS4KxAVf
nUxXbthm1rdASmrd6OMwfGia5b6VU4E9VLCgCTYliNzuba2fQG8v4BDV89PHKHcY
4nM4a1ij+EpKINkGKUM+dSE2Bd1s9JmPU+WaHVjj+DLXkU8mwSq1V57fD31B4UWc
ZPRPh8dC6MkAxanheLTX4oXCmbWq3Ygzm7SnoOuh1lEEYpJAzebEeC9Tep3sOSZx
/FBy64aX7TzZORHTwnhELDcFaIG3PpEggehXELuYzfOMpQjXLsBmT+3apPSSJU4h
/JWLjIB/lvlfH/CM0/hAH+MC+a4xgrDLVdUMy/mGJiQ+7zkXylRVL/a5f2D1xAMY
qdkc1cB4CYAkVu1vPmTHWDl+AYXq2dKzlda9MSdiWtMNpsyIR1UKI9SBHObnbJz8
tAGYk8BvOJI7FXy5772CVKSu4AsMoQpW7kLt8GSSOZFq5tVufOJx6vXfQahHLK5h
nodyVZGeLWt9u1SPNm/5Hs4t419IQ+qbZAublqKnFxxu5R1teSiV5ETCv5QA5gHp
JXl5e89PU9mvyGzpxnOdIWg66eab0aKSL5tSlQHPbKGTh12AtPiZDi3t1j95nB59
ixmP+O1vR/OXd485UFHrA5BDGkq6QhSvQ9VenTii735qitooKRJYdksaoo1XVH6E
Us5M3/UHxZB6Pmrepju/HmFzK4jbmQAeaaQWWJjuOwYmzRqfucCAcWEWNsIrPuqC
nE9aSL+zKSgWDGStwpkT+/XXlLIDamh/1OdcKZovfs1Z4aLHpMLG8mz4PoiWqEz7
45TjgzmTumcnOBVo4Kp/gao5gcZb16MBeZ45644bXSka/HNgrZJieqX9WSt07bF6
1V9mhsQk4ATtkIBw48aIv5XaCfYjSjsrdEf1IwYaxbsycxm5nbu4UoQPeUGUCHKX
sRo3xjXe9+q7sMkYfl5+10FwCBBSNcamytNuhsbf5Wc/o4y0swgMdO9wGO+1pvhW
hgUy24O1sjLjJU2G2FZlPlBrIc5NieIOufFxuOLszO0H4OuN1QFHbFP5BaI+/Dw3
A/1bEF+aTpU59nEcptzCjDL6mE88OS1YXlvoAQzqnAolGR+I8apXc9pkxH66cwvA
bA8ROgJHoyjwxjnc8o5xvsiiKVZXKUAqi37OxUhPYmwFBbLyjUo+BzEsDWZcN5rr
VmIIdQA7pO8H5wqrV+MoiDHJi+kKzaLuZyD36FKPL/l3rrLiXNP7B8HLlI7DwAxF
Siff62H6jEuDDFL9Igoc4mJGHQUU9pypeHyp7ORhKUJyfBkAsQem4PG9LF+KxM7K
yC/u6dezPSW1u8lg0SoX5esF19CJuav/7uIDODRWvTWewp3+iqvn8RcQIXfQto/q
NmQdKBg74Jx2r2vTuko8xNbBHF4Yk32qKwCwdL11RfAlivLIn0hSajzfWzbHrmLC
0oR/9P+Sj742uDwh7tPgC1qbyS0HKabkEwGyz9oLRmbMWkytUx0HgRL/o4Hpzy72
joRdJD/X98AG4jPE1wQ7KBv+jebZB+ngDbUJe0PFcnwqxQwYtugBDQNfO66ynUFB
kb46TxE3TxRnf/ltZ//m0Ne6pn9PgAWMIljPdAFnyTL76Zk3sHxhF2E86K6HOOOg
H1lb0VMNBKLcfwlN51Mot1gZ7IYtmnGcYLHcbOGQuZrsVOJctzUjWHPpm8q8cHH6
3e0g6FvT8i+x59cHdx4D13iIa8uNWMEmTEYZ5wZZl1ViZDBPVrRqLgPa/Ey+yjiC
Z7x57RtrZYVZCkLlQGOR2lwozTtGODIU2PhDIIr2SI+rd5tvHAF7cpLftpqwy7iy
NgoSNi7WyWUBLQOCMGqyVDAm+v9kMih9CiytBsuwonUuqNDnDMYb+WTNfKZgepFZ
NEfZ0fcbZFyn+wZLhi2SPOSAw5kGYuMiUIATJpkYxiiblVcWKaABGvbLu2eUUk9k
tUz427vpLXNIHBPCLwVJiK0BbFxSqUxCW30uKS3CBcdcxcpET/21T95LL41Ba75e
38+N0z1LqM6DhL3V4NBOd3axYarz8w+ez2qwJiwnk0dkv5X/87IJhNZzcya/c+Uy
viyfWuwTwN+esU6oUDhj1h0yGAYk7Z00Z9Dv7Ts6Hx1GGTChObQxQHn0cTbm1FGX
DN829Bzyoyh+4LHxwKaneNGveSpNPMbvLRsNApKnGHfr1XbgIT5Lr04ls4UvYCLF
NDtEfh+7y1YU1yANnLQz9ih22hSVqNwrLrv6cDLzNuhZOXdHjwom9kP12fBag6Nu
puXdPyKEl7T5/mX/bhONNVNrTdO7KcT2Zuu3KJT7nNIwwpZj7gddXe4FwAQmE0Up
FHg1h9QxiRq9mTJKewLs1byf/gQW8MN8OaCg21KvJNBMxLZOBDps1ThNonrtFpsm
h2v0vb/saR9QgCJKQAPTeRqfG5tLnHE4bs7A5QNHCfqPY0eejYPX8yMvNrCgOWII
5iDB4+MUQt+Q/bGrx6eLevxqwcQFCTrGoFVaRG8SqBKrDXPps7ijIjBfjFwe2LZM
fFOhyw5ukFKAe+az5t9zKC/cTOCr1y6qVv7x2eQ5t4SlLV1G3QVXb9r6oZaupZUc
fo74PbXM+5YkYU2wUirA0sCRytUpkezlWLMQcbtT2/l9XRuqaLqos4LUiZCSQVZm
h5gXfCqiGSyqyoKRRG2yue1fV77q5kfptYNntzyprco7NIwvTOiSjv5EaJ+fvrDK
r1CY9HBsu9pIluaP8nphFpEYMp6ou7hbCfHwlbtCZmaD30ylRfrQFlr7gqsuGHRr
ZoE6u9Usmt4tr7MPbFpcHOCExpNy3kFc+PyziVnxv0DpMT04Ty9JLY/hF99xijfP
23/iEkce8g0ZP00DPMVUvNu44d6GJIwOPWJDKHdEsa4ifaMD5bSWPuADLBNJ+EPq
G3UpGaGGMlHTd0/fVyOhmT9KS+NZ4BuGfhHGa0w9eairXBmU86dqQ/QN7ViMFjYs
Syr6SUWpHHHIsWuOhB3wtauL2A1YxArCXVYcwfdEW9gSkivuHPys0yL32FbwTL/9
vlRV3GF8kdQ1smLFoUr/IOTieL2Q0sP/lxPENHySNMmeclJ1NP1v+hSD0EKRsFE0
f53sDwjsu3kibeohK7c2fJIkie+/tMyEV+aInWYKuDwiZ/d6A88BpPXyzNz6GyXW
wKJ9aYX3mPG4MuKYGv0/jiNmvYNYia36pxyaw5LwOZNjzCAU18xLYW8uQrywWJsZ
Q1IAGxjSW+7um8L2Jd5I5xTfe8SXhOTaPHDWpF8tKS3Uf+Zbgxhse9W7EIrCbA9N
Cv/4ePBUSOjx+ODND7RFlHbFm1qv5Bzah/oOH2hQDmG4XW6keQthAEqqWaGKxn/J
ejoDtXrr6J/sitnqTtsXNHYTKMfJWECKW+4ufhQABCnpTkiqOVed0k+HkVT6hCop
tpyDN0ffpm/Ys5JE+wr8wxFrVLS2FB2RP0WPbbrSDUFa+wa47I9OCSetyBYudv1j
ELPdydWbuWHSMzQUUS1Atcgsu9GKH2awBMS0OYT4bmn7zgF7Yxcxw1qQXtRk4hWY
pt0A4dW0yx0bWxW+gDN3xXdDskZidLFJEhN5Zojb6Tp9/UpQILK95vJwHKcxKoIm
WOTZ8hby3soXLZRqND2HEz1yFaYvp4tPag/e1dzMGKD3TyInFvaQZwG8QH45HpIo
raxh/wS5rCmtF9GHgLJ3ENoCMXLyIIdLyUt5AcdeX2ncH7LxGFEPUBct0U7MrJC9
sGgFRJ1vIJ5nUane7AGXpucVnFxkrfg5PM8Vs5THpeGMOlzliyMGdn3b9ftsT1z8
AGYHSeaDkqoE4FisItlbrbq1yvlyajTXPH5tyYoT+Plc6QWdeMi8buqkETYhx3Qf
vLPuAkzzwNGxXSlFlpNsl3VYTTuF8oDe4+ZJOgczEMUqMFrjhsazXPaL36saxjcq
DzyHSXBJdr0fBOzBQwJp9zOL6uP78huYb7fTvnbTiFFUNoiBK7RHZaO8DK00Q6Yx
t5rKJ6sBRNYv1tOi3g/I9z4BYPGyLpaqDznEh6AzKs5nPkPxqOep/iijZbKtjaLA
xnBSho+IMMb0NT6XOcRzUja/Y6u2dR7sBzszNzxCiZsNEsL/lJl5POrQXnAVlGrO
yC3xgwuh5FzGgHO458qxyAj7/aGTpoVmhq+cskg5urO5pNnrDa+N8IZroKNodDUN
OSQ/LUs8UEj89jbQCWl84o4pEn+AFX+Zs4CegnEH9mIpLZ09FjNyE0CwoGp6+8c1
oN8bmDrrItWMycGzwlBFha7ZJy8T5ta82J1zKVXhsoVTdjX4BTQs7cF1w+lz03eV
FjNdcAWQ1PYq3BI8nRRqyXkxmoLHgKRyBj4EY0HRzy6W7eWIjpw38m6acEhteEb6
9nMTgM1zVk106b/sWXMUuhzog91dguHEUkdKsmVwP4XXUgcsPeAlozC4l8wVffJ9
Seartkfk+m0TUfwcjRxvMd+Avb0RUvooHCsQtevDBy0ZdWuf72fw7WAN5nBqY2vH
tjduIFEtgJ44dxPM2lwcRUByKGuQ73mDNPfrRfwz1B53PWO6Wms6QQi3zqeAUne3
noNdLaTCJMBT7BixGP9TvYsE3wXDYcReKwnklLeFI6ej4KGaTNyU4kNBZzEAlfqJ
oAPLTrMc/lTFJ02wBF+cnm7vf1Rkg9ql995fYdRYy6Xcn8YJZ/fM1FK/LJkaEs0a
vlWCCoBnIRn23I0elZ1TGBisz5oXJs1CvuxZ71M90CEN9ba+pNEbVMyG2W24a0Vt
Owub1ouOrHGnb0MOUW3wzxomDRfLx5aZiNSq/fgKsTS2gv4TLNWCt4O9CQGPm1nI
rT2isWbO9gRCf8Z7I56SE74WxAOYL2zr5y3J+sToPXe8fMBsr2tUfDp7Ypaj01Po
orqHQXYJX2wa7EEiajCgyxo40qxxZYlWwZcfTn3Dz4x/p9bjcHcA45EZzxruQrwJ
4CCA2ROYQfovNwbBVVFdGuJRBpNStWIlnlUWzX9zzU/AFF1TB6W3dZ3iMLiwfL1s
A5SI+6hNSo8Yuz+HIdT+v8aJce/Cc+BOR+sxeF3b+gEqEwwn9wG9Fl0MWutTsrle
k994nRTEXqcQnfs9alQbtlFTnz8VrHeAwgGVlXqyoSi3PTICjPknbQUw/iEDl41Q
OuenMZO2KVD7gOoYHrvVvoj6MsDZLfVATb/aFfQR/6Suv+R5//0Gje2C8MBE6nUw
stsmFKix+qZJSjUmhxJiMHjL5N16iv6v7fzvnbZO+W+AkWDgQ1J9Pk2cSyczuwg6
7WppJRlTpB5MXIgzuhXihVKU/5mrvwh4ri5CsRRR/91G0fU0zEFJdC8NBR6/GVZn
XMbp3aXf8CE7tkuTI5buxJmE3/maBKnJlAEZgG/JZePrBuObt6wqJ/4CpHeHcIAg
Lo8KTCXtbbZ0PL2MZTBrTDv8Z4DpLXxIRBjMuNqO5Juxh2OKwVCmKA1ZwY+84qoD
saIel8iqw6npf1kn4FWacGXYOy063px7kSMc4AfCg4MQVfENUxuEzaAZ3hTg6h+H
emxpoex0Xnr2opwGO4Eg23CKZhMM9hS7ngRvRqJJlWS+exHbaiFQzPQKhCaCFREJ
LYrj/Ymq7FKv7a5zPaTyX7foncHb+gIxD1cJUd2gXJat8oxA09lkQv2srrPL+kcd
/HI2vjsIpaY/3GTJ8ZmcRUikZyr68fiHLraiONoHzMIFtY37HfGNlT9bIz/CHwr7
cxF7HEcXQZ57IMdO19BKTkM6ogd12N09Hng4EVq8+Wq21Q5vAmMU/U0BlbPTeLAz
xe8jERJsWQdKxznaOGc313nJF3lzxnd0iF+c8KTEuQqSJ0+65JqzAShgPJ+2wAzF
390+iU8Uby00lfCV/JzwOHb32Xx+Eiu4jaxtJRVSzeA8gWdM1fH9GF2VttSAnFF/
Gvrz6YZmC4sxpEWy1mtry80kTWf6M3gVKRshuOt4QQ9y8RoWzYbsDDToh2eidUrl
5SH73avYjndXWFdyhJWK8ylvtRAYr7LjrPHUNJJ6JK1/7V2WBJ24bEYFIUZ68pQA
U7LvTyqJECx74HZtWS0FHUYWMk5mGZSstqzTlQr4XnDj9h1GhgWfY21atH9fZkIM
TgItxi6uwtSSRSK5ZEQwUnSKMSQxA10JZHmeMR/SyJNkgxOjs/iMV/G6VozQxAPd
wFME1zXJFAGQeZwiTI44R1gGEM0xggczaje4PXsv0T8Ih0uPIJYSiyZg+GVRCXQE
mtO4R7M9wAjkr6oJavpj4Ych9J8dFZCz3tgdwLMSZQz6BlekY1Hcs0RHjmioaOMw
9ok5aHw+2xFjt5YKD931MbbhaTlNoFWjLvoxHhJehNwWvGKul1ZUS1uqYYldaZa1
2si8UXmhbsSSLKiaiDcK+KC7MFZ33eA5Rk6MwTMXKFxVjr0NWBn577JcWYBUPXJY
1cavuI20pEqBzAM2RYlRL18vKdUlDRWGSO8f/y2J26AffTUiVtjYwUWysn3Yr6BN
nmmvWX18NPWdAJP2ymzX5qhUZOpUR6Dj5uuHy/5A57arO50o5hUS9DqQJ+/x3bE2
OgmhadKfLYQUYgaJ583qWnZcwp3+roEVMlFTXiHQ5YJuXpYqKcOjdh18y6PB12RC
h9tQZ/a5LSSJ+n3yjkgvPgT9l5jVZ19BTS7NhIRF339FpivDVa3J2LgyCsQDbwdX
XQxlrov3BPvnsZmPH3zCbjlLqXfE+QeEstVj/wNHjXJmiZnSlJVatOArTsfKF+Yq
TSe8D7zzLSyPaSxoU6887FpkuPFqwCWzD59woujty09K+hhl991tQ9mQo12Xw1Zq
IDLXD9o14590JJvqy2ZkvQntLKD7VF5zHqgIF8KnGX35NpodHcY5IBy//KDvtJ8q
15mxuq+XrRmZsYCkbXfpFdbioz/j3BcPf7Rcc5ysn0fPQkVD8PKjhoVGLqtiv86J
llWjmUpaILoadfdnm866sIw9qvdo9/7yA7s44/593rIiOuS1xjKa4dNTzH08kvWG
StxKVrXi2ByThoh0ksSfen34ZOZD4tVjaIiWh1WGqZ7PyvBJiRVvUlt/LCQv/tEC
a7pc1p7R8bdpcNvgMHcDdXJKuDM2zgTCNEd5HOMGFBmmPciEYCcsNdNCP9X5R2Y4
RktlEVLC00uE2HhbvjIPdjcHQ/FTFMED/5DFzCOwyoSxC0s7/ClLGzdbfYSoSsGY
AiMaDCFCtidgDUto3NuME2LsfJDHekqlslDptasyXXiKBguB4Yo7hDvmuYDsxvyF
px9CB2QiiECrMZL8mr8N6Sti9kQ9eL9HEf3RKiLuGTSVylydNmCADwc4KJbfPrRS
xef4oqpclHMmDFlbTfABClA2t9/MVfijO0nzGir/euSkaoAlcmlyVHvb0h6X+PwH
iyhDTgo4K3Up6RsdgAZCNQ0WkgtWTs3xG/bTMNl9G+RDQ9mdFx/qg74gkef0OcUO
y2yfsmxNuh4uBJAnWEa6Q2fazCYeQZvEU6Uc/aHltrGMyzYmHnk7KSroJR9zeBYF
smEa7ED1S3SzBZvllGKk/UrJO1Ds5p5dE0R93UY1QEXeScmkphksZ1sXPAipwJZt
i0kknzAX/okcFStpLnvIb9yxnAArm7HuzNUHJAWTD6G0Aq5Oufaobz2gSyYYx+HO
bc61xaelZS/xdIOTJF50NRWirllfqEl3RvIuEGYf92fU6Bi34bKbSKppxQGVsbfY
E56rQ/EFIMRp7voPM/KB4TWQZIFWV3FVpLEfHbr75ZdL0OhKFVWbCp5KjulyRFDz
t9J1luJNffZAMH7lyBtVArSAsDjZ2plq1iQSKbYCNEBxH/OPlXqdzPkYGLfzeUF8
Y2CgvyfkfCYpEV2hWtz3J8B8Y7kvi86Rw5uxOgPjs1+/smgFR4u9wuXOqUagmuST
vicEpSFLbk1a8olR+fvCSLGfqPt2EWcMUBQcKl/RKeMD5JE+a4IES1/aQ1fBiObv
q7+skgxp1SHYw0ANY1b9qUtPDaHqwLaFdTnjLIb31Norq2nINKVZM/4U2WJV/QPK
4dLWRmneTJL+3fKg6lyo+bBRoE9DLUTUpncTykzFxHWlz/ryu1mKU9rqN+wyVTJO
o2N4LFN+qV0uaExNNOCD/qiDBoJSAFimtk85pPjsQvfalTk5Sq3XGep8YHlcCKRf
Z+mfVjh6xR8H9Y780ZfGlx2w0NXABvAkDD5lJXDfHn1ZodyvjZWuspkRfZCiXB6x
reDsOK/TTm+z0qcYyGE90HDIBrCX0Go/tt1kI2gOqP5ksXPhUz/6eBjospHyb13H
pSZIFQ7SBzqgRHmGindRFXr+oL7LFdhkfxnZRUyfbHeg5F2TD35lWA7qUUl1n0AW
F7chMZU2SomoBU97LIexTHj6FwA1mm0XwxkjKSflQOJWP7GjmOd0Xdbppebg+Rto
EXNEjXVPO+a7ffgRhXlJHNNVAQuNw7anpLEz4e/TNmu/uSoq5b78GjhgM0qCMuea
XZxqsozPpF7wYhP8lOMOFYI5ltULDx4L/+4EQIZasKY4HojzLABCZXfVq2Wbw6QU
7WXZgWzJz3QPjLAcThEfOsyR07sjeBo+XnVyRt5IP+R9hch67FJEq1NQfHUSXjAT
lzdhbWibOt3pFzIFea17Ro6vY5mT/HvXPkEUUJeayIvB4tqmXLzR1e0jLa167GPa
e9c0NT7mYCOUI2sRgWXWTUvyHydd/qowMnLRpIEmUm7SC/jAIwI1j+7ZPM1Qd56R
5k+kueBWMno4pJjGQDLEV0GOnXNqMOehCSaOWWt8rHh5wMA4VVGkaPwgQEai2lWD
VCj1cjCmzMiKuhNAZrQqIQIWSB9lbllkIWEPJBLrFr+fYslOao6uX1kkjYx5TXgA
a+FxiIq70ZXEk9Ce1VFt8lu4J7CwgLYHwHmx1yriHuCjXlPt2N0jgz39eB+oYALE
k7+qxOt4FQZ+RRbmrPda2Znmn5QFlI0eVEAdhSR5mSFD0Js+N3kmok3b8FzeZwNn
2igjJFwsBb4enfQB2v5e8Y/4N6ngBoa70j/lUEDug6wnXxnU16jv4K1eM3k+AEmN
ONzzjqZGOAlZ9aFRiRCLlKOE6/WWCxuIA1sBjw0S+ZU3Bdwc5esTvQIXduQzVD+g
RaMlcoM/KOUU/DhIcnq/DFHZ5rnzGkI5zY4iaPxtgjanTLOYRQQAw/01TEKnECie
RbCzynfpzQltf/B2THRiTq25K5FU6ubE3sVJKkCt4MTPezXemeCEWM7kXcmk7fYU
aOR00pkQbjPQjwQkOUiPZLuaQanyMlMZIYRZ8B8EDwFfjAijTd1McV0SgTQFbl/+
qZNSJQlD/RJphVaqe3KeWBmPmkmgemYtbbyvW0us5Rh5NVNuyaSJMe1LJL/+rAD5
eQrqhPZUFG8pw38yzLIA6Kvvazj/gm2OEdwJhA7vAHODug/GBG6Q0XPwzxXV4dX1
MxVvorN+xlfdplQRlpFTDJDW83vgY6Kw7JywUdBu/tAyxbY+jRyAzMS8Cq/RY9E6
1mjkFFSvRx/uafENfAPRP3ouOCYVScuwzeyWCSunu63g1aN0JkEHUW6ESlg0gwwZ
syIzHVLlvSjGVDG3VAs9o/LI4C5t0nDi88ZIiA3H5RMX05bLGEzzLLlH+gCLfzpw
AcgxXC1soS35tw8d7n2KOLF6U15FHG03OVpZUNPMoCPKVRQQoGEPgi3BF/F6QnZq
8Ukxc+7SeykI/aOH0J2mdSsfJi9JkjBMTuTqPIZETwaGi0SKVqsXD0J9q++Zy6O1
nuk6cX3cGsJ5xKCwsWHRf46Qkea8a5IR2aUvtW5cwNf+1eBtNUQoIAfm2ZvnwYv+
IO9i/x1kzkKqW4CnTkDGRZ6dgunl2zSZzRo8MMlYL/YrXGvhyJnk3YFaENvzk/bY
0zrR3+ZfdGE+fLwjAiuNnFrxIgdZf3bu70SAqosOcGTxfcIa0g1OLpZeN5QT9gAy
YTocYBb7/aDB8frUQK96t3FqkP51hn4/ZL/aoo+x+USHxpZ/8mgL9W17j9kJzGAg
7Frxw+/caBICg5JD4AFJwnrmWsHVvTB/hRbmzSJ3W1NKAGueW7WEtJCMwgyCNxXE
ovRRIuZgZMWs54y+dyNDlwgmSm/i6mVSA22dPofkAihP4KyAdE5ixT5ngWfwwkV1
F5LAXfwy8NDD25znlO9xEno+oirzAnY5i9FVda90UpGczRWPWbXYYUy+0VCUsZuL
cTeP4oTjxHyjwk1WUplpD4GutgHEMboujLuyK/vcs37ewqe9Bs3Nvb89VQVI7LDg
d+qoXdB1K2CjK4ahT8/LiwkcoKFdfCppjLATjdDx5qYTZ8BdiY4AduUSDmWr2vBP
00Ao0UpzmrSNA0MyofVQk74aXPjT8Q38T4L9SMVmRv9avYHSnVUhq5Vdmfx8dVfJ
AHc6dGhtvaDSOjvdHjFSAMPI7XYddVMswMvzQTHWCjFfkS7Q4I1TWwqVBptoMD0W
NboDWvv449S9vZmI7AhZREFXA4rsYW2QwvDpSYZqwEzmWoKc/ECWTavoiHoMF3M+
PnpSx1PIRY0uRd8GNW00Kg/CPidtv5MHL70ZZUD1EANNvpVhcD11vJkcpu/RLr59
aqPucxK3X+GIYVNyLl8hWNSWEct+PyoO5AyOv1cRiJCKmlCq1znOisRrRzpevrZo
FJZv16vhpJFp1ma9VPentuRcfSDpcVBGm3/GC97cSte+/WI8RMPAxrz0mfFW+yjB
lrSqW1H6Bk8bQI9qbeiE4EVoDOF8xV+7d9A8pFcAk3dsGtvddgnxcpwqfXIQleWm
AIhhfAP866me+NtnH0peVirueZdiEue4faGT3o/mGjAnpYOgVUltHrD0S/ZZ0WQ6
8Tg9xJgF1z2Z7Da8b5rojMVTl8ncKu3Y9Udk0eJ0aBU9bhoqpUi4tcK9HWF1HIiQ
O+r0f4EdXsa2/Tj+XjLES4suLniNH/1fVfC9IqYo/trA8nEB5CEYl4t6WejQnFoj
UvRvae9/1DBRcpso0DJxBz2DzHhL1xFZdje1fkFIjHlVRQgCCU6n8+VYH4xzhmGb
lIbSUC+wo8Vd2RCMCs/nltnnCl859fRgr9Klcq1JYP6A9bvjORxx+4Sv6jswPlF6
0GCRfpECaecy8xBtdYqeeIVQlYQjAM//kPPGeAM8tQ6WlZDyECXQspyon081J3Uf
qbmO0s+NEerazPRpvAHfg14jz0bWnI2czQxITU/ANBk5Rd4QiZD8e9vgYfYevrXE
8T93uPhYOtsYP5t4cam0LUl4mNVRnkBnj+i7QXLyhu2IFfWWhGTb5DTkODnn98Hb
nGBbhQFCrDzkkHIuBtgS9KFntUg0hbkH++oda11JhU3Z2fPjFwWOGU85MNPV3mq0
Gly2mXKAP8el4C2yB4ThcE1dK9U4X0c6UPJTUsXlc02sArgmoMIMIoMGjiyCIw+D
EciRBe/tKQTn89McbUfPKAv86TT8ViWantTgMRnF8V02SAv14L6/XF08i5hV3lfa
LRFBoIUVauua+xKesGLwEjrMp5vXlKddW4VyarIKGUJ/iECmPFCvoPp2aDI2o1in
bhtGUPzzdf0Qb/w4GMmvC12cRHVAYL4yMux92zHxha5zKHPQqGXbkou3zPi7T55R
q9F2TQDIf6QoZjLnmhNWCfZpmgA0H77jVo1v8OO7T+ShgEQlAWxUKJXT0W50Ywrg
7e8a/IjinI3AjHRqZ2yeUcvbDmA8Awt+HISkmDTC3jB/jOgm/acZh65d3GhtGf9I
IP3oIDhWOsjh0ppRVaSg1253NxbJbwxqI2sCSaBzR9UciIg2F/EAFmRQo0jzjIHt
KlnZ1rUihkSFPktxKLi+C/U1aB9Bk9zRihR4+wwNDFZKBsIcum7+7odg5pEwUrFS
MCsJPYoHS421ccbIvimaogjjBa4JjRFTuxlURu1ZRPdQQ7Qu3Y7x7JJP10fU7xNq
8NW0FbWO/R3Udfa7Waa2l4DitDP8V8k4Kjlv9eYb1nf07twAuXtY7nWOAg4+Tw2Y
PYhgDBt4Tr3MqWkJnYKHV6Jyi8W3TCAV+j5ZgNuQ8dYde1LYOvYP+FBaeSyAGbT0
AMuCGVbfweJZTmSQp3t44HwPfA760imkhRmaodw3gKaCWLrqeQrO2pblgwScWGnz
QoDDwGtrl5MjjXBOh/IKXLObqfxjPdX2uNPFi+CcaqggC4gI2VkuWSQwlE6odgrh
Axa22fcFyl2jLzjW9ouaoCXg5TFDhAg7DAjIFyn52FZICNnTLBpb7jPnWMXdFM8K
BDveglai7TkJRSDDIoxdWW/NaqDH2WqOeFH8QQDPw4d3cV/2kdDLepNZaGTIPpz3
BRtmZ2BdJ5UMTBtnAQFswchnDKMPmokhV1nkNeWUy+riZG8GOTrFxxCZ4brML/qd
vKN3HisLR11uCWOxHshgXzibBmCEsroSKIbmmJLePTXJJOQLtSKaoXV/Ht4fg24W
1m5pFyZyG0inz3+A161lV/p1SHrQyCW7W9N8vWRYwPoN11znTA+PN1SHuLfTD/0L
VTU+epqs5KwCBV3yWuFLjnD/kgtvL9UsY6BUeAQmQ3bHwT9kSKbyIKOwtVJzHqbx
qdcSFFSig/jjdYxeevEmgOhA0XCZliLoydnASICMQmWm1OA5KEHaMshJvOyr5+Si
VRIjhtZQJ2cnS8+C2gzy5rFCVUBSGYJbWNjFVHFsO6jOjjHvEaDcytRNTb1Pl8Fp
TI0k7YJDKIHf4r5IJanuwSnxBL3IAKaYrViJI+gN+kHh546LOz/rOXos42T73/Cu
KI1OANTOMncJpkm2B499UlyC7AQ66LMVaN6ytBjbLDVdogqTqTnIk2ZHDXrFZn+w
mdHmdHS2dd1x3sbFFqa4V3PaXETDYjI+qYu2GquL80zvkAnUKYnMrPBp4na+CmR5
pHTtUI1AlOzkvecp7vUwZmrCu63q3oW8X6jCIKLXFYLs9INheULy4wJ4UBpxr9k8
nD7M5MSNjdxF0g6uTyHzxAmhIUXpeu2ZoPwDbpOuhyOVqiP+f/RtV+KZMzp59aKQ
cOq0vlBvPEe4RyOvyqElK6PkPyMsv/WDS8tnsQHlb7LlFGGS2WFR7Rcz63ityvex
S0I1NkWKWcFaMEPlTZgT6VAFilX53zuLLdFevjCpcmZmt1w40VtJsoe6U8y5bbms
tQdwhyZ8wi0HtOB+5QoymD4/wLXz2jgacl2KTUAw9Aot3riV7NnwsEB3L9F9RTGc
kTUfxnYIpisrhVdrE8CuzIswbwcQVPPWwXTtSxgK7TPKM6qnLOCqEu5EaTGWuxAu
W9Ws7dch9Fhm5eDcUGU06HV2+aSt1qalqCiei3A539FWPpEV+Q0VrUNJfKgMNWig
b0Gw+0WMEcPp6TFrZC2kd0s9rJcYfaWmnzeb/iJqHLk8V6/YRmRfVMd2Z+tmZtw0
Hm/gNFHwKLXB4HkpXlOgYhGtCfb5i/Yq4eVNK7lUJ1orJy8sAR639DHYrdnBXyew
JDfyr1DvttphtZgO/gVSHNxG/P+IGQDPxSKcqlqv29x8c2WMGW+9A6K61w0rMcIy
Dva+WpO9MKBmYc/aacgHQ7TUoH7LEyaqDRDovh7DxEvthlFDUKq5DN8gdSZxxaD7
tb8gi+n5ePec//ewtTQe6N4nTC/TnhJ3gblGA7sjxdfOTaDRwWqpGQGzdeKTK5cb
UQzEh7uCgFKuvilKyScT6LxbxXjsXLCJNQrI4mB2aosJrWd+7TKnSZI/zy5sOp4q
r5/CAz0oQfGOd3KeUWsK0/oHr0Iw0Zvsi4a4oMCHJi6bpacqzhkXBmYBDDTPpvIM
zFFsEf3QeMDt5KMD75jpoZF3z7VoEadKzetNfXLRz8QK2x91vocjR9w/FdlYalNF
/gknE/SxDsC97XISAgEk4F6kWgrmn9oy5NmhB1xAJfH0q8fKaYRfXcX0YaACVV0P
nRuQrulbaPv39owfMucvpVKJ16xyej4LOGpREDqi+mcryWeWb3YiuNQcpacrbgoa
MWcDbaNh/a8yHyb1sf6uC+4esGHRhZE9MRCvZZz+P3XOrp+K5txPU7LcNhcXJz3p
9Mgouchnqikv0Se+TJMIE+8JlmN2YmVcpSpnd1oyMBIM3HP2pVGYeNbLs7q2thgW
gRuaCsYn8dlMvT2yhGc48a0T+mKMyK3nFZdkS/f7IQmfXLEzJG86EwO9qxY59WLU
bXJRzl8nTm0PZdRe5Cji3mZMCDhth+bm2nBiAaEsMyJLeyCDcEs8YAJ69mWQJz+D
gkhnDMvtSv6xIs3xMuoF36bI/spfeNlBG1t0ADVzrtGlfoMYP8IeUag7eFUept9B
uCSg/MrcYnBGvEHocSSZyOu85K+IB4FDmbfQ1r6b63i1a0iY8dNJQ+Gectlp03HE
RZtmiNwKM7+6wRtdMOWiuFd03ITJ79HJAE6D08SZjSkaYJmSgl0GKyDOKPG5eaEF
QzvzRnxLICQslfBQV89sU/p4wBF3JsezFwic+JmM/MkCmyH2VNXA4QY85/ajB6fb
wtOfAarC4W12AhhV4DMBPXsh7FI7BBOXzmm3eLbXZycTp/JhAJpk10VayG8IpXFm
hQvVVq8lUKp7cPCqrEFb9Jt3OGbBeLmDP4Dr7l4QkMUwjTtcfT9spxBlkvoU5aQH
k9eWzC85ybSRni/+BL3g9WJ/1gKscNOk6611vi7vddtLc7rKN+iFSviCIaCWIXQm
O6kTSdSSMZpKW8BK5hzcvkywjQ8mfv71XY+wdGopX3szOoZU8U6kxkVu9nJRohO6
ealvmWHzYYKVnhYTitwQS4PC5T6AIx9DqRDxfzjduJudh66CByiFq72GMh8xhz48
Nejg670v65aBtDwgrTmhLPgavMltj+yJEW1N1A7Y8Z9p/S9oAU9fv63Qb7RzMHYO
zBFf+cMU+I83KTL02pZQFW4QjVd9Rl1N8oX8xxe6v6vkQHWg65m02jLZRBebabSV
+PVuqSwIcl3Z/eMYNbYxi7SWXzKmC7rnOLzGvL1QuViP0FtBN0Hzx9ouuFS9TpwK
aQ2J9B710AqunkYsFl+MZr+R1XAwGkzSmupvCXVLQqxgxTop14+rHDMKGuW2nqn8
y7gv5K0yEMfAfIFnRL+ge/i5ddu++OmfMNXf03LcU1HCuyFul+n83OUeSryuKToT
Jgc6lqiGtt/nMzjY6YzNQ8HvwleFDTgFdZ5pkNAgfdYAVhnWd/RtR2UIeeHjEbxG
nAo5n0+4GBAus4WmH79CC+tnsvMNpvd0QjNl7bSxYELrMo8rvVuVFRO+iweIcbxd
xWxQkU2Tjp7UO+nljgGTxHl9Fb/AgvqqspY1k6CXlr9scQC2c8F7ruW/d2SdcA2U
W/KJ3y0/gyyNc2n79kHbwKQmFZMxfJsY/ns8I6H1+my1OHYWWYaQZ758WxARWZJG
UgxIxCRHIQViYwr44rfcoE+qBOVxdNFubfGmZyEDUKO0BqFZx8xROz43b7y+iB7P
2PXiWRSedtVezYRsGnWT7hIEzJwLlsqPqCDqQx2prosjP0dbWuuG4GOet5U3sr8r
dPFlk6wbz9Cw4Wmqv2/bhqGflFbCcyawfTc1KMXIh8NVAtEsvDRv1OxrCGGzYELD
SBBQVaJajzZMSJ8FfnFBggQKL/lHqH5SvFuWUJ3sBasiKMUf/oCCtOkjW1syeU8r
k5kSN2RRNc0N6DYAYwIPOXIyzk3Tcmsi1OMD46GKemy9bSEyFzXJwjHLetIJobeS
O2TkNnKf+A+UeJEeUoU3XBxGHFv7k+WrQ8sTMIHNmSCnvCFzhQH8OsA/kxi1SdHl
8Agg/9LorStVyoy7HrWd2rYiompq6vzrx8pkOb0yscAtuerGNeg9Bkhw8wnQzw0/
RzCh5ISUduW1ONvCtG5buD2FtDnsvTIGDgNlPqwLcYPSbjXzbwtEIv2iCoZtPoA1
dhAX+WIUpFxgW0Mge6FnvfuW1UAhrLxHZtjzI3vTEaYcKCMDGQ6zczsJ6ncW9J6H
qHE4iX0oOtWdJXgCwr/cRqcXq+uHrAsz0ARmDARvxIVco5T8bcnU0ixjrVh+fjUp
PuROqpJsKObwL+OPz1t1znaA1LEU2ZgOOcKs8DXzvz9JeC9SnOmwmwRaGAnpAG5J
nNeDp1zac9AF9gK+u+eLlRMEh7heZtpQuzuSH7TIAzRxO5q/KJUW3DMwVGoHwk7j
bv8UhlLg2GolBfi+g4I3O1PV8rcx4Dl38bP+TZC3JsdJK6L6ZRMiQc/9ygD9YH9u
M31QMxJCVVUfaSudFn2ynMEm6l0DtcD7hVOINdM4NIV2DE7TisbcnLxwSBgmOFMY
fykr67QAa2yYGTeBtR1Ny2PoT1ai9U8fwd8z3bNJs46vAvRB8K1mmrkvwlazFInV
crkBqUx4I1FROV0YHhyb12NtDZ0mFB0pqdwmW4xABaugeX/yZk5d8z458FA7C97R
Ixis4I6o8tcA3/8tVP4QpV0y1xbBGMAfYLTs0OTll8Xyfm7WK3K11xEEQJlgRJqt
H8u4lmKEy9Ck/t0r8e2zM8rndv3WPKV2xR2Em+aQRCTAzvlVUmf+awpR4g7U7nqU
08DiWWVoQzK4gB3olbt6oi17MlzCSB8rxDtnnHYQhiC6vXhhBu7pZEy1DvTkgags
F2L0nwUHQq5G+XHNOcAWg+IjyuWkTrYDSqvHGYy1Z6OtlsdPAN+n7BHnMccfJoYY
EtwD/RTdmAyL8q21pblpuJfVgvz/edoNyKh92etH+pdQgso9+iGkrKOWAgWAXXwr
Z60vovQAE8t3aAbLKIaQY1dgVPS6Tefk5vavMvV3EPaBt8TIucwCgwiX6CPEgras
8JjSOKPrZi5d3bc00g4jNrV1erwmvCbLRyPWWfdy7OY5udNDzb/pjKxIwtZrufVs
CqQycG3iWMxW8d49LmmmeRk2llDKaePeBMdVAMInDK9XpsVhA3K7X55XdgM+F+27
vvoNmtIpiWhTy5nHr4XfBXMQSXG0jvm3dyJbXtpzjQFxvp0Vdz3ag+XqqepYqyWE
lUwTOcVE/WHgIkvvSUVXHRIkLNBiAxwSEB0X33ZgI1WCG77YmcfVoF0vpXh29Jd+
373xpGknuXLWvWket3j54yz0tpchkylPVTuRYbVsW40ra+c8VMvJVTT5T5DywEpA
WSNYEZHq+IXiSPp/qOOY9LvlEjM+FF8OewWEFfMeGfUdeT2ew9S4tIpAUcG9jT4x
kZ/S4yYbzAz9hveE2rorm3c225dXKNxlPabRGDu8bxMS1mate5gXgV0DLmclWJhM
W+cxM0oeMWkpMn/9CVI6w7zB6ccIrReRSRDdf5lYfjKCeLEb0q/GYlqyubDgMvfk
r61I+3HoFWEDWqmDNjPI5nql7l5inoMqSYxJFJ8XT5ua3qYayFrZr55EM7Vt5bIM
yo6/SZ0Ecw4XLqHPEV248Lbd8BRGpEbJBLtAmiyayvhS8qRFZD5S9o9wqMXrdIkK
stPXAIlnP0ujvcdvgyYmqEQhuTpSrwSBlDtP5CNY1l9n9cgwmGwXZ3kEDG608USp
4PeUl2JBO5YtfUegocr27ysihqx6Bsj0Pj36+QBBEYgGxuPfJJEjj8allLgR5Ga9
tIuEV014cZks1xJMYh+p39G8VvGNw3oM6fCAz3tY8EfmzvldFW4lSG8Hmz6Ri0WZ
UoqbB3wRjG42H55qA699D27QlLVO7L7qRlfOR/gMwk6olPMA+Dca8FiDiAqHmzU/
KIgg/i0tbalV3Lb0CRUtIg9mFhvKh32ZkdbxYluh3Dl3vl1oqed1sE4w6/hcJp1+
1DO7Jy4P2xl2Hk2orOZmq5wMN+dG0+QWaUcc6AbB87DPqYUry4vyKi4ZiNa+j0Ob
/NYEgI646LAo38POrty/9np950/6cHXu5dhY6XMnL4R7WBfqhwUA71Th9KVqSVqo
VUjH4QtEN8KddRLEg/0k9hi7G7Z0GnBh10qkEbHRc29jv/v/vLW4TqeY/0PdWTXL
NHI3x5dkU+NwxvZHvJysdc8y0Y4hCbsGqcw5MPdd8xBt1nbyHuQYmzZyNepts0MU
nZ4+QhX81v8Tswtc3ELjgK0lRAIPHSMMZGri9VUe72w0Mkd8fkNpVi+afo/Mgm3h
tAHze9R09G3nfvlL+mqLNPPYZ4mXq9tScBwQzX7jh2/9yLKU0rMDLybOFyeDtm/9
+U4mlvsAdmwUiIRAwYDzLCAsq29W76LmhZOIFpax5K1rYB7UppuhZfdRaXNSQH4Y
zIBYyqcES9bD3VzeOgPwuKhvfh+0Z2jxvrCqZGL1/74YD2zazcEjdBuZ2nboVHA/
dzAO18D1IOLNP+6IUEwaXg9YK++wPPhZfXtZRhUQL4eeKlrfEdqsvUbym1bNh3jQ
4Fg9zmGvS7QVI165u0ahthooVSKf1fSidYhm5kMkw3whEvNsB/g6ks1Ru5Luz220
egwxZbjVeBT2oFFZKycV44COIj3JnOtdUg2LLfevRGTRr51VvR4azxl8ZgTnJiSA
fbNFHTRZFhRt8HPNKXW0E/a89P51VXKkBd6Alu2JfEJI64ItvdzctqIIx1EMcrZ0
ciiPedn0ykHKZwsZn/afTZm2FZXceQJTz3QadpeFJbUfdzHoQV79fVXzknGeHW5A
+psQHcNJckfi4gMr4fAtC2Rn1pdIEka/BC6drcr2Nj8qjEB3flQUJaRRdxNHLft/
fZjAne4bT9M55LRnjdAjW/3WHJ70Mk8R1TIgvjxO1X46FA6zlXXzCcAgDjzvwuPI
tPybAVsBDcxMGHp2cgpMooq6CKgnnQWOJaF6ACLRKgCdrerp3DP5lt/Er2IZJYuR
+HAJFB5Z20PisKNokrCMLRj+sOm5lJlyVeG8ao6X3Qeh/uiq5jWKkmL2xZODyX+T
i5SX5cIt1gDe7JrZfbylGmrhZdeu1lJ6fdndUmswgUCD6kTrGfGZZh7gggpH8XI9
kGffdNc6m+UCt4N4mCSMbzYcvFefd97CxWJ/1gdv+yh1Tpxw1shqmdQTCWY2omjW
2L1I34qMToAZbw35qBBNPHZD7CVQ2rS0/ssO9BcaFQUpeR2N5f5vRZIJ/lwX+G3z
7ev3ZVwFWdsHjeEEeoNQsiDAOM759vpipjoi0uAEX83/pYwFDLokRzsGbUnlVs2Q
NMbZyiC1sQTsFViNORNLLcXBpsoKWi2+uq2gWsr2RZsGRuRzNjhLboBVBVBc6WPw
+778gg/i9/g1XHOt7I6LXcwowgLgZteQemd+SZAE5xpLuUHbsmZox0kISOObACI/
LjCyiWP/41g2V1+tIWV2F77pcAwndjDzNGZlPTeYupb4Yq0HTZo/k/h/5lavoLeC
0IajgvO1NGEzLBtWxt/hVweA6FTINHkwWFA6gcHO97YnACvFDxgx07hYdlO8k7Xt
YOIh/wboneKotTUFHgFl+/gAWk8v6D3w8xAnqLu6P7EgAcAws8xaXzK/I7KUOM+u
lG94+UmmovAP0OPAmvr88SORaaNcgUQYJaqoLh1FBQhXv6My0PoAND+AJkz+N524
4CdaD2YyvnT1QO0WDVR0muhxP39jscGraXUH+QhNVXLiyBIlCGz588PSmXj61KNF
d4czDnTbpSTr5EDHYqVZnRoVOa59r7XIX5zHAQQQJLPciu1RAq4qDf6qUXzzB0lQ
Mu224JAAUvoaX6mAflymmjsePC/u9OFMAtbAgh42mwG8Mtf4BQ+hDqIkdiGag6oA
vtigFQ/awsw/SspuzDiv9BnSlL9TvBtoY0EizLzmSbwAy8aPMDgphEusaJvArvv+
7dRzuRtMbPzHAHv34vaLl3hvvvZRAHRBMSFZDU19ixW4Ue/5oDXkOKtp2qzW742o
a8aAlyPg047RKcH802nsjPu3Rrwy4U+qSlWNnvKAQRwEzZl1HcYZxZoaLTPV7u5e
sL0KuIkAXhx7F289tEttqkpSZPuAk2+IEV+bd+XSsHY/bWdIMwwIaNfVQrhmutnY
oWgGLCkcgtjNNEylsLLhVwFG2VhxJMVXUiTZjzH6LW/0+smP49oR+AcA2W+n7TIr
HiWpMHiRqhoQyA0bbDb6rL+EUg/TUNQrWzgB8bmJ70Pn5frqgUTgWsIZSDLAgGzQ
vuSktTcCuOnttYWBPvfqSNiykuKSt51U9GJePajEhMgTNucDH0VBWWp2wbk1xHT/
wkb9PmHy1R7LwQqIOegDP3udyrMdUi0pYRVpDtdUqoswf5mzo0Z0PThDpa4UNLbG
D2KVWfF10W62J0NbXgrEkrhXemytLlCx8mlxrXdrPB5NOseMHqgiVVjTbggBG5kG
zuL+4OtdstNZyzVRJQCxfdVfw8Ta5PBCW4F/Zx08Cm00exwD/9/m/DiS3XBlL6pn
Xp1L7NjK7WGrkUtyrUzhJwR6kLK/aFSeRrTXqct6RgiZ/s0egA5TZsf5pD+OxySv
CoY7Vb+pGlT87Zgnzph/hl1dvZC8rqvq1xcRv9md10oMehufudOBbBLA0HR85/1l
ckLYP339YVVo2xTo3WLawvuMQEf6HrAv2NfBs9P/bQTfwz9GGxkASf+ldd7f8dQr
OUPmO+Uprvf24vCoh2hWglOIRmtgnHuqRiwwwtBL0vRn1edU7If4s7UojGuvsiH+
/vijUWg+RykUwBg+ZjEgRgwWcdjVrn67qFmsphlnf0bPMjeIiFRQSmn2VJ75KFBX
jxRuTk/7k0fmcWnWde09CfMnM/FaU7MXXplGDO5drxnt82Ak6GNzUsyjVtcCnGPG
raiCCA46qtHDicHeG4iNDQaNgQMCRXAHuBPcJAcUvwCwP4vQwHn5gZfmddnc3HPO
Gf8ijXy/C4gtFIFt+6LDS+hmkqfmHKR4oBFRlTZEkmfjD1/Tbya0LcjQKGaqzWrS
b7PfMWrUOH7EyiyJRZhOZ4yrtUqIcmKCwb3K35H7kS9EWBkGXXs/NIYv04MvETq7
zKrLvuhu4WHhma4NKueBrGGQDetL0E63GwHBIVB8y36Km7qemJyyXU2ZFbAKqQ/O
7coDGOSPnnUi/3MidEz/mIvRIB/BvTQvcx2J2Vb7HrE6UL5S0yw/gh0Klx9wf/ln
lly/bFz8da+IWMLZ47UYxdgYvXUtPjSjo+rkkRaW3euAUghyeX4Sxwaagd1qifzZ
s2AZfwKvDZ+O8iQBgIigJO837PjnR0kz94jNg8Fz7z0RyIJbNnAfNfChqWNY6i85
Tj0XJcqXqrrzynZQrcaSgl0Eaw6aHmAkxUR24jZB4TVB+QhkobFu0yBVO7QWtfMN
14e43YGobyws3lC3r8kXEHCE9+zKUZG4hqwc//wzKh9h1s0aOsi3lUiImK64z8Ud
SkBO8d53N+KyiBL2+XniNubXZ7bzoJWsFqHTOh0lUpWdmnczmainGBRJwBNaqg04
nwmA8uiA91tzNbT7Ckv+A6ln4412Z2vkwnQouIdUJ6nQbltgcc2dF/446+xuKOZn
6LEsLZkW+NqwLzE5iilmIQlJi9Qs/rsHJBJR1UN0pAWAWrL42RlKAMgM2x1CcVqA
1ofXbXyuzZCRThvqzayviFKzk0igIV7dlJCyYxkN0m0ndZ5dxaBLHBVTbebScoJf
Brxsf3e6PXcrU6PJZipupvNoRY7xEWvx5aD5MN8io0+GEarXobv4QpnefXLbQmvD
CYTYJ80hGfm9kpYOi+a+Y+o41YhuDUFkKtwHFrlwhpDYofowHoq2WpRSNVr/8Pgh
sYWQZLkfe1+2dQrjJoZyRzwNNg81eG28OXYQDirwNANnU6AirXmFUpO7NfsY8cf6
oIaaxyj0M0e97Plb0+VadGMXvzqsGGCpHvROnAqTqJV1qrUZpcQn+PJTMFkA9Mm3
bIW4255+A8X86Eq1eoT9kSFvQLv0/++b+szX5kMPnMKwuYiHRQZQgAy77uYlb1Fo
l/cJ9bHWOfdcnIczeAVBB3joELAr8D9pijAToDpffssqVftAoDNxt5VgI8my0YxW
tAWind0xCpMR/fflvVmCRFHS9l9gjmSa6xKQAzxGxz1w17wD3x7dABAv86WklW3o
AB0cuKYyJ01JxmOwQglKIoaxpV0EkyF1UqxAsZO1ZhnCucroD85mPrb0l3mqmkvp
eW1d80F7pZfciMvmNf+2mIixRHPyvIrGFtPrhh6FEf1ZXNW4CgxhJeMkDl/3ruZO
diGDz7tnOXN8vB2A6JGD3J575JwX7U3PK5J6gf+WZpI1p8Zd9j2jdOLG+U8RaQCV
SxeRgBIcsXxZzvkh4WFRctntMkcJ0ByYVB5nozhAR9SfaX77CyT333B2uRPq7761
oafgiWb7+Q1TnHp163IsIxJx3/+Ur1MQBSGi3cBW1TEG7odNVdse2PHUrseWPt4C
At8ixe4jJOTBWxpCzvcQ84sgo636W9V/TR4dzMjRDrM5PnIktjJcvGdmJvwJ4PVO
mSU1MMpFOGCAx5k66FiB8jpz8CRmbDBLoiUsPbsmrDwNrjKEL+3TxcvCATkMkiIn
Sy5y5JzYP5541iOrNAo8Pqv+SMxf68BmKtGKeJ1LfxOKdJuRm/jacHEubxYhJUMV
tXPksrDNI8vn3z4wlxSHjD++ciXhJsABX90Fj/1l9mBSjlwtrvuHCfgfVpXhmUG6
FSi7dNO5G4wduYskl7tbBe2US6+b//Fcx2B/8aRQmIUBo1TvN3tEHr+0hkN9wyWI
FXmtLHsTbIGYUSmZKMVqkfpHLHmiw47tkvNAXsb2vDVtK6HkKuB4y2cqLNeCgOh8
sRDe5LjxLHgkcIhmTIu1aau+ClXrBSg3b4HS6zj+F4O7ZCgnYughdhPlchb2fOSP
nw1FGaZ5mue26MnQ6mHa2xCADtZ7Z0sHwq+SycCMrk12LDf3tVSfMZ/k7iPoNE1D
X4kmN61ZmpfWSfYzVSBIjEewtALpnBCouPozrL1x6Op9jeZOxn6iPpSiRkRx3S1r
fr/Uzpl7QwWiatfgEKB7juFEf0FOqwmO8fK35ng13XDMm40+aXga6TDWOIXwSGKa
zxKGfqGfS/ZYdnpT72kDQInRrLw4Ny0BB9sZ4T4/bCELQ4FJa+SHbUxsyebog//g
ionUpZBB1eYOZeMzxmINjYcja3TlXUGy2IzpG83L/gCS/cSTHZ1TdOUzBxjnFN3k
PzX6m8VpQtHEHMexlkdJPQKL/OqFNiUlnv7avl8bjc3W6R+bc3Ekfl/F13uZ9V8D
L9FNHF5+ZZJ4LP4GfBD48ARc0TRxIS7cK76MwI4G2ipkEIWmFI18QQPoAURnn2tt
9wpNh3Tkxqhs5BxJwzZyoQ9mNvh9CiInVp4nhO1wHLHm2e3iL+Nn8z77aTbN56eZ
6MPRSgM41JZ7eIGQbg/WNpAZCG8AbcC+CqInCNSrds6mOPPno5OuVSwytsFm2evZ
BgyFfF+GlAOTOXWUJHgtH+Z6N3lVFQ3unkPs8XWPFV4mOiSYyTkmLumCZaE0YbE/
l2zY9+2FAwEIimJKidRvLEZEVtnCzFfAL6TOcSvbJ9wMm/mZ9//Gabifw9y9LQCm
er4ZixXdVgYkYbIuL5l9ZjvrffYyilb1IEWydFYRRje3wTD7DSNLy+jvUOm+fqNH
5KMbqdJOoMZ6iTTtoM9TDb+K0fQjz8xPWLjp1vkPmhzVoMI9QjMNjY8ma8qQQdRE
Dq8Z/WWryHzNeR5LgmrCZ6Z9XdOOV8JuCXj+GzaZsod/+uWiSC0RDdue3bxmsgPr
6NsdaSZkbznLFT8OpQoGZGOrH2Lo/GQ/4I8OihM2k0bhl5HpOl9fgGVdIdfZWApW
XT6+LMKUqwL2/wK4XXIks6Aj3rDwEuZAapEvfb/ZytAu2c0M46L27zmI+nFD/GKe
TBKevW1glo3GVyhXXvONA1vMdSjK/uYg++aogy3+UUb6t4Hj3fSYKq7d8e7zPXNY
lv3kXNZKtq7k42x1CEuk+JCJdqNMI07dG88+OLW0Sf6unURFa/++DQS5zSoF6tLH
Xz3jMFTpj/BUapv4GPvFJNXGgBQksJa+o7K3A65VdM4IsB0uaLz7rbk16ZLR+Nbp
OTNqpTaKmetoAynF9T0LBPNz97tEmPmW0F7qkkK8jPzSPnwao4xqgVbO1fI/f5m/
eiFCpclNsT64RDqUZ85IM6KePlq+Ju/srDhKjyOovuHhIQ8MfwdO7l+pI7af8cGC
wZQ8XD4qNKFVhcmXuLYv3wSqpCh90X7YAwjfGKR1Y84wLWqWWX4yKbRwljehuMB3
a0hDzVny3jjAOuthsP/MHbnSmxzKAOQgpjMMIT52mgllbncb0X90WALbRcaTlLfn
gDbObGa2I53MJfHfQmO9QehyIfHlU3X8/5ceAaSEXTX8BVass4HxOch7YY9EHHld
5jhgpJcvM3b4PtcabI7RuXlAPTivHedJwfEcouBv2/zFhNrFMtAdY4gTO+d1c/Ks
hsjmLdoIHLhedG+kXeXKNNg5RlfNJME17m401acM6K+Xt6tTjMTiCKNcZSgInRbK
fJkVsdvF0SQEzFF4QwkEhWTcwOf0zg2chDqz3dZJ+hjH3SAd4PrJp1bawKGSll1J
i9D33fxNztFqv4vUb9UOjSPo9ldfYlB3nnOVYhJYEV8AynJ23gYFzau+lh5Nwksr
LZpPXRuo1+wnzgJ4gRThWb2Iv/1UxI4yq76sQbrm/jQ6u8oOW7RKyEDdAdsLcAZ5
cduuMMBk8ygiNGTvO+JjeNQGL4S1OBPbsMfZ0Yu36FWfIqsaA22UYndxVJAof/HZ
SMP5Mj+ls7jT7TNmxq/efkFor2miwfWy6YmXmuQ9kclwHYWNm6lPvla7hhi4RCI7
GnNZwAhJF+wDQD9OBha0dKQc7iqqn/BtTrL2r392eLUCI+93o8AfdOMUz5fEeziW
fM5nRgbORCAhMsphfwyEMYaclOJb94OfLkL7noBeB3gh3DLN3c0LxPyOJQf70JFN
LFbBwd+2Rh1OSksad607Bf5th2sIoTSbZYo8E8e/BGbjci/vQGmu1gPCFweMoao+
6t7eaR+e9OaO7Tifih4Lsw/XZPVGys/FAcStvYE1oE0kzLL83kFwwN3BOEeWgOsR
RAaGTUu8Av/kDFO+AM1fiaIONI5KsfzPbcatTS/ei0qGbKoFE7Ea4pvn52B+6UQJ
XqlbrJMgTDIDyEgs7mSsBmuogbqUd2s1k4UvKkV84xmAZtLuIlEElQew2vI3OC6H
+wJ+rEF+pVk41TU6gSZ35h8avtkPmsCC4yIDvB3okBnjlF2XHNlU32Ykx8DikwD1
sFgbRFI8uSbSS/ziEbCyDFO2nQisTL6F8R+prNG8j8vPbrNkxOyaAaTrO6fmqCpf
UaFTugGqmrSzoOBP/cZv8Tx6VvjGJ4aXzB/TwKd8jZ2lZxt8hwREHmwGF7t1CaQI
2dHlEuZEUBHvKXhx6Qet1kYgu3WcYcC1ukjNDDdKESxtvW3ByucbujrWp+vp8IlQ
5qkcbz10CiKaxftv2kxUi5xiE1OK1kyB9abbsm59Mxx4M1Zu4UDNNbiS+hmB522w
YZkm+SC+1lO86Gb3awq8k9RrCW/jaJSXHDOmwDoCj/H/6mpJdFIXKe31sNhSddMy
4nx9xsNuj99nCNinGy+Kkc/ui6clwsHHvOG+7pGtDttuRMLFDCdy6Gvx7Z36TzGa
QEs2sv8u0H8O4WBb5rXQNczwgqPIcytJfsNxBHClGfUjvTiIvkzTDhLq/9M/IWf6
etmbiosr253aUdYLoyFINxMBD6aGeIC+QOmWmgOvluZpZy3XB/gG51ZHQxUqAmiF
orlOeGy/nQ9EGzLObcKpKG2PLAUcHJOwT4hcJ6k3t4jrIeGLR26bK9NhWk9sCSIY
HA+lWrsPDogdVz3Fv++neyHGsGwOu2lJsVD3HsJumwvb4KQRgzPusTM/IHUdGtp8
+32NYWwQH/MvD6Km2oqdrtvbJ6Ys/QOYQ7v8eSo/mtJc2V9q8no6z4xAoyWTw3pi
Pwz5bIDybxZUD+HETQDFwmFZD2eB8cDukNDMp5zCfYQw5j74s8vIV60kO1xrW+zy
`pragma protect end_protected
