// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
j1Ae/BtRw3SKjTGg7lT7xRj2lA+Acsk8P5y5tUMSbaMVMC6QbqGCY98wD0SH4HcW
rT5q1YqhiEZga3yXi36C0azk68wWygKkQx1J5WSxweKNkzt4wZ9pgL5FHphMzMJ9
8MCZF9JPz040nCz9NATMjj90HIdiiBU6urVqFP67GL0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7088)
dIJ1kFOvSbeXXDoUj2z0nkuI7Ljn0DbNKoNzB2kKSFyLzHfbjNFS3r2r+B5Fqk5/
49OoFPcgqvgVoQ+3NQpqIT7zby5NcMM8D8O22ihfcRiJY971eTjTy/pZDDqaEV+1
4qAJrYwcHn3sNBx+vPF8bdvOvPsWVJhnPtBsZhvfnMmeKZRfXR4oopxOUezMVv1q
qNDOivZlcjUY/7k8HmhR9SFkpifz0OnSDPCptsYjkRHtmAlQ30TXZlYatDXcQiiv
gF0+9kt/7eDYxkEPezg2hPHvOy0ySHr0nCuLjYIVtbHWMUnAZT+Upr90YKSx5AZ4
YzduU6t4p8nRMrJBWaM6vMbIKQXMIMDfOGA0MpndfWFQVMrfneaeF7pSS8PxQr5v
0aIRTt0JC74xJidL0xvtLLbJIRCbBejay8duEazNL609F9PlZSF7kMe0Kqa/JJ7r
s/528L2lP7G+KJ4T8mOLdul7+3wLkacSim4vWuU52gg1vwooVaz2IDxHUU428GS7
HC8wr3AxhnoGnb9o23ztmGN0rENk+DyxS3GCLu3SOzfqI7lHxaQ61xiRCBU0+GKL
md0EhXxyTMjB808WYp8HxMuYYQo9irIcjt/6POh/EA6Nhu4T2gqfL6ktXTIu5zfl
7iziqVNmpoEZi93kTUjaRG3J73CfgcHVLNyBbUqlIUR9K596e9EWPtcPsoZsS9d3
wiF7FOs1Ac37BtMCa2HI3gzqiV/0ANHmW7CJrr+T18pQo6or9tQfqXxRPq94Sca+
w1+54TVwYcNLoZ7GNSVIIYl5oD9fW4EMlRNteuaTYTeCglmjuXFLLnKY3MAxP75o
6kLIVAIz5Q6MJpvJL7c8h/c73np63AF4cjCepvFeTN9Nk8+eabs1FRiZUBp1Yd6j
vT2dejDOqndCK2qB5n6rikUL8Xi7EaGGtqHjR97TARbs7AKz8EgXQaNCTsps1NH4
I5XHTQEoIkMW4jTMarwkjRtu3cSzEiN9nbLuVqAQB7Ct1EC1MFRz2HU2XAD8Zu7W
Lu7zMcEMRYaCUA+BEcKpHzP5Rq5T4dNmLOXTXeDE0mnQPUV6JNAQEb6CgxYQFS3H
4Y+4nj3ptKUHpQ/jnbGFQGz+Eskq+a09gGX6WM9s91x4uci5Z9LOb9tvZxRrNihq
67puelCa2Yfu5jFDg3Mu2TXiOe8Ajg3wrWm3j72J/hSYzppPumI1J6ExVNDNI5o9
dCRnqKkY2oPcgF+sxhP/bRgg7UVNRzesVAQ63L/dtKK1Ki5uNIUr1L2M1B9WdNMv
zm/NsWYFP/ImrIoGgV437Dj4BTriYs98kfaWnr5ahNoQbL8aUrq28xb40u1V0ChP
LPnauViM2n87o0pAFFCgMlWfJF7VR8jbvB/K7UlzDYeak5moRjTPfKTV17vcNpXx
CldVkK1gkW1RsYOApDXsCId0wqZ4A08pTz+P0ch6sduhmogI5jg9zDrqylm/T75p
N5/L7h5fw5NMdxG93qpPOso7wqcy/IPMODNKCn3Rg6rOgfnrW/9XBJ9l6jRQ/EPZ
C8gzqGakJjFO5VlsW+9jgyPXq46Kr4DQgNmbONi0DGED8GcexVaBcblj+1+dRgha
QM6rJmZTMiynglM9thA6DnUoueKr42KV6cZgIVGGDXdI1JS7KA7/eRpeWjDfm3Bc
KPiTqCZAR/Tcl/XyOKzZ+HU0aGTwpQn9OivtDG9kBp0fo2WypnLhnb8Z9ABNE9Ro
IZw3tZjAvl/IyIXMUuKvuurEiwO1dNugr27iWDVRcoqaHLN96aSpgqMsoE5MkV1H
AfHbgEDFjFgPlNKuRJtnJ8D6S+oTcWRrphfowBBzvZUzsrmGz2Y1OZPzY7T+3VIR
ihqTa5j3N+YzHNFkCusLDDQ4wB81fSi24aGAEu+RmufeCm3ZCcc2g8eVUIyPp4K9
f6rrkiyzI2a+ETXeG1i/xyovLiJowVtNZYfhXqR1heBY013VbzqL+ypBEfNtIXb3
/q9a5AqLyBCYZqSVvOeaYm9m8Pz3qBjCkljVTNjE7W6mrN9vZkjjaGEvwJJDPrVq
9+0J/aH9IJ6ZwwZxJj54bTBSwy9x2naJa2M8LWGdysIiVEulVXZBdFVb4DinQoRY
aHKTO8ycpVB18QJCDIaGglphAPNBHFvoAgsXCksIIZ4DAkTyyfo7NhaSVQFIEcph
33lvaUFpxOKApSLgoRxzEUbHjHy7cX8OJw9EZ66Ja13Rj0SOcL1nETaQjU8DpoVH
r/Q25jrqJgGwR0lPUmV0jwVL9/P8FJYlPVGf+NVFs7ZXxaHq8ADjLBeRvAg27f8J
NomwwwgmMnu9jRIJYc76VQMDcItgC2T3sjyU43sQQLoT9j36sUYWKJkxgZHyaD1o
Ctma89NNShfCdGYs3SO+PG+I7EaxkwyRlnHBfivEfZfdeGYX1WNWFsDHusK+kAEP
wsyRsN8ukqrzI/gBKhufO24mJUHZVdWBTs3vjR3XtwQCgGgmN7+ymDnyJbeZtRWv
Jrauzk8OyV8q0AjWyvJQIMRk+L/pYF9zy7Wx9YNt4GXDOjBd8eDOYYLFBz7V9+fG
iP7N+C8GRXV7WgM8y6DO/hDrlNXyfmvRJB3GVMOON6oUzJ+cpZ4DJKsio1brX/UD
M4zkEJhn+jNOtSD2tVx4qaHhBbrNrLqDNdvhK/ifSC9t+GK3UT+3vL6ZKzN26R4I
vjjScZo6V1giqrzUB1UGLY04oU6AkUY3y0pRvWXgEBTFWbQxCAFraBhRVPjOgPRL
FTkT13NECyPuPdFOmx1Kjj/kX1Joulv5MxV5+1KuyQ3VYkWPSHr2/ewIgILvMvNd
TBb+/R2ANoiLbmyoZU3t897mkSFgiPBJGhrUYUE8cAH4XYUp0+hBtHEK5AncgPYx
8loQdYs95WbeMJO1SX7WMreTJ/eHuH+CwNr0c02i3nbQ2W7aN4wtUF3kPKAOoTVR
HGuSAucrEWYD4akwl+jgq0TbgG0OqBBYK/Fw9o8sn36FL1z0ZuSnwtcKJgcUD7Aa
4+worBlUJ047XGMJcLNWlaLf1Y8/vrzhHtvYmfrbC7DWRirV/8PwDV+76NhYUJXB
MnfUBAjQGDv65WZ3h+kNgDTVflPSbGURH75RfLOtXRAr7nQHSx6x+yzX5pro46BI
Fw/aPRRSwxuG1hid2U93JEEiTMZc7O1T4FP0pABnSTIGatqOp0jx5Et01Fbk34cf
gyy8mHlqR8COJCGi0T0x7mGPC3WgcdhVo4Ztlo03DujvjzwCmEFjA4/KV7ogPKXl
SlfTN3t93cCYDsO+C8qeiaWuih7sARipnmNmufrVcQXZ3Bi/y/1AnS5U+Or80AbV
aXbvGbTrq6ehdyx6g1SRZTBJ4/P/BaZKmJrP7oFjlYtgFYPJngy50Q7BvWZcZzwd
fL1AIMGXDL2qANBFwD3JAx1V2yXt93NQpOilXHAjBaPES9EQlK+elLq/ktWChEka
+6Hl6Oj9lvF5s8yqJA7oYv380LR+A4rylmijw5/rkcw/zRwAgxnLN4h/FVrX8lpq
+xNARto4w7T7ZbnJUMMuJklwBfJ5Pq3B9TnB7dNevRRvd10CDMJT5Cyj7sPui+Ku
NFlPQruZDcQj2J1Vml3Mh1T45aOIOn44aD7Y+5vSatK28aCrxpONqz2nqRbkxPD+
WmNqopwQ2Uk3y1FszrGCxhQcMCOmg2GvPg/gT8Y/LZcoepmdFeJNFLKWn7uwDefe
20V+Y5M3fFkS7CcInClHOkQMDMqVEioIBefJVusIytwwSctNiKU7i6bBCn6Gi8/0
VqXWKNKzeOZY0wZme/FsazsOTiDQy2fI6eZ7K8EuNUhhAX2o3oIh7HvIH24nxVfm
g+Aia/WdzxZk7DIGAC1XQ0imRm5SaCgSDjzM/hnVam4UAK03CeJH1KOW5UHoIaQE
IR1P2op0p8OFjs5TVQBHOtWUV6+e5O8t0U/dsmjbD6NUKGBJX5yRJGUXrInnIznH
/xp3fCGDJxLdgC5newp1c9hdqz54VNkdgE04cVfzZ2Yp3A9tm4soyCRNqKPrVaNo
ldCIeiV/GZZ8M3/eWHgBnRd9x3Si0WvvNO7LP2WR/jwVjFptsROfOwUdAENcLtKb
JKwJ8DfTYgH6N8uDoSzQbJMH9DJ+1PyjU4WU4HwEss6oWBpX4lNadTTyOSUaRn3c
FO78DcT0zqWnXymD+chQ4eRRH+3aKp+pLdxP3SwDxcHemN5F9y5pRDHInaX+Ub1v
uaMQtlxKbFo4Q6SP1QawaVu5r6y0YxzlVYaKo4DDxmoxBq4L7KlQv/Hzvzr9x849
UdEnCzC6ns8zHzgnBm2EqmVYVgq854KjFjoDg+rxZC7ZtyErasMAYpCt7q1SILXg
qCZNCchKH0CM3SPzwirJJEywFd5xjf09LwysxwZMGTFvPuIFYyP9axw8whD4T7ZE
SOdDkwynKleubNHWpiy6bOrzwxX+6tjJ5Xm5+X3lyQQhkJ6Yv+r6CM4TIFU5p/1L
Di5imqwQpqShYE5OE9AsNlJ6/ntaspA+oMRSRQskpr2HqM0oFngC2uoA9b5usnPa
wUTFvFyzn6tvPuK6BNQwHsQysTkGCzp5PWNuDbptW/FjGee1IY+oQiu6ynYLPGfT
kGilf/zCRzown5cPGlbYJy658GBmSw4DplhZeyG87jnjHGtLFaAb9a/hoUYxqCFy
3WjQnUxGOH4mKDdF2NROtBgBK6pR4qyZ1AvBubYyaXCCJFDAONaiFsk2BKIQiO/R
Q/dSM419NxX6qY39yFq71alFWMTnN12aaie5ApSCxMlSJ7LPkCJpiYm/XN0chhOt
u8JOPux6kqvjtmK5qyA5JZGbJXy9Lhs0AljvxgJHDi3zYvTc8ZLdX9ym4APjG6IN
yUhgChd6PbZpztA/3QubB+tVHM5kUj1essh4wdohsfpWfJhfSF3adxxS77cG7pVm
hR8tAMfBgJyysQbIJJYtBYV3I5hZAGwSS50wF6yjakOrrHVsIPk6nkUpfCqknAbf
eyvwYfTmuDB5lNiaQuFWHvWP98WH3uyEO0pHngEBIUzzRxBeqf0T9XtL1zfdx1iD
PIDtOBWbke2sk9smF64T9vdvNlLmnLCLRF4AD75Sg20PO6UOh9ruxDGMu+jg+6FD
FuaQHRIUMAXYYEroi2soNpuZKmgExrzL0fLLn1x1p2omnqoGvPok2QktCtsieo+n
D2ik1to03boFq6zT8BWeQ2ZgjIx3mgYgusSd8N69YQvX+dR+b7xuo5Kf8/fyrUxK
0rniuey1or2cr3LSpHlfNP3vQiXqVoFf8I6oGgePC8l4wXMmZenc4AfEua3JOqtL
eKnw/2lb77CEz0IjxacVRg9djGwMtDp5V9nQtygIwU679W57x2x0rrm4+H7KxZlG
NOQTb9I4/Ps938Hfv/T0Nra3OPm48mJjTXK5yV2wZOaK4Nr5QeV13hbtnFHAgCwr
XteCnyDTcf0SNg6ZJxnSfIOHT9kngGVVGPmNVL9yuzht4YJw4DVqH7ALLlt/7XOb
g6+u4OKduuHwStBTwp4SZi6SuyQ5iFoRL0QXDLnXUD09XNoCrHZ2hnyEj5FVJZJO
1ydKNqZDyKNCaIKQ2mdehAST1YnA6ZJothkeN7IPbv9TR8I0g1Bu/fQIq/UFbXl/
d+eNBmhFsD/Y+xjPH8HH+yDGJkiDnp9mUlUqSNddEydtzDSbAN9ND/sRsxGAAxDk
sc7Xztn2fMNfaBq66WZV5xH0lVu3o7NnlDzB71SZX2wZ+OVKhzNpIDtPKXcrRNjJ
6x3yYnpAlDFoaL8ZyvuIVjzVVeCKkJt6q7dRI0Z/1ffHu7e4DyIRsprlfwNwSJc3
C7ZHW1LluYyHgM4U+VjcFvbiDa1gCUj6+xj0poRg8ZHv6K57j0eWaIandqv/3nT2
8hd0x2P63rygLUIDrTJ8/N8+YZmWPRRwn+H3W0B2plWV1Sysp2lIjZuqgzF6OUwM
WnihIEjOsZtsXGpHLZAfbJi7NLXGXKOqWJC0UzUG0wVFCllwUcwraKds4N+TUj2O
xc4T3Z5xQiCX+kKYZxYTxH6Jn9wgX8nfsJHoTAu5Bs3Vv7MPYJJ6xwMu6uob2a/C
tSFKXzgYQ+idUC0kPGQ74m6IbEQKkgctL3pgtGPzSHYdv+6JDoogNI5KtyTOe0KV
9P20w+Zk2nTvi46NXJgNgv5FG6yIhb/r/ryiNsyGmfRhfXqeNDdvhR5lxE0hwotj
GEtHcgCvST7W8qIZMpkWxcrgv5MPtdn1GGBw9piL6I3LpSSMFTbI9ZdH+rUDRsfP
IrGv9f4X9BFWTFJ6xug7zC9Mc/SDCNaVRQon+oiVBsjCzgtE8NP12UzDlOrdazXy
Dru6F65oGaBAwdqmsQEpishaHMdxk6OhZSI+zC100V581EpfpI2jZQ5uB94z7LLO
d0PV1dh43mo7if2JYluqWFJ9L/8UeUL7ffJKBLPYrb8DukpATjW17ZyMpdzjO+zE
ZXEQTEoXE5UF3pP6slb2sFJTqtVZEIsHu8+Bs7faUB7K6BXsxG4CMcfy1PL/zBy6
8AEpTRQKogjHPj3sERiV5GzXASZC98wfIuTmOKPUU1WvTRqaQvL0y82N0MKBSHqe
KOiOYXDkCA8DDACqa2fS6QHBJuVYAT6W8Y1Mphd+Pt3OT4JAxqDxnV6LLwWK9ztY
ZGzj9VTygk5k7cr5oBA14Re5OSFgNx5/5KOn0Rjo4RITkPPNLnwXLyngGyDXHFWO
QXrLQ/fqIOXKhlSUwlXr4FCMAYpv23okzsVbmuW7mp+/MikTdwzDc9r8gZU4Dp/z
85yl2NsqkiXyRxStKAXsEM4X5PYIpgBB2g9HrLofWvnWkao7xvtc83WRBPfyHoZM
hyyO/VR8QNJYInYthfgSsSo5HQqZEWzQJeGAhJIs6P0ZvMVyM6XSSrFu1qUdeMZr
zg1TTK0MhGyjmhi1DGqmxDo4zOyx+nyXI18K0cvP41Lkg7htHsdiPXdGpg9dwBE9
v0a5M/ZvQ6OhHzvV7sWPCLwa0rUKtMZrxWtXAHs6TmJZajHhiMqgjpsNcP9JPA2I
lZ+bPfZHwo29E7RMWc8CObwxNFoOKNr9qsK7VQWxxaLK3vrsmPR6s6jSK3kLVTFS
C8diCSwicfhlXec2AgAWElH5iyilZsCA6JIpml5nLVEg1jQBAg7YtElDC2JJ6GDQ
XP0Z8T7LUSrsJLYui7mJpKRpjK2OuIQ6cIKKd7Fi1vnQz0kD84yTYkz+fuiDW62Q
66QrcbnopfUveF0s2MTCcToArGBArgb2/3J+VnfVXyr0loIVmwQ5QYlWMq4nwcZv
0RP+o1n/trxsVQz06PfW6LVhCG0gTzpVg217H7L6pR5vZg8LWcLBOqAhM6g5Tcqn
PyvWrMBvYMhY9itInadWmuHHLs2CjfOd+8iFQndQJ2Yd/epMEEZdvlhw2gHHuPy8
aBQrXuRmpmFcsLpacaXfKCbjJT4c5X+wp8UEBAmnrRvsGN9kY48ALGdhpVz/fdop
iE4AsNldJUQU3eowCiMjlH+jI9RPD0DS8aiUHF//wUJDRVefA6V8dBL1N9PfVPWo
bEjybPUpcK08ypQA04MyNR0j1d7m6nrjVHkLbwZUZljMQbwkxLM+NLurxa7kVbhr
OQTrhENfHTdzEdZB8Hu7ec0qvPpLpI9gNiU6qGX63RpaEkd2ijWjDtbK52U9MyLn
4rNRt2N+2v6LP7KlV/Ui+tvXmD9e0gLiYv4LY8LdDL86y2iNQ4Q3r2HN8wRn2Z0K
a8Damt7nhyq2QzN5ie6W/k5MZzNCxUeS7nmxg2d3Qhts3yIKC0C5U6r2GVuropiJ
iNEGvXpaMU/ST4dkxm9XNPRJ7BjAKqibEkOoq/zLgevON2b7BVeeTKqeyXgdNEMF
vLU2+giSz5zQTEx/3GhSk8/xU4KrOW75QERu5a46wYNHdCcM+M60m6gWPnulowPL
s6S5qnqbKxsbij5vd34VwMHjMnIPbVHoTQuwPxErcLp+EZh2YxkWjE6R/HLg4n5b
rDn9fJa1iXTCytNsUK5SdWVZtp8OuGKbvZeZ7W02szJ5UoUFGlsJT37VXOyjY465
EbCBiG4jukihawy6N5vpH2UYEkpdtEmWg+KriK0t1+40yx4E1bmZRgHKMcaKkLBN
Z530GlE1K9v4QilzpFP7OT9I9GMeSHdqcTjr+UfnKteNFfO2e/S863oSO/BfUJ01
yAJDpKf+hmMOrl9mhyNwxWoh/znKwPAuizK9uG6o25nh90PXrusHTF19y6yIxuNf
y8a5AqPY1riTqcpI31GBrI22G+3cQOq0DEoh2B700HoVsYmWIOf+SfOU0Wg6tX2e
pzvz5xi4wSb5fOFDfOWFmBokxQ7WE5TugKHWUxmKlHSECSqMXiW2Is5PuVmFdifL
42djtG2whLYY9OMqfCDOI1UfyImAHaCL8IeB7jUdTsmSHr8VajRmSJWSLcoFLDg5
XYKK9LUNznETU/2hN4UAKomNCQmrTWb9QnBF242wNroHrA2u6Oi5Ib9AJ0xfMQAM
QMbo9wCIc1sYzkXgtiCktxB5mIQ2mUrsugb7fadzayRkETA95ArdPZmkdVmCQ6I7
lSCDzqZhHfaQR/D+c6uQ7wNwFRa3v/uoLVTDC0zg7he+5IipriNqBq5a1J9uSApI
/bZPsHC0MEoBkxvIaH3qvrK0g1lcw/ghEE13MEYBjwIrhDzwwwc0o0tJCo35xG7M
37XwPIkIZjP9zpRUdtxpUqz3J0xz+2wKVh1s8HV7kXHrVuP+wH+XY8J8PrXgzIeX
6m9AAvEv5B6HtoYKqqL7KWXH+STjDfbrvSaTb41zybcy0cJG8IsMpnAynU7XM8zn
Dm4/JBu2JTbJHMS2aAS8A7xDnSztzlD0KDwR5GlG8gT8bFwtgXE+y9Q4f9QqJzf1
B1Tzw/TNzTXL5Xs2QXE131NrU1Qw0S2Z9i6qeSoPK0Y8E2WQcVBmDfaoX6+8zVlb
K+62FAYbbuTt05wV0USCnKUWdrkqIXvEM3MEAgPGq7TWZtBnea9w6795GqgYjp6o
GFoCcAvir13DgPmOFl/XPejSoLRvmLe6noN8151pPq/95efJxkTUxQrMqRiYEBSn
v2jBXKjVIai3pPbkL4Vn+iellYaExVNtHHsx2cC7R5reF4hXELzATdOEJdL1rk31
CqeUHBfGvU8jXPkFFlOVhoOWuE+psrIEX/zRyOA6Ud4rqS0rH7BvllZ0iT/+PATQ
W8MDKeleJzdUULzIJzgrzebj3F9Khgc1Ebq49+Etlb21NY0Lil8I0oq031iLsg1f
bexFdZ+2/5l0aRyZczPU5oyfUQ8H3sNo/mAOuzmYLxDsJVblqY5TzMEcNxfi5bdA
MikSb/0eEgprotwH3LUhvfnpfVAAgvA/991USa8JhfKO8bAl32ezhF5g9BXlCqe9
zRBa8nTfkXl/Ey4eUYIRqA9q4IQZxeToBXJr8tNhCA0=
`pragma protect end_protected
