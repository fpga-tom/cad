// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pwJKqqtGd6VSf6G8d9zoKwFUuwg5JX2f3FGZ1C5wPtBYHAxhHrWTUBeD240e7jZe
mNPEj3Bu/pp4WHJQW+lstizJHVOKcLqayZEk/V6wKEmT6Im22Yob8B1cLIAZm3eM
l09lPK0GBHeOq0JdpPFQGOJ2N47GhhMm5l6jOThrIvc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7088)
DkHbIxAWJIjsWMfOJDFA1KGRxvl3K67ev3yLn7ocaGNudofLGxJp4FoLIEhE3uSn
qSfDPaF2OZ8npgAp6tppTRMGOqbgRgGE6b+AHHtadL9pSsxNuU4qGmuvsTZFkHKN
RSbTjQcm/3+7RORCNmCmCbCmllMJdIEM/vz0kycvJMRr8ZX4asHPNYPu5PR4pfCq
GcDW73IbBs190k0qibOYA4W3o/QuJcg+2VYvoC/Ed19zfEJtKrP432nZ+nEu4gzU
unK7tgDiXxP1QaQAWynH0Mo70urYNqODW3qp+wGqqLMLSLDIBRI+7Ji72OXyp6UJ
On3X/ZJXveOZC6xhlH0MnVWx3X9yRBgQX76stC09SlYO+ZefCwo+Lr5w6ugVpbgv
epK0jr/Wi82mNrZQmZOGaL13do8BO6FASSWB638K6CSGsbiP3OCk2bNa2gogjnoN
O7SLSULYUS7Yg/sC68qMAvu1iiULCOaQjMVQA0V6tzb/uB5B3LHJSfrf3a0egVym
D78Y1E8cfRwYUJOmbO1fGFYNxFZoP4ocuGiC3oVkYMrtswp1zHmEc8EU2TZI3O5Q
2iGvwCsLyIlUSuSbLlsnE/L5zJDZq4EaywKsRW3ELpfNu2cyx3SiZBrhsCqWXAnf
uereLpnb3xrZBSZyfW2+i+0E0qP3UmMNlsA3/DLVrdjZ6rV8IQGKJPrIJdejM0rE
7uv8a/xMBTOKGcBnHvyfjICVgfCKf3MRy0mCd9UyIcLmkTRIAXnIJbMjf14WhTyH
XP2Vhkdq6sAxWQGH3B9sPKwclSTA9JeMfscZguIfP1iuKH/OKwM3goM5vhxgdVbi
iDwcHXQw0NzbhlMUiBmk2Tl48hh1G173MghYbBDf7ck07Yt+B5CeJ4r3ypt19o0E
3eLxW/fKdAkGAxiEo3bfqtCvu5yJB8WQkk2TNlmtMwxK6r8tIwHIISjr21UYvYsJ
xsGkSwKuZ+g/ZmMsb+0jbb4wNAQcdgKEdnmXW0R8Upzqh7vFRbQHMAy8TaN1REVv
yNrIt+DY0WxjjS0bf4XvCGOtfu1i7iCep+VRTp2SdbDu2UY15IZ0yEd1uQ0ToGRv
+6lexDj54yjjGhb5X0OpnjEL2BEWMDAGvpYLkzr1K0m8DhiSfbGG+sNAdCCGG6dx
rdICE0eq2ViTIgfL2w6k5QVtNv6QR1W61S7gATUFOVLTgEDRajRHg+dLP32CiEtd
YrAnnK9A3MkIECUFCs3ErloNi8U9Lr0fvotpdFIQfEZwgNQUfh0yrQDg5PMI2RjH
ysVqV7wBCzuvhYLXUg5VNQAtokvZtZqN6g92nHwRYH0NGKvdECYUsEBa9bV9Cc4V
ZTzBTR2UhUHi1KQsx2Gd3aBSQThDIiSrKWxUAdLMawSjc/4H/FS/E/z76hiFa63l
gOF0wyEiwA02d1bXjFOzr3gCYis/b62bqqjs2xKGbZWje+pc6f2sw9DU2U+M6u3T
eKSuHF8zNRQHTlzYB360XHtU0V7zjyqZxs85t/YXy3yDpnqZHOuChpgnufe4qswe
IttJU68teC2qRMFvtBCH3Jk7R0SyGjOHWouSqISykQ9P5LW08J7FF4b+iqlLglgX
xaDrr/fPCps+KGBHCnerRZwLQnGoAlBhx96QjyCcqbBTUPEFfD0AEjVYadY7bQZY
5TWPxZrteLEfOXe+E57Bz2428liXOLo5tYe4ebVu4PscxTrqwbNOEYrUdVd7odSI
X59GbL1RyQJsNp23HYs6ozdzzfizmQWOfE9YAudOTQsTqsnRVSD8f50bnxG++PIE
WygY+VGCW6eYeMPPBfoWRqjyzt2hVqoNeuQ2IA3C6J5/pycopDAr1flqGMyPBqrd
JDipt9T7wB+OUf+RYRPoBKAvUUy9sOmmbuNp8A4QNdcF0JEDeGx1dxECY79yYXnz
tLFr9hhwP3sAb5tiuXt0DfRFvTl+CEC4WJhiU7VOCAFjoviuA+64Zu5v8PI3vppt
sfzH9AZvRQKQZeQH093qMuxNMThqPVPjVgGODezuozGJRGr7acqiRlzGQZAQZ1aM
hjivCdcwOkF73zOMcilQpZATowf0c45XE+hfhtaeTDugo+je6iSFDjx3UX1NTU6a
LK57Ze4tuTohObHwtsl+vKeWnMGztPpgHgqJ6beI2aL7jlc+imfRixF73InJ4ecK
qMI5OPYqTxkAg86nb3jbJ29T9hKo2MjKarePPKGAnGEcQwiq8dNBbSN8Moub4FIO
S4FYGnddKASM7+ECEEne3dudM5oKpMq31FdwFN5zmcdYoB8eS638BdKsa6+oBRUK
aZgWeGBHBhv3cDuhT4SK7MdQtChWBUOWZr73Xd3kQ8FHpsXGTzcktJJdHSY22h2b
yP2tSECas4mYG9ys8NZz31TqBLVZyJLciZPRrvVRKkGxjh/yXeyrVhZONeJ9Nhw9
FwTPOR7lY1Kdydf2CXm7jSr2bj4ujLtGbEeUjR7xTaWJw21SrU0m+Cj6EQHuRcac
T3mkxBXfr/CmpXDpvEYlF+ZwEOU9l3A4LDabNhItxtvZT/sUDkCbidocLgGHj+nt
wOq0/YUUJ92dIhJJb1d2SUUNlZpngp9peBvcwoCkMFfjZmO6xp+yjLEgzLDkRxLu
/uwgnjRByezkBHl5lW94nC9k7gLxyw3G2ThC9BmS3odYL0rLwEdSWF7rr6CPJXdx
dr4siaFezJR0F4VGVH80WvPr65GFi+B1PwGdxBVdOE9SoCb0fKJ5P7l+BlQrVIBJ
gdTNKTK6sFM+9ZAfIp3S3P+vM2+2QUxEr8caONZTSrm+McRrHnwESSB39p2gl4qp
dzHb0kqI1m375px9LNSVGdBAC1fo7dMXzbVE9EceXSW5Uyfmd8J2mitKFlyFVHxt
soVLLbGtk5xx8Z+keFWUwz0F4qSnckzbXcXdcHnagnmGgzzhPtGjIK55X8H4xsSU
TSTM3fQHESlBt1hi4XPPY56E3Lfh9pxpPmvMnNxbvbz6g8nwjpqjRMzSpXUoawWi
Qs0UjQzwOBOK/Fl08Y4vs/AKYvrvawEGtTp8cT1oiS9Iub1j3zH9122svqgY2D9W
8DT941lLU/T39Fu5DuNHi3uxafDBIeXhej+FPhg9IhGjqhShyaCS3aVhkRGuwlZl
oQCvLfdf7MhOKjmVr7DPXWYtr6DS49uYeMF5g8ss0FjhGRmCm926R544aa9s53kO
mh8bQp4By5LlWYmPhFYk33Zmo6rrUQ0EaZFwR5+wOwKEgp01NxcT/Thig3e2h96y
SsPR9T5IDcg5spQVeHeMf+Uhd4Mb58vQ5V2scyppA/jn9QLpGDOr+2ZpFqWvv+sZ
E1NDbymo1SIZvcXaS0xr/xrkCU3GzoLNyqvtFuFlf6F+kb4msL/9HSv0QIUAHoq+
/QLCcAXED2Yjbu5OmvfOBwxh4YVSxAkVK+3wi+uUFz9i95s9DvfMrOm4URgt+xWb
SW4ejsGrmxJoLCDaPGdwwiS6Zveo7Lw1p9p2E6bE3RCdE73hiWlFGBBgXA32d8bM
QZYQqeL5Lnt1HsoJZVA3XiQLtCxUibc69NJ1eluDtucDHBA1/qx79AKSd/7T66/u
J45ClHyla1nq4r3qzaHFFB5UzYr4s88EoXQFx4mco1Z7H2/9Is81m2suJCDZB9r4
3Yk+qfy4cwaSH8Cy8Dppv4EzGcC9SrgW2mrxzTLwO7yHrTrQ7bqM/L3mldX0wVmh
0WdGrCMzkuD7pyLzKkO4tY0ZEk4dfxtj3PNU/FP4vri+IBV0KFSI7ggVpWhdof3e
qNNYjkM2pDZ8m1biqG1YFflpWmiMNyJEVZvFmt3WDCZ9Kd5vChSQmQ1AjzSlVRhJ
8q6D+Z6HnZ82ZlrmIkwh/QmXB2PxlEYLQpcdXf/O/KBI5GjNEpnZEITZm/wpW08N
o89UKK+3cTYLVfv0hu9MFtaf5MyKWuWSmlT8txMROjJ0hCuORaW7/7ZMP3X40f2P
/MNhATQ9DXo7+wJbMiyaG4PS8Caz2Zi1afAYoMDM3K82CwuTO0tPSvfbNmlKJx+l
nWn3qA8cHgcBhFoEfxsfttHrPMtJeCdfYF/7xjpyFZ6OyN7tcSiuubrIfpnMoLRy
qfNxcxAcI7X++nNfpd5lP7/kaAK1vhslQv8egDb4Ko22qN2sZg4MDxstoV+AGcdS
gw7ulbsVWbPDk/CXhX6WVzR8Oc9ezJ54fq69jKBz+fdFgjfZfQ0lU8MDBTU4Tu3n
R7Ip+KiZ659IeTbG0eihDU2UPuNMREOE/MCnZ9p4SGwTUVkagYNKaAEHcNkPGIXR
3mgQ69PboU0fOzGTpJQ4oAiVrV+d9F67YqDrrtb9J60+a4RASXAB3UNgoiDGAWzO
qBOObQYsgfCfDIqKbcgL+1tXLBEM6GfQfTZs+4ilEbyQOeA74fPrupd7upUIFlOX
suRiC2mCN5ooIHVvQkbpbbqUhQ9PpQhmJICiqtINb4flAWjLDydxYbGMc2YxoJZl
HlbZR7UV3DiVIGqhfHlycObfzmpKoZDa/THJiRlUomVS6rlTbBTbNwcA+7NREr38
tqfl7qMfFKaUXM/jWPFsIHQy7bqfcbtxpaj5uv+Hn8S4Xyy4stLeTrH56OlMszlk
aWRygKuD8nzb3opjLLTwUZ67i5qI51VnTif4K8MSTQRtlomcFoRH6aY0vC6cCUz5
YSHWsUAUYisty+25A//ZlHfuVVWXW2mJq/1d2JYqScfEIlZcBBg2Lbx2dGQold+C
6NU8Ab5pMx+6hyDTGfBkW7BOSPz4RT5ZFtDQxc9c8Qb7e2jSMdOIHTgLJao8cBUD
C/naha1a+f1uicUc8PfVj2KaM94dV8JLDKg7glXSmuqNEMOwfKV7Mq3mjEPDq++E
FFzmreqxxYSwy8rpgzbaaeGNI3ALRJf1jERUCj/ZkoDqMzm3WRw+y4/yrmhUxosb
tF5dc3U4+UgLcQWDjhPFvO+eFJG+eQAXLmYhZ2IooF36OeMAXhMZUsULYzAGLDRd
45YKeu25emNGNqmedhQGoa1MOppSY3FoNFiMXMvydevpcAAhoC5xajoxBQfFru9g
HS+QiNGkBV1awW1brf81A8E2Fx54mTUQLr/fHGQGI7s0+UMhjB2jAvfJ8Ujhdf5G
kGj11BA4k1P6rnmfrGqL1vR0FSf3N5rKBkqVd+ebuGOvmcK9fIbKayqqj83aGF01
rWKcCvv7o1srMCKVKnCJC3FDC8z0QwPXWR8sxpvyHIGpBhTs5guGS5huYdgJ/nLA
jS/E8n9A33qWxBZHkLV29ihMihLBBtaZV0c9du/qR/2DM0Q6drTfR/LBnafVW4ZY
DH0HDvuLqI2/kQm6E2HTKLKGf5BjTtoaQgSwTyafyZ3VVFm1UPAFUTbGjk4GXlqX
+9kLRnmQfjaPCRmoA1l3nfXBaKWqjvL7XpysmN2oV4/rcDtFTQHD8FrB0gAL8pQx
6kfcqjwREplyx0koKhBtZ/4smEHHJ/9dVoiP6CdOQVa4IBZg99Oi7fCk5yWpt+61
r+qNibMt7xalJX348sVCjLypLIc7DDDssAwVg8Marl8TBvfqS9q5zz/PQLbNV9WV
KFyJp0Gs84ju3pb19FWH+59ENTWShsnOBICBk2zU1dnthUU7YkjbD+tRd0S1E0Ze
aGi0ln2zSzdozqJLovpOZdfEXgHVzGP4dtyqlAetckH/fihy/OPSDaM4hIfJMxfI
/N1UA0zXiHfVMkpWd7XE0u1i/FIuljgZlGVKURimlk1iVoGZ572mwuR2L3OWjkzp
eI/i8h38A7ufsZeWUF1qfAUDHiWOiFFFXJqkXmsakg1oIUIWn/lhW1Rfu2k/rWB+
22Fc0HLHgQ2hzG38Q2CUTiFYxZhj5z7Hw1fQS7StCFTRaRbQ+fZyBgyVg7OwWanZ
029ooLFTt4djxwbdND29sgvnSyBeCxqGtMQcA8S5DlCOzkui9Duy1YRAMhQd3BUd
vTbVBbuROmzx1RB/5/JwUKeXqeVADMEZj7lGydBbfSLSLPzMgKNv5RWdm33TSliX
K7LIB2JjrPYcHt1SYKqwlAAjVibY9MmWNhYiic517tvTvlSy15zVdQCvQhhdL4VB
9gS5paoxVi/F7IW7zf0XwSIJ8qdJ42c4pojKPrU4+kyy9BKGjeANCJRjBDDv3g1C
USsKMbRh4ZJywlsG/HDd7JAhPxhSgz3w5opNEgOkYY5AGPw1EIHHrNhkC9hC1Icn
m89mh/reQ5v1FOE5YKN9UBptDwuLmd4DmQp2pOmnckIGDzZxG6R1BwzIWzWJ/8HM
p+tcq8TUtT5X4ogZh8jmsBdNcQOaEtQIG8pAgaPbzRThHxuOg2/77zbBLU3k66Rp
1nlWgWyWNR8JyvQM14vnK2gB8OYwWQHs8/DGkJSfzMtFT8u4upfbcxhy2eys90QL
WMQIJVjO1iIVSJXde1KnlZnivtqpbv18QY3cM9Q2YQz4ejhcOeYnS1Zkyw7Sm/Yi
U8RiKsCXrltbxV3dKY4+vtQEZ/swpYvw5uY74BBtr7cSlJGkXNUsuNMiN9vuR5Py
SzKOMLSwwEXcXbecA/H//8ZF6ckF0z7oeoR4+cuE7xUS619FdRt2G3HdpoIPoC7T
nHCcLw8syypZxN5sxavfiZvlxXewK7hKnc29bYDBq8wYn6xS25E9jaU+nIWoO2PF
sCXWHUW6BqK87rhMfRG9DzbMmcU+mGM38XpT4Yl5N0X2CwATlnvTAbFK39hsDUkf
9o/VrnswKUTTTeEAsGPcQs/fIU1GUztDYTiWryr92HrfPUHgDYcHGjFj6r4PL0ug
yontTPmJVPubeu1q2xc65fJyeL9GuOyZ/XpjpZLWz0WLA9egFF5OZY7JUF7+OEJL
Qolbn8nnXmKw3KOpuDYUhf6JQzfp3Ljl+Qp2OLsAHkP8SW9wdyR7QhyHanU8PGin
5igKRBi9+HWQL9B3K9LHBcALt5jFCEpk0vvlazi9zF15WZGJEoCc3xYSOX7x2EzZ
+FzavKS3TvDLoyAkOe7P8uNpob3D1OOTTJRyn28xHA5woQ9CVaeo88YrKnT5kTUG
0bJPJ1B26qh6kvXPkNFWRY5UpIuLZV882Fm6FQ6p4PkWl51m+QVla29NPoa3wkZW
u8CXFtbKtValwKJQ8s4uJmhbpb4Q7SrkzvH5KLudRyhVZUS4aby5qrRUQjq4gm3t
yq0vh5Nr2CkQhI3t2TCCxPMnT9jbrwBSE2Xasq9m7xUVRMfTyWK/24ZX2wfvp+MH
S9lI1x64elqsAexS1NBr4e41/8CHdvpiTIkax3cHhKMbDdhFcmR0QkTYvFRsx+qD
Ws52WMukhCOkKv4jmI6EheXtzPrvhAUszzigDZkAXMfArJx1KI7oQX3pr8G6W9nO
HvueHUa2wmRetEeARF2YA6G2Bpgdp4rmIlGRckIvDOZaXNcVYLB8YLSk2n8umVxs
K8RyBCxtzad95My2NwIAtWOJpSATmLCQm/xWQTGUGjkLxTq2kote7pgDYZ4hVOjh
zy4YpnJVFDbRmXvzBXvA+VQPm0KuWLEI6vDm9kEaIvTLJxB262p8rQQqBBNShvmJ
cs507n5gqK/hlk1padXYJUb6yW7DzeKlIt0d8qa4CkK8nHuPyBLs3O8MaFoszhf0
Mlrs//MPv4MAcjUg6nUW39BobCsiXxpJrWMnfleMte0sG123FGck8IEGatbg/Krm
/1UWQQQhIvQ3yXoM2WBMfc06bBE8E2Ks62IWi0Cnz63jf1uRT4dDX6GPZ+CVf00w
7VHsdcAcKSmnVftEnZaarW/EcWx7+hcg+CWltyWMHhrRSB6BtktQ569cLkY0N2ru
0/WPlFeyhWWx3TGXbluxJo08C/qXwFsF2txm1g4ir74RN3vtU1iVjC+cUQoM/Mhw
Dfv2FyOVumzjY1/TTfLAQIqt5w+QF3BEid/KuiK3z/Qsg1MVkuRvdJQ9ELrHys36
lmZcdxq5+2whLF1ndqddyhmzqs0F0DTjpJB5hkfJOU0aSDAYAJH7PRxuueyJ6xw8
Y1vt9628t8p/+89wWmys9sRWkZFSfONXtp2SLV2PJY8hOCoVI34OO2Wv0sHjwZrr
hEh+mOfY7GQWpFQEETkAo2M9kVr+omRKVZf2FwOSKdMhi4pNqyKOoFK9E7A6r8D0
A2Hzb9ZbGeSWs990hhHuZaM6YGO7pB/Lh+SH3LnJ3WDHhWtQrK2vCweItBoG8SFT
MNVGwPWm5H4K1lFTiCQN7oTA+gDeo7OPIHgTAXxqzVAwAfHArkkjW07gw8V56U23
HHYYlmI3lVRwokrDe2zyuBX/fCehV1bEPmR0Wq02jWidrV6PV00aATaBe1ArhzLT
K9hbZYtbG0hK++8410Dd1ZQJXt4Upa2hzEX2ZgpAzHZg2tK28pRt10QEHm3zcmVk
wUW+9pxvvlsJFx2CbBMhlsDaKMz3bOfSlCg18paEm9VRQkniiG2HxuFfglcTMMW2
mnG7uUusBoP3KFon+IiwOKuEmvr6HeiN7RFvvCrEG4AOUBhl3riXZ2K1QVbsA/gU
Munj+WaME7EPwrmgn/l3z2jEBO4hAKq3LkElv0UV0WAPJLgwe+xDooQD7T0L2U2D
zJ6SwITK82Ub/ovh3DdnAybZZDAWouShFhOQlKfYN1wTHzFWHh+mORVMHrMtit1Q
P0V2i8L3sEa73PJ+0TPjQ+EReg1BndyUVFfSoaCeKpmsCloxgHbnSqiF5fvJFkAa
P3i9DqwwI6RCDXN5ZAjrXb4E0EBfoE/n292x80x/UJl+PsjdJn5X1Vowwx/7EUyz
dcQg+L2ejGy3bu6qqw6R22BZfLAxmoEn7ebxMzeH6eDGq9VmACKOgQjQjHDgTl/P
/MXIfDDe8emOV3WYrR6dbYN5E++xTKu9pROHAO7U02hO3+ZIeatcL7ld2cHzDTX4
5qTMRPj4tdP0aEFfs2NEIBOKr12xAWdNE1NHY6JAxxIfl3BMVr/uAR2EEoQTgQbr
5Oy0p5zkTx967mVDc05oQKFRQHezoep3WzpiYt7kSFCQ9M53ys4mop1pZphXdAVB
OaGKsvE03fXyvbg1DT/zFGQtrSLQgONBvQsQrzdLFdUE3rbKodjtkXgyfunlHgjH
xS8CLDtfg95apb4fhYYQHI/HWD3dhf4lTGZsfXVpCA9nC7y5sD3gNvwfhgowDBF2
k1JfW+M+/v8/3W42uX92FhHd9WZRJzawCWMSfNHQKwEqZRzPkHZ+uWg0DOqNaePu
IcPbbDrz4/JcqSCB01NS7p6S5ZSjOETy5AlCuANfs+EYo9v1T54TL/czJjPAIZ7w
i/jbqVBK4BePFhQUtL9bgAxu3V0NmfoSOwTRL41rzl4K1zQdQHYhvC0iCQl19wPS
XaZh+t4zyVxuitsOq3qTGre8N/NQ14UWxy2KIyncNSzdOlLUuc3j3ZW5hvB+P1Pt
fNVUgyf483Oq7DftJEAUmMRs6XZoTvzj7s8y4XyRAtM=
`pragma protect end_protected
