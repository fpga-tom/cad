// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
p5rrbPaA9t7jEXQ+vw/6cGwy/awwxJSjUywJ11SDWYOXZtnMU/sdWd5WEtH6G7S/
8sLetr0ytURDZfy1URl9Y28JMgoQmFBzD1fJ/LqvKHgoXB6ccqPLH/tlqCjaOppP
JX8WhFlIiPZLoyY3Oe9fZtNTnyswPE2GZ/JdFHVNNPg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12176)
Fercu2xNUlEQlHFGXJuchO4n+iRQw2Y6HPCLgLZ+FK6x9teeLCe1F6dQApGQbE0s
fUWm/018h3PB44zSUW5fGtBCtWxhhfielsy04wimFxjdw+QEnRzlhN7jlf8AN0Wl
3m9sfTT5bGGiMNSzh91GOy28PiF0otn4GbcqBirYjzRT6ieuVu8rdq3YqHpnWWqz
gCDbiRv5IXaySkTc3saF67Thkmq5Ozl+xS/IYUbURt+FnneTyTmzcSFvOimPDgHG
XWOIJjEyE5RliD/WeOdFRfzZ/2baxCfJ8LEY9jifF5dE5rRUVv98CSsZaG6+trpa
3xIHT5DwCLCzS+KCkSZ5khUfFlddvSmPKFPb/EO6GcM/X/E5vEVvC4fVLDbhFV1M
VKXqy0sSg2TtvHUBaKSq6J04ujOpTN9wvIafEwvgxlzBkoQcdi2NtVNB8BTOWXMZ
dUX+eaqyevMtQ0bJ4iC/XBztneWmPiuu41RDP1XrFCWtNVF1fE+sBE2Wh5ZCmg8T
uuVnM57x4ODCWtcvjSXFIq/KttHB7egWsqHS8gXJgVL6PWqRT5fCu13dKXMFHljz
96duMWFscGzUx+2WaFEVZJTkWYtPlukwm+PC3v7ZXyBcaiS92XFdH0fqbZ8mnBYT
O7+J6GgfoBw+FpfVyC3JhmhDC0Jop3kuG/i/RN0wlJ5fpfzqYn8rHt6IM9iJHlKR
9xQ2ykV6eLT2CJn2rIA8EeUySx0u8fZsxGercMCP1USjyIHAIEyMbr3IqsdkSp5F
vpwdD2YUZ0vDiMD8zT+E44MvAHCBGTEfWdLlfINfPLGgj7CIBku1rTrnzcOS6h/L
Wb5/Rt4BxZ4sQt2QNyeehwSRMON5efaDcNq02OXAvEfOwsCV3pDUOgf5qKDet4se
PLUoatgvmlz7LD+JfRlLPaCgWFF4oOeNckEEgHkUyCcgIeR7omLnIpKGVMeOf1EY
83YsEApoNMhJYs5G7lVi11hHU5p22+YoTMGVhDTftXdw4FwJ1fef2LRUY47ad8/S
MqwxHnl61DZ94mj+6C4DUD8cFI/sn6WbZJlH4sfmJvX43cyM9mmRCVzv2qIPZkq8
zWXzopUbfcJo51Miz1I570yBiTnQyNPE/etPDnQ3gkwjsfr/9GJMQ59YMVRIKGjm
aYtNuTc+4ZSbn8ZluxygbOgu86jKFP4NZdNkpcYzJKcVkrdPPLA13VFLuV7lFzvA
fNO10qXuRkS18venW8aPqmyqFsKlHwNqmVwwQv20psRckrWh5qVRjNdhqenF04AQ
hFq2Fty96EFHKWkM+B1WSn0EfZCqaWDxP7D6ZgIvMvYj/Bp8oDymZIMXexps55dQ
WK/TTDv0ptuv4QSWOZXm2DxwLjv0xFHKaMDeWUxBebjNBeyPUxKt00bNr1bk3H4a
KAtQa6HhrK51Nn+wpTlIZiNfjXbXNBBkm1EQ6tZmlOwC8591FzykFDceZ0qGvUaU
raSrceJIyYp6ovBlipc1h9hw7cTt4eR4bUbdwpl0JDg12gwe8sQtozw/49QFsYYG
qL5u3vjy2kBfCNrwSipM9WQQtGG7M1+DwG+lIONsCg71UNGjbGjsJH4ACc4gqf/X
PEald/GnxlIwbopEvX7NxUHVEgmjh0mTzWL96u6K8aZBHv1wGBg6hwJvNvU7n5AS
h2tRg3THYYq2diJbmRoMCv9l63Mk0/3Zlj3sP2rwvNt3nNIuo+2R2fEZpiUlnZNY
91m+meGVmOTiTe+B0L+fIxONHuyqFTQabVzMomE0Fs+dxSgaXD07jeGhV+P9OM2O
Q+zhcnVRlUotYF9s7lnlb8bJDyzQp1SHXsBEMKxKkoJFQx6gFyNPR691ld2hMASl
XJmzbO2V2cYNZBv3LW5y6maxgNxwXdodND5EtEm+rJyECTLx266u2HArCrCMLt25
WPTsSgDi8NIewq4cVOjt/WIC19aQkGAMvF0Zs37P0GI3mVeCFBzx4p/aQPbzWMQu
7vjviOZhQ1fiiUD3+dCNl6EAGf4h7k7uyIdI59Xrk7W/bKQfb6qZbIkpn5l1qaIO
xuTW5L19YAs7LH1Bdd75hxa+Rcv4heuqhznipSAE780qr6oEya6XzdQhZh3eaOne
ooy+euWMfb/7h3pFzCgE9Prbm0e/U6kClx/zv62M7d9LgLx2LQheKKNImw7NICde
O3A1d3VvG/3uCwHOfKdtmuiBaCUEgTw6cDwxsg8Hq28PAJZmiduIQhv8s/lPubdZ
nWmMntN6GSQ0HneQcRqEQ5ZxSXsZyXDDhkyYhRAorAlavUzoMQXzUGQ7lM98Tt34
kwCNSUF4pyVFM6pjI4lYiGTvvNGuI0BOctCNuEwS7PxNGOnxQR74UsT7FgDa6fI8
D13izq6+bnhlHcZa5Y6oOEkTl3vDIMvaUjNRiTRtZUKrDiuQmg8uk+8/pEQsv3bF
FtVOkwSPKBC2qpwuJDKfUe/v6LoAjfDNwJ6Xzr1g16kOTP9w2w5GsLx3BFCpQUfA
DUm4qIMQjk70fDtCT52X/9Krl2BPN1MnDQmXx+eh7VLUPFhbn3EHeZGyyV0Nmgut
z6ib6PG244VigxzCCspxUADIOwgIeypKG3H5AdmPIjnW/22fFC+SJFcIq5eQdBiN
1fWcnGfSGlHhxezn75DvVflKpVeXFmljKQvsZ2R/SgO6qdpG1kxY1vhwprahKk6Z
gnLTGo/XakrdF3aUEE/cejb33lqOb9SaDxmJXxpF/AZNmTD8jSWtY9Ntn9qS3oMH
JpdsHT3p3x/dUkmYTYeTsz37fqtNH/qv8B3Px/hSRp1UqqYmrnilfvXvHB/lY6dU
g2G0WrZh6dL6zvp8CHMytin/iuQgF1I+CpUCQB/uWZdcLdxnT92u0ia8gkWcnOnG
M4Z98iqW/P59692heM+XxqLrpzwuQnO4rhl9Rkgdu6th6qRm98alr9Tyu3KHcaEV
SFnZ548hVIMz+Gpxde0bUwnhtat9utZZdi87odska1uaUUmb6lcUCg/OZj815Mft
agrZOlxuquPiRCq4OXOm1FZMuz1xrn5KV56oLP2JsYL9K/BYWYJZAdRV1v6+tav3
n1sbDnbqLlAwNJ3CCtFpzFn2uG46Z1hxGiBNk7LATJo0kNlTlEiVxkFCIZrDptmj
YYREKtN/foErCjiFY08JHUvzew2AgNcUVmlJqQIKuGocnjKM4KUSajdbSZA9wNge
2EA/e1S62q6geZjgcN93W5pBl9S4L2zqq/N25yOQh0WLJjDOBmUvOH/n049slKcY
Oe71BNbOgVNBjACEHBnZ6tD2UCTTnewA8IZTJcWFf0odEuG4G7PAJJFhufO9Rdp1
b66pLJj5etSwpJIlKoSWhuZAuJmYek0ikBqfXb6mj54NCo+oqyu6d9WHnpmSt6gg
cJoWTXmXKzyNaaNztpalcV+28Z3ExjRgnA13NI5O8UPeZVbQddocaKHxPIlHzHkQ
hGiLX+G3vpRbizysNiUeIoKCbYCPnFnYPx3xjTpojS+aLxXYXY19t5YDhiuCL9lO
PvrECQE09Rw4BiM4ewnS6I7m0TR0EF7seh/JkXbO/G4eEPq8W4GQiDvlkEwGCeMp
IdSnvSJOYKZHwZtUufsmtmHp18PhjR3P7ivxhCcLAAqS3KG2euz0AErHPLRyPeZu
Th7Eslv1EE1gpcD3NuLc3Dq7Cf/U9SxKZGcJ2XGOxzbAalBSeD4i7CZOV0hIeVG1
A5OoCkghrmzHofhc4sNvevMze4vhu5Midw89h1kLoR/zzVbzXVk0Uz6LV/BJ3UlP
mku1ffKhBKo9weYd75lKehtchjwHhqYuE7eYmsSGURD9QFANt2ba/RVyjr4HBy60
PN4iANM1dXM0ie4nivLub+4oJvL7ZDyuJA/RCNiQKNorgHP+KWXV0NWLKVX5SYbB
KKNgJs8Icvt96/4cjXv6wOdD+e6AyipS2EDs70QUNOsL/J+kL0Vf6xJ6o1zOzppJ
4b7/XPuxEszskGeS4hNAEwnreLtTtqNUsBTpDE0zC0CqBqz1voEtji54KXWjufid
M3bVPRIwChD23zZc1cjvgowj0q9/p96vy6LbDZ/9NfzCATTmmyV1OOwliNQraoK9
Olpdf7YIHz0AOTAeWzSkbEDV5mlndcyxEvC01JbBQleXmLG925bvTnDgs3jp6Gsy
CHfYE/N7kQsi97zCteY3qnYGk2vGjTtmB+CjYc9XKJsfUVqaQT/bRjfbVSeFHZZU
SkKF4KQiDYQgTtB0jA8nrrG7DxrOq+Km4wV5xUPLz2uU9uEdEqHldvSkJmZfQ/M+
qWlCl+dszpz4Ri1QmU1h4gen5pxsaPlscJsFxFsynI0fRMEvhvH82gYHuYDOZDfL
/10MCk+2KStlsKS1JyRGJweRlg1S74aywYtd2AD5t1XMsyT5/RAlHJnOH/tzxfap
jWd1uN4FKlOXPfFXhGCfU0H1HfZ1XG6sQMeZ8wAlrXrGyOFV5PQTpHvZe147xgAB
JEAgNfgELyCMwnCHF1ecRtUS7J0FLUlka2LBy2hHW81AogJEJqgX67tgkynmKVck
YbN2SNIQPtGppVZIepnr1zdbydnwyIBQM3l0oMHHuV4OSJRBHGuziuDRagBI+t6V
PHz7Wff51r+wzyAC9sft39y1ABnwgBAQ0YF0UK5W/g6FCkoeTbeHmaxR4MnqmLe5
ar+oPuNJrMJuqVcUoFrEdE2J5Rnd0KMKA271cm4hQxTF1STGZvu97zRg0W3O6M/H
wGyDfFUHYyiDyeHg0m0ySbGaUDhJ/rBr2+JuNZ5DfYfNKQTQhmPwwKFn1BcQvYI+
P2WToQ/HoPyzF4T/9JJgizy4BwxuURMxpYCtjDG73eOTft3EKsUatM6nPvC/EvMv
n+nqNixZqbpLGIb/CWAi6mqCe5aSZyVtuB0PDf832kiKnboNkfRK3a3ze/sEn4v9
o9X+XxQT9FW8cZxc9jgX5D/5hKZXv55IB1x+fDTF/qmJ2GPjKXox0CI/fDEFd3fQ
celNgHHK5JTalRthS5ShzWsDkgUCT4moxeJiWca5Xw106Ezn4XVbestGmWRB3cQK
v9BP0nAi0WYKb94OsMxrafO72a6HrjlxW7JQLTDzYcFjaUR2am78wf/8tG1GCClI
6zaYbBp4INQSI5YwIFgkmTq15DSfzYj3hdgYOdjWsZEotTT73+P6rggmQS25hxNV
n0/j/GDw1s3/rbNsMXD/JKacdrHWZ8zmoWdH76WD+pyAFxVkcM6sOs+q8Z0c2wQc
DXAFkbZydsvZRucYXGNaEcF2POeV4uskmx3zi1Bv5bvROJf9A+qLYzo9IMC964wU
XHPZvAvzB8D8+aTHGCCgUMP3H1UXeigeN+idJU3C2YpkkwsrPL6I82tc5s6vXzlc
cin3J5l7uztAE9UF5fImxfWQEf4Q3wtv7NI4zVFVGrSnELpO36J8NHgQPltY5J4q
6yU/jPjP+wazG5dkKtuGkYJREN8IBpdrLMty3xC20hfQLW4uPza8+gv7aV20iOns
xkFP5Kn6WBIIbuwFlr4wp9ASUFzmiJSAtMOqJtfOJYDjaf9HPWniEFdE13eVHOPd
0yJvfYAu6EectH7iuSNPxtS62n6XGeed1rAzGzNH3NIe59iC6QMTV4EtrEjJi5qU
1WfHz1Qp5Ga+Mp7iXrSazz1PK4w90OAHq1s76QjMcXuWhSCBDB/evLoAcsXB30nU
Nre2qEv5Y+e+WJ7QxZcizr0ye1mo6guWiL6zF1uCj9+yMrRi2eSbIqLjvgae/h9+
Q4PeQ0iU2PK8vCK+TtGAm6++DznGxIAQm8az8Nn0m2LiC7Xzny29dgiDv/BbjKH2
Ew5eOYxm5ZYrVNhrRkbZZaHoTtWP6nkqefek84Ro/twktZYnGhf8Cw4vzSC+G7Ng
Q/ijFU4IeZNKJbW5J4N8n7hyaw8n2RElBBuvS376F0jkk1hacqKKXpHLdycqe2Ao
VIX4jWyEuBt7Wim4XjyubB+xQt2DRFfOF/DgpzKKpq4mPwTqnwKIItOBcHCPAhxY
uvbjgT5FJd2AseE4dAGOBmedv5wtlbA0j897nlJXrg9Y99hImgo4erqX35dURwwX
6jy32C/wOCtByQOvRCHcaoZ8YgYJLhbx7BQdOc8QuBPlpYdIwQgvcWpPzRdXUhnB
flV6jXVD7/xEJyFJC/zyRYq9MZaHkKo5M+TeKDJRRk4qcg6H+SfNf57/XoNu2a6t
MZFi1p6Ciket8MzXLPGMAvYRWuLCBmXSLyhqJDf2BX+21CZMPMTJzMTJ2v0GzfxZ
3LnIrdb0FG9KMTclAYVfZvofFvvkOX4ilsxP8vqY7NgJLqlFqMPRYGYeBVxuJuED
Kbh8IgqptK2bPB/NznZNQL4t9qiUprkHeutejp0cjz7/hJDQOwKn4+XlIugTdfn5
2xwGPJ7SLGciefuHEnIjt3WwNnYL+Sof6yvj7m2VVW//u1oYaKJtuChKqp02bMal
ErwVlQLxq5XbfGCfgMNhBMqc60KoCvFmUgGbIOGIK5crH4MN0QsKY75v91DA/pcC
uMBAF+QZMLuWN7fa9MErxYFcSZtGdHSzDfnIdvBbjVV2foeJuNTFicVap+wtHL7a
6voy4dQtZSfeVpCABCxTpl/TrR31MXANxq/wFfjjxLpEIPjJyGOK3BZHRvRNfDKT
xRF7H4Ac6AculOmbUqRl5UKPgIFZG/Am8GZQSRj+IeqAJdeHuEcgvB4FpdceWZOX
y5W1AjUwxXG/f+QDrdYdm7r2tsXF92mknwcOVScL4c1xuu7FDjBiWv7gZX1mPQHA
8l3yqpbX/wp5Y7SBiMlxK8SG8uGf0sGxZLAA7oQjr1J0La94XNXL4nHtfqADqBZn
4YldypJqD6/+DftvCCcXl6xtxfySsJYADfmzdLnmWiHzmdj7XCQcNAg2t37zpWBK
RdrnxKXLaX5TOERjP6yj4zj0ocGizTp4YNecVWeu3wkGAKwxMhjhOB0sqeo5W+1M
MsYCdsKlr9zaPp/jqsG7xCYpaKu13+YYSieBQqUVaHgCV3JXXykMvRcVB40ig4GY
Su41BXE4AqXH1ks7RH8Vo+BJIIR6i/cA3HQHM8ZXSce1a8JLC3FWW6p0/kZNlejB
qV1wOzbzyzpgKv8YOfrE7ucjdgf1vaDoyrmKH/7MBsZ8QmLVCIwUQQfWlY0rew1Y
JRbDbJIau3yWMchrdEmtr49Azyq4rli1LeShYVM/vKCrMRq1CyXI2Phm4o8I01rg
eKagQc4/VMjrrj0/lP6u6wyC3tQg7exIxM/449Kv8Pgi+g1X/0GeDBBxLzZWMrTV
47yMMCr4gGDqCUMsw3By2Y812yVWVZGQJ9OW9WxAMb+ViHA9Yp961paI6aSWH3HJ
zl3Um8Wmn1uOHGhTEm5Gpvq75dcwxfnV9qqJhN25CDonMY0uU+Any6uo30fT1f0j
ZCmZNRDbzi2Zqbh3LMPhmhKY9ljHZ6rCUXSKuKUtAcPW1sswqF8bOzhQYIXkOQmO
cugjsLBt9tTXrbrZhC9IxHFJqysW+nPh68wD/WOMNkLgzPLU5PLWNYDfw0OLlbEv
g2MlHApqaKPx72oNlczwF9VGc2cgLbBxqDTSTHiJrYA1SBf8YSX/Zeycduv/IzyH
Oxx7lk5z1DyrZCx3su1l/pv1Ycwu8MEAFsOYeSfajx+xu23O+0of7YVe6rzSxxIG
8w0XRvIrlnX1yUnZdxRKWCow6YehM4pl51p8wr31mYH6Y2y/nupZg/RfaffmrrAw
Z0t68zSP1U+iXHWEryeWzy0V1l7pcdQMLWPrWtef27e/MR0qR49JblKHBq28W4Fw
8s0ruU0l5TX2YDpQkVD0EmDKzcSOg+IHxoBIu7uoV6tK+u6XwzS7UiUBWn6jLAul
CWsHE3pWbDpjXQXST/BwgJXGXIaGT0Z4hUWUQ1/d53do3/vWO5BnWV+RioHZ23Ra
QSMX9ZjmQJHYhjXITthA0AeStq50/p8e5r6d783LsmVHmuVXTxoyn1eZPsksYNqO
Udh+WnTSyq9x6nWtD+UuemwZJa4w2xUlKM2saxOxUPfHIC93EQj0uUVLJfZi7p23
Ghd0ou2lXMTh60mpykRMVaJwRbJD5ELsVqKxTxP99G9x7S/pRuIjz89CLphsFrl1
+D8Aaol+yU8nJcU+tko6Y9lg4s0M59+TSnw/dhLJOSzqBj3hk6e5UFlclIynM78x
2zmOYWIvPK+YwT86MwOF9KvI5iLEDPi4qgFTahMdhFwdn8FTnkqv8dbBC57Z62iN
54km9ydQvR0smOi119anj99rB8E4kopx9KUGcz8mHxda+YS6J5FAvkHXTYL7vSdP
/Hs0xlJcipQBDZJeStv4jmwSE7OmLl1otkCNRMjxzlc0TPr8v9fTgl5f/np6fhA6
xV+yCcB/SyPfREaIhDWwWAr7RAHbpMby2KI/5ipRvdc3luP3gMm+cajAsfGweWLL
+A0RbKPxI8XG4nT0BAlYgCL1vAPJKScZvqMujV33qOqDyac8H6z9xROPY/ZPG6zx
+2HA8mTi7/ByXUxsBotdtQC/m4+e4oOSo9LQdTAwBYpQN53KBrlS91qFsW6xLn28
Vtbg8yJ99+Yy2nDz2fwnvdReEi4qHMPgxRCaLGgEqqZXdrly8C8weocq7H0DvfT6
DhOrsF4Hd+Kh2uOPoPjDcmqq7U4U2s7MF+/NR2KHeS7N5lebL2ojiB07//sUsWNX
LspV4HPc3IPp1g7WF3myE5X7DUnz1wpJ/QGNLUgy3C2nzNvQhRPAI65cFTeO37Vy
h4ilklX858EUaX1tTP5Ntd9kzzG3L6kJbnS3p08zqzDdA5hxcz9osAntZpc1IF1N
rzEcEKd/e0OIGQusq0Ek4ulFAxCdQQ2JE9UES7F7NUyKJMJNeZHshQtSi/F/0s1M
q0Cx9/W3l8pR/uqu9pbSA7VEoSuniia3VDa8Fx4hzh25NbuLVthjlE3c/l7s66kX
wi7/KHyC0Ov8soPGTxdnqXCuK1nM8LLcaVahfLvmFHqfcCbPsahXhE7FqEt6AmcH
NQyiNzPKnnfWN9Pm2vKEaYclbJA9pKeuMUibkUdvWPyL4XVOn90eZLrjJT2O2ZRL
sj+T92Yj7TdEvee7yLyd2l3hkOoSJ/s9FUX7siQ2MbVKWErvxJCLgZICCtg+543x
qMVW3pHn0P4yrRX1mVTL3q1zASwNp+F57PrhQfaFmFOX5otbEWRV3OywwGfDoEjz
kon6SWwUcQywxSLbAxIyksUuLRdwhg2jZMjmyhL42q1bH/4jQnquMI3lwovWsaBq
oU9S8lZom+YQ41I0gjF/jNoJbMfASxQ+MTN4kvdBtwcLAHgePQJGP72KEh9t493+
mCJuvf3HObdx0rXu9x8epkyVjTV0oONtstPClKUt+OqMnJBZKn2cv/5OLCLEs5x/
bbQvNaESd8lkjGHEc7hqd4rMDjBP37arNLOJUwmjfKMdRgJ4VzF5uh0lGxxi99Rm
4hZC3Ewb3tPwIeQYzSoz3MFSaKVqFN7NE2JDA4+j5pNcMCXvzZaMyo2UcsM3YPuI
8RIKB0spgYxlfUnMQ7Z/qTbf9oj5zlM53IVRbxkN1MAqlWpuIvnTuKPUfwkFeTg3
eK65vOng9rnoSWX0LDWQRmHm8gpxAS0qCovB2GGdUeYNRt09jFRIP4OnIE10P6KH
ZZYIl/zdMDzg6JKd4aOOjecPqsRxAj550G3b6bjNRrcHhhDrY1A/+KGD93VOhk2w
NGvkibGNcPNdPI9j02rlNIk9o9gYSotquYHCex14O9zSxFOyMdRRzKIp2XeXahzV
Q4EdX9QqviJLdu/yuE+8PWqEFrGV1Xy9hMxxPpr3iyQi7pPvvg0HsjOVmvQnm1HP
B+jR+DTI1g2Pk+4nuzOTPYnaUJMd64vIPuF+wTG0jbS3Pp6e04v3T0PIKjFLe90N
jRIq+Fs5TQB2XZuWd/dFUpO4yEO5e07uRIZHmAJBFxZfAo/1sNGePtu+mORHW9YD
v1/V5RBpWhhkNo2dTPez/Cx/VniS1+8q1Ud2ifwq9UOV1FGt3WE2o7ZzBL+/jaaM
1PRWk2EvhccQz+g+/A3TrERKauvF3lrtt25gSNCMByZnTWc/bCQPSSvTmn14jhLl
yMzx+OJEEQmMqs9kyZS/WCLCscH3fmV9SH/R14ex0/NnFV7DoVw7QNXB8YIJYEtS
OQBXBONpRs/nnhhiYfpdfA6VsALSJtc13PeZ3Mfwpe+W+c92ELnhtYzipuv+HiZ2
zE3YN3ZdK0n4qeWTY66uNFBvLdLuk6RZ+DVH2ZyF7w35CErJWPEhp7P+ae1pnHfB
boXuotvpfuf2+uUHnVYSRx4paNyxy0c33KW/V1rEedVLlHZhysbXmW+24fR6922i
QbwpIxO2aXtINuH47NUOUlZhQpdZ8/9qNGJafvo5T53YnZTEb7eiO43tEzzLQNlT
0uxW+9gvCac+yyLYTQuAMFUHdtZrZLUSHgkYn3GkFsTFAETIjJgE1Fdl/cvRJKZD
DH629za0YmhLxR8sg9wOlGkBpbSOrHq9od5er1UYA0Bq455O30CkmrrrhsFfdTAX
ddll5XTQcqDW1uNuCXzycgjbtTvaCLYRSSczDucOj0OlYAKfij6R24n1hp6UlxZj
WH5BCci3BI9bFTrCAH8q9+5Dfv1lSzgzPqI4resBSRJXYym3lAure3oDSAiIxY1d
JoHMmcg4DHAzD/E3VPTdcTvjv53d0VAXSlZGFa6wLUMgmVfGE+UbB9mlyP7ZEgrf
lHBlq66jQjH4LT5SOO83ADsr0kezeecTCH1Io7CAOKKQtnSaK2NPpQDKoPEJvxbY
JVMA5vonLSUlYKXbzExHVW8+ndiZEckmlzPVZQGWv0eoYlYtPM/B1b6cN9olYnnK
cP9aVQa2yE0HnuVF4jDKJh1pKUGvwKQHFkRKhSaUWaue7MM3ikEicGYNmy6t+J56
a7Vj7p4a/4vSAXp9CD5jpX8ix03X69gIjhCGOMfLVFKA0+2gsFBwupSekUV4XPQv
4MqVo1jez9jUWGlEb5MDM+2yt7UxneYVWA7qrK14dqD2sGxU+V1BksbyjOTqRYwX
pSOgKfmCYIf95DkZtzYlccOL27seeC8I9ywCB523he7I8aW0LErdH5/lV9F3PDeu
OVVNTsgOEeM2MLGWll7ir9Nz7n1GqcCXG1zfAnGLJCDYI1P/2ISufZqu24//h82N
J+IbJBthhdrG0ReB1+XEYjdsP+DSCOOkl+Lt2GrqQKPOpsu7QXv6aMAMrFSzhHJh
Xdg0Iy2SQ3aGf4oWMEsKa+BTy8UNrx0ZzngFz/07DY2tmElkiHroCaGot6xXPUYU
7GG4L4gN0CiyQ2HNedabLvaeGtE3oT2qYTWmNUco63gtN6rG5TMoQ3WTH2ccKG+s
qNog3CItGCAHjXbOuw02NZ76PVoB1rXEYHTq8bky1TzJlHVBf+9wfXmcF3WcfKSA
WWcHC2eFtIHcfGyGEb74pSlbsOcPKGylTTBd77PfILy2MosfXrBQJtU2c1/uXd3U
KGiSFWRbYTf/2kkJH0ee8zkycUFdk4I4k98FIO6+iowk158G/X5HvgETTL4Roh2r
kc1rZegr+JwcXPpEkZqn5vkjdDkBolxRaQAoZ8R8+1gmQeQwxeT4yCfN6UaTuFcf
mVIpeb5E9L86HbXhwD12/tWYzitXly24TrHZxX12ZkzsEdNdhM54eiqnYyIQ1Vl0
yIr7My2GJkAA7bGM+BQJRFXaG6d9UNqqMUYn/9l540Lw2GhgT6yY7IuYm0m+83ML
PJJNok3P8HZJU5V2KKqwvh+tk0ZrhXk7ShVCnrGkHK0yUyB9OG1jykGwD3ofPlQY
Y11LUI2/7E1HScaBf3swVp4UxXKqnsnJa3t3kClSL8FLHInKPDqr99sp83zfKBBX
ySZfIOZKccCTfAxPc/nGJa7Vlfv+7lT2/o2UDIJBY0YMJNvMotTY4UR8KOxsN8Es
wcb+F+/j5s7Puwq9JstifnTxDNPHzbYhWiPnG0jLPK6r1hw9sF7wOeWTI6MGhDPq
8ZTBc9BKVEy3paDrO4nzJ+tOuTcILi+tG0gvLfOsZP9qNY6C6oLvNPyT7csoO1HW
zh+Mc/q6sKg5ZrPhjeiD3Pz0SDHX87gFYHYMvTrbwa3q+LvpLtk9+HPUtWRo1G76
J1NUXXIgHUoF3hlDqHEfgVEy2F9iTvB8YnQsOhUDteyTTuyt9Gxb5tyJ4AMBrlNi
ORwcGGiDlehEr0JPOm6Gyvrsg5FcuoucM+0KigmDS2pUiyUowjW+KB1vnyHfB9SR
BMfrmeieBSTXLCzJhz+quiU9mGWa7t2Xaha4VsERvW6qoXevAcD2gnQ8usqhI0XF
K0qDCHTuCrL+O9deBmDdq5UBl893bMcItbJueCVfhCarOqsYJOpWM0fqfbVi4xnl
suqobwJHdnLZXpzuQBtk9MrOuJVPHAR2/zg8sefmyOU1EC+B4By7enZmmLXcSxtR
OrIO4NzB6xQnLDmeIyjDBuNF9Ex1x1flEAMJUMaWehLdvWwiHEVOHrj0KdFcYbTv
Yp+A7D7OEEOnBscY4fkUSI+3IQidKPD15UJpmacU1qgaSmZmxaJAdnF4Cpv3LtHL
w2zecZtMe+gHiUtpZ2kIH6MUc6Xvw5vjLH8aGPpvelNsRtsiXcr//h9xTeuAiEmg
WLKkmmQsPkscJtWDg6rIEs+smYBtGTEJUTdxKJLX2UY9bMl2ckEKzi2H79zzZqOe
GMSwhrR/sK4XIBNziiHrA1TsmoyPYBNeanmPyCrN5JzIMo5cs7kDmrthJjPJOtPz
a0zSs9qYRfb+3ulYiNeukdYGPOb1p2UiAeXCSb71USfLMlGkQcnwDT2oMhSgQfD2
1HRCoWBpr6zPAKDc5BYsDAKOnXH3cVuyNbprhQKNrK1Tusefeb81uI+Wx9Uv6edO
iQ01vwxGQ0SFitdE0Cgqzp0bEAc0qK4bFblxS87Y55SbJBHWdge8OU8ntHNlSlKH
/Q4Fa9C5iWtswWRDg3zKDAGGaUq8Xsn9xAlWBj9UTlsSnvrbIvMi0ONF5SZWj46L
mENToTjO68dJCPfcICp/Qs0BRi+X5waWeF9S/uNVK8qVw8ISKEo5TJkgTGOKGnZU
WmD+uX5vLKJOpbrt58CHL20enpilqObu6Q4nZr0llR2wncZj8ra4ljfdrkvhgwe8
9GTMtaiFilOaKz/kRRabu4uj3GQxXY8QXDl3eEEkwIGN/0diV4NttxZ68QVpFdps
WIJ6MlO7ZVyb77aG0XKicJaqC0sEU8fGT/bPAlMszIkpaxVNcdUo+8RsO5oUjAdD
nDG33+f6OkwwBeTHolj1JZ4wXOQQTAak69nv4zi3i56CpGqTwBnXoSDwsxHlHs/G
6PjfuDBoMk3+qP6mCWNFAoxAXPP2kwzArbOUng1a/RcubIgQ6Omc58aR1v+nvoxs
ibCHLQLkQR+xWmsk1w6NE1zaweuNxSClqrDsnqQ0ouAEYZpHDiLQZyWvOs0atT1f
bWGrH6a1EGSUfZs1m586+5Fz9qiVEhXIyYTv7g324HfHExSRjoVbK0szrxbLAALC
OWg9tuzLWdzQGij9HNoHEtBnoTtFK+LMEomcsld+V9GvzulelO4pdA7W/WOgxJ+h
wFeMTzNUtNo37HFyrSWZqRJItJbjozAuXgSxOOFz/brZIWLXgCGDxN4Ndf5L56GM
tRH3wXS+dpTWL38kpyar40+vGt9FEJsPKF5CKZma/jk13EB/qzBRmV3ee29m4B73
lVmGtdidGPl6+JB8ZJl6g3HubADVE5TL4PNPkUcsYqtr7huKdEZavYHW8hg88EB3
s+LTm2iIeZ1X31v+qRz3Fg11Rve6ys0/6bg/vtVFbkKbYQpuq9rCF3jQxpv3EQtA
H8ZqGSw7m4z2UtiSCUnZPLBkwDGQ6lVOPXMNzegZTUiMtxTpgbKeSnajPKjygpp+
PqCQo4Ni0KAxQeHsJn397qFrktTPTErTd9FnwgBdk4fqw41hQZa9bskrxvvW7SGp
0anlJ2u/5VRMGHY7e0oHPZPGsDua+GC2WRZQspPgj7d/YzOj4gRBxww61ePNIO83
mYyGKF7owD+9AnPgivvzuNJ4bO0QkXYaEuhaGx35sFMt6aqJIuzRS9dPcDEsho9C
vEu8KU2tvwYeblBRkdOLO1BehpVF34rx8GMxaLqU/4HggIaGgjGCdGOrkQerfztS
dJZb0gRuYnuGZya4LFY2N13mj7mwN1rzgdXYP3KP6y/IYjm1u3vJAAczxciZhCMw
/3KX6UuozHWRmsuzLQ8y7ly2oRtWIOsb/3KZbXz0KgoRyJeTRamiXmBE8GU9WVcQ
Bgjyx1Oxyk/gDxxco+5CPRPBf3pUK+3SgDgtGDN8AqBAa6MBUssixFI5UoTMD4OJ
G0CLxUpsi8MOG/1ib04cSd7mqh/rMUei9y6DnQ/N83A0Z58e2ixocOcTAi3dSB9i
F7gR7OuzhGKQ3RHXLsDZkq8TlIphoCLpfI0mCYlBPbiHUp5QFaE6SwsR50fRJhp8
fpE8FNgFvWcVMewj/MDzOVRmuk59Sq/a62s/5xSYzHKTOa0ihE/1doAC1x8XjA2D
KZbdopAlx9kwWLjxT3WFolgP468rkrltmgNTGyRVj1IaAOpUGLWgYkwqiTNCP19T
5/t6YM4PtOGWLdlgqD8VUiA0PZv1bYaYr5cxQWrchgqS88MahLpgtZkkN62qrSNC
xH34HgKfhaIFZaTvjSFJCEY5P1xHRHDK9t7dwmUtNZcD/eiVlZBpFvnvx5O4Egmc
RdrpsGckQmf9bXoTviD34XRirXzPiklIzOxJ7Ir0VsYkRTvOJCnlB01UvgLV9kPQ
r3W8E1uspCBf6SxN1zHvBzeLdPi9P37ue/Bzibta/fdFe4vX8u2oP1kzMvfVGNOc
gTb09UL5Kcq12FpmjJo4vBjfGe4r4+SQxhO9Df+x30bfYOZ0ngLvEHwxk/yLK24z
/sV9zsDs0W0PbBdSzLKmO4yF8Bjcdjfs6cSHogMSp9w8idWq/qk66HMntYWJEaGo
+XxkHBTbG5JefUIAoupVV8owLHEVlMV/vz7qP9U2I7S0/zbroLphBJh/Uyj46QtS
LWUng/PEE3F9p0dlsyCL8SkanuNxLauRYotz7stahSN2nZXYi1HOniJeEp7pNxkI
gfMsOzQwRoY6JYyMxUacjOvg0FNmi21Ex2pVt7JdTLp+8DXs0aVTt6nkJaHFKpdy
bDawcGGmq1z7tsCyv+ylukORO/i4j6+MCjZBdnKOGZ6NFHUskyb7/TXXzrvVI98u
QIZ9jj4fhhRi4fS8xe3jYrJ4CRVChgaME1aCs0f9wpG4WrDoXVfJdfp9gd4hT9EE
DAcN4yVLkRk5pczzL6gAv04A3O7PmFeoCR76ZrJWFUj22bWFSFSyAW6+UgishU2t
HhsqZJZqNNlP58FKVDbzmTPOtolCmmDcAdF/tjxRRIwUekFDHB3oY8x/LrWqq+ml
EHPSIDOMoN3Sb4lnm1RHv4RrXgPDopXMYMDLNKdX+AAMJyRCG+zypKAsxt3Jg2j/
pPvb+B8Tx/5dErW9WLt0rGCZiEGoLZAXI52JGGkuuZ5dlk332cFTRR8+2bsYNYDd
GqS95G9BH9bwaFm6V0rMD5boviscoW3Vw2i4fMe5RNIapquEmjg+fZZCOUt49l76
4tnNCWUyp7hqoWTfIziyxJQ5kTX+CNqayIdXo7plnhMtdlM4NOSlmOo9gKCedMw9
eXELHIovoa3Y0dHJzZa6YSDZVM6yKlEqHpmjrTC7EPd3X3EF3Sy4Z7S2rfCLWx4c
otFfreEJuU0oVyYkZ69k9ixIEyuPQNsPZrqeeKDhGYSIJXfI8wN1+5pSYVentgKM
WfTJSsBo6kAMK+jljfr/GZUpKqBrwTAm4oiLKn8Kq9AdnHE2Hy65K/yoZfAS4wIB
ilgIyQLn7cc0qV7BWqQRVtz+Z3c6nUtjIhVXvgR1lBfqMsGyesMNZZdXHXM6YVgB
vfuqKShYpEfcdVr7pbqPup2e1gfzuwwlhMK09J5tv3LGW7gAqEwdHvqHbwTbgHSl
wgOSKz16uc6nm8aroKlgt11wI7ql94UIDBEc4JnVDXoH76Y/iz/UBGRRdYM1ajtE
Dli8KG+e62Ux+vMJp/6GEQSTWpyKyEadBDOBy7cXA8Mu5HIffamD0rWHWP9p8wdj
LqgJz91Y6mFc1r3z3zEpbQ/kBHMFNvx1OFKKev6HWuw=
`pragma protect end_protected
