// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bQDbRiOxBAwYkC4t+57kH1PnwyjwKRT74LS4ImEeZs2MUiL/fBOEcZ47GwyewBUC
FFxVFAjz1BaGl4q2h8urH4kRJjKmHOpZsl/2+aRC5ppJiSSSJdlrgWR+c1RyxwA0
cgSTVrE71/7pRR/rZLsDl7p42XQQ+82rcOCFiq+eqrM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 125472)
GwmzS8fsFaKZ0zoQBRgXtRTNKjGJv8oMbYR56qaQvVDXmJ95ueEOm58XvN8jdbsw
fltgU/kFg52cgDx03B6DK0z26JKJpeu4Jx2V61L9h3oP91muA0wbQgS+ttuMrEFl
gO9XU4MeJhys6vWnIFIyLYQpZYs6bbGtZ2BME7H7UHndg98YTiH55QEA3gHR9ATk
sG4Flcx5nezeEY8wbB/Vb9nZ13caWFgnZ+jPY6Fx5sSZII2KyKE8KV4FZo2NdG8V
50zO54ZDeJDFkjni28xu4DaM+Pwl1cBvMO6VKKHjVsf2UkJ0ZoYZDebjZlMjWOA9
CQnSsSNe4F5IR2QcaiBFZeBM1rohop4WILF/a6pmME+nNeJSxoPPgrnEvIor6Ha/
mO3gilz8e2E5tDGjBHwRp5WUuqanpIrj/5i/p3FFjpTSukTV+y5HNzjlPL395TdF
pV1zGeAf5ZicrHPDilpHAYnCkB+NI+aLGp3RH/XlAA4Ej7KZXFmJWgs5N2lK+M3d
psdIMxwRBWpeSBNQiAClv8+/Rso1WGzjewAzf+1FlFXpMxxEFSlLVk6tChgnqZAr
aoapsqjd014+lFjLTmqFAHFm8j/WckhU1LXayfPjTzMByYGC6gj5qIz8mUIAvmd1
4wNtMcaA21tI0nBhZJXgTVS57Dpgk8q/ReTqwGVztN84lTipK5VwbUqNCSMjIdqw
wyyvaDaOCBc6qZCE4jC85W44kN5bQ6O9Ze8zepka0InN7LwK9cRYya90Q6An8VoS
6xN+MlSTEF3MlaiMa9+roxNtIcw0h2IojrbXwn72xYdLO6y7nUMUc6ShAzYwqAI9
FHohiW/NJLzejQrC8IYMyygqne0tIzy+x6hZ0DjqCqcalIThLVT6FPSed9CzIGW/
uUN3BLQGa2UZf4a+daps8UUsHJO12eDzo4zyR59Stm4RjyqgmC3kBcLLLdBInKmW
TcWr5gA2FXYwancjJSKDDnx9lELmQQlvUxpln7otBQEr2Ez140wqyEJjKRe0Bc4w
KGel6Omc/5N9OeUD8Enj64ZyvjbQTgtjT8TIaqZ+emWGjtUbtgK/xqvvCg/op+VX
sYUhAnaGyUrZ+Za6LTxMH/WokmPqARzcEcPGdB/4x9uDKtlCcu+SRwzmG7kPloYs
imnrPsWc2s/7TjjALji5KkYR0/4mqd4Xj8/H8bD3LJsO2z70PNUlwi86HfNL8ImR
MESYiUj3eO8FYzEtpFoCjK1FwwaUVFoA96PoLU1G+FAN2obJlETbaPPbPTzHu/oL
PvuBHJFy8kD5uNBYqxxNDI2k5DPPmG/8VMAwG4rsUGYqlXggn0YhsGZK7g132+gA
eRfr7CSG61si7iDHvrTbtO93y6X2qt6eevmRG/0YfEYzL5DIATqkYblqN1NtS6r/
qj7n9GT1gdGI1jA7QPWVsyrivBePqWEKc3U5gocM92NAYMPWSAoB0P+Ml89FEj1B
mMbujHZVd843EpmoiQ4isX5eX5RCfvgx1siPr7hpkNVnZ7X57hXuaypYVaxOPQ/R
+Kq37LoFT4M7ubUD94kxHUkothqvDmUGyjujXC3lb1q22UpvRqqAdeFJaFoRNJV0
lJ2k4gsrsxwH1ih2kyNVzjhHHMf736fXjJRQoubxH0eCex7DUpp8DrhcQVlaSqCW
ajD1gGym/LLSDHk4q6diiOr0NR8qKrdjOs++iLdluz6FNAyt1lGg/M5KHLPFLdH7
CXjflQuxwMnnfUh2onl8/R3aV8Vv+aQA+iYXjMbBbsfSYRLpLGgoNDIsJ2Xp9Sb1
rR/OxA/66c0nzwJeA76jpI8S+maWWXCesOg+4gkvOr8VG7X6LD0y2yuY1N35988q
Atue68xoUWlTnM2mGldXwfIaL3ut5zvasEQI+PYmwzx68lor+oXar8pycWRU6IFM
2NHR3WyBSSbsFL33uvy3gnvvkl28G08EJR799QJx4B9XOGrXuCSHZlnrzscmyIgK
yUrRgqC0QkxiXFC64gjbUqfr7rE1OkYzhSHbilsA6FaxYww++lFbzIjnokDuJqlO
GMBYSv1UxLsulxt7GuLxPElf2H47aOJJ1320zCJgJl/FxIgt4tU1L7z0w4VMx4+a
xQuHPZ5ionueE5QTjXQZXQ6VcGs2PAtH4QAI6J4crXSHzmoMlBbF7kV0q6CLUDrv
LUWIIWq+InoPn4FyxNVX0Xhn6rijUzh5jeUte/J8PgLLyXVFs1AV21l2yy7cWiSJ
FjSqEIjhses40VyrnDF1/CTrhSvrsVI9z6BGsT4jyVTuXw65jq2qqpCm9WZ0eN0u
/txWYrcx8Lns0OEe98TJlr7yGCG1oRut1jAVI/nk6QK/9Vx1UF7hbz7CPIJbKW8+
zAwawm4w2xeJiaqkdIcwW/BlnalUvqUd5qUYFIct17jjTYLbdAIDf0zWAT66f6w6
/VKQG7VE/AyBdzv8OegHmtrSnsQ0owpaG1Q/oKqALcTuuxrZCMh05qv0EValkF67
heRuGQ1o3DYz9rf2zvVAdVAuqZAb6DOOFej926+nIy2cyyk3k55m9Ka7AxLSrCHW
083KOLpZQvtlcj2f5gaRLum6bov/p36HE4NrmgGp9kKEsjIqgVin+UFrPD0tj+xn
ktsTfOD0DWXVP3Cm6w2zFIz4hzNGqUSNtbjgOJ103JGMTcLmDx1X/Odl3KV2zeW6
/E+ezPrUQMVS3VzcQIpo2hp+Sinab0CpqQkFXq2Kr1C6tyExnknXTd9bjVcOzwA5
Jthk9pUkoZUcjv2xablIO7tZqG/G8+PKi1jVCorN/4NtyNOD4afihe7xSa4YN+Yl
ZE6cdD/yBjTlVJV3jHpC7UWSKSU3g6U/LCM8aZi3pl9rTjBt1ZTHBxgk/z1cvfDb
l/60pncONWtLuomm1aZhy7WRCpdNZoC77JscaY7sBLxuSfnM5HIYeGmtvd0uS92i
gOnW3oO5GiQGGrCD9bohXozqchuiFW5Vj25eVdGk/BilBs4qnSuDuyxYDeVqU98k
6LFXatLsvrXiNNc3lDvEayPCTkBLsar9apIcUe6LiWShn2O7cyXdbXKt0hQkEdAb
L4Ume5PwVUTJVsTeD+nPjMzGE9bUKCn4dWtiL7XUf+Qank/lJW4FJuxmpJZJ//7S
rejgAi0npH0qGKLOOXdRS1g/1Q9AiTBc/JgNqNCC4OuBaKQ7xs/BVZ9zthiFvkci
TayxO/xp84SoIsIWBYghC1sAL0BkeokYZq3rAgovtYfXXxRMpF77DDpf42aPEuFG
f6eQDwOzqkJM3hog7Bf9j30Gmd++u5xqMJVNM0hloBXsl61qLz40tmqz3zdUyyRf
qaELxz7raukbmwnlPlzMrOxWCIzjZwt60LtnB426GMMW2LSYes+yyes/JdiDj318
r6tCaRX3A4NJUmXtTUGgCKXfttB8uzv8PbdwwM2h7KYcan5taDXseziE5b3NmI3/
nkDYHnIgAHaeY2waSx2mwMwP/LKNN+98wvDjv1AeFLoIlx6zT4LrlxjrW98OYE2O
STKibsM/ulPocKFHgW9ar4+bLK0o81hPy1QIUBYKi5XLyVZmxaeEAhrETARUdBhq
DWtPQosMo6SX7ItJ8i2c92gX/Drv/K+B8qfkBe0vfGKA2ssCvugx1q4J2+MSx7t7
zE0gjCjdRfIgOkpC0eVml+NvovMdqg0/mC2Xv5mj3GE2lC2/sftVrElXdnurQXDd
3h3yQ2Q2gRcK/KZGSk6VHkk6BBDIY/T6BULB7wU1+Kcxdt0NN95O1Op9EwJoS596
+x9UI586hn1pnQRyINSaLYgPUH4L36m4P5RC5UwWn4cOKfO+qyFHqyQVhu/wL9Cp
Am+/d875grYrvu87TQZn4UbnVRHkZI15+FPOCqqtmFQpq/K/7+FXWLm0m+LJMp5W
RBgLxBhYLlLxi9YeIWEjHdFUCvVXlRI5a/qM4mh82sL7fJlp/VZISHWyWhVV5VN9
YBTGdDkR4oaqDpUYqiCr6pyQR7SvuPMet7fuv9DpkYEH8DMIHwxXeaxD51cWp+Nh
uWs4hg0JBD6yg7gphv61FPC9XTsKZIQA63G3LS7g0Kna5f1JUPv8F3scYgqc/4Bd
j/xLtsl9/H0MpM6Vh6aSo6C8CUWTFiV7xk5U8/NpMw3xS2o4n+RTHRGxf6fCLhdi
8ayGGGuSAN6NVOUthzfMVWHiXOBeRdyPWTs19BEBsQLyy5f5PoR1RrWyTwyjyq5s
wsPrkGgbBkjBn4GSNxcmQRDXfYvmqBN/DMMPKeYOqcQpf1UFwO/bLRr2b22SX8EG
mFR4mlo4ZdLfTrcagKlATeoyyfZ+D/VpeG7nexv5MOVGPkflGWFAXvXUuwD/vced
tbkYnMZOXOHUvxPEIshr2EEdWmn5YyPatl/av5VJnzNBxFH1kt+s+wsMV+GNxTJW
QFxBLteUl7DYf3YcOq9fQGhbfSso6rjY3WxFI+CvNqtCF8g1r8dpStpcfwW07n2X
vRNElKs5Iq8qcGha0/ng9ZlUOgRYKTquzGm+9yod3Xmf8oa7g7Q/7NjvY5Jy48Yr
gi5s2cCuCHV+0JCdrK47nA7bjov+peZS+3lV4y9VWrhJjRlygINRPGfInKG5WfRA
O4UaOfmOmlbzrBNBn4z0UFIRMb1JhmaOFrRMZ5n18DruGCRbp1mzD8PARDSbjMlj
/tLjemkyMSKot1iO0BcpK7EOlwUeqFX9KPmShXSg3uKatbI/jdgPpRiWImE6e1mI
27fJ3ciVyXBeZLohIBlZfPuTbi2bNkDqjAzVBy26a0tTWRXXlA2wPwyix8pkiB9z
mP2Y7/DcJ1avY43499vx31wRDN7Acq+TAaX7gbpXPB22D6Q8+vmT3LuN43A+9QWT
nkHoc+7rF3vWLtlaHZdUXTQseNFOxIl+EajbcMnENpLcXESduNtnfRYCKU+20UDY
s/mBHVs8a9Q9dLBcDOLZ1dQ/qSW2ZHcaoNg8+/KA6Bj0h1qpYAO80JhUxQ+vrrsA
Wt6Nom5zMoQgBBSSE/VjajIgfyiR+Qb/FUywjbOC1JoPNK97BJy1cn6e8tVKBJKP
CHbV0j+JVAdMf1yUqRjQwPy5vXIPckhmd8ytAAn+1eGDOTFmeI08yaJTbxsZWeFt
5IRdK0+v+6xEjlUudhfd3tYOBO0bzb4P2Nh3MbJb0bhpBi1PbvU7GI8xIpA4jE02
AdqL7Ati6+yizCAUtnGuMQjS7hg92IvMzNuZHN2OouZvC96T8F/ECmWrqRhsRATQ
XCQ31P/+uShsWlnve2mCCDAH7nBQVKbk7TMO8ElNdVpq8sS944OWH7iSGTFpaMm6
Oux9bh61eDdCIKqF7SfyfxsBZdkL6QVhULLnM9EVkVGRU5k3EBkn6tKX6YbncDPr
gcn4bwNSCsoPsxK3brkTEscDjo430DuQpuF8w7v4kr22JBNbwPnwjcXkipou/xZu
CGixUJQ+o9eM8mFUsJwqbeZQrYoFFmgATmtzDpKAU7xzvFEUeppeypJ70A8ES9Z9
2AdlIE36o576VJLAnllyoPajU1qVVt8sOen8yQnPJJX1L91ui0KOXnktjJPE6Tw3
sp3Mo8YqdwIKJ7Xe/xE1VpEVgOjb3+rhrhnVdWmfz8+0h/yAlJi7D3TrNJ6cZUWp
RmwL/7EEjIO5GerJq3iT6uODoGSIofBfIBGkzGUmDEvLxDVAbH5OKIrKimuAHb3g
JcWb6LNHFzP93kC8R3gX2IWGlJ2Fw2OD0//BSTcS8qiiowoZOTK1a4iax9S8ji8S
mSyuNIRBmQ3MR9otyLnZcCCcEeRyiI2ovsYbZqoEqIF4NAqo4Ud36aJe79JwZnMK
o/Z3gyD1ppTXERnDK36l2Qln1tHsqOR7bpGdV239iw1CsN/i3VqPL5F5SiwLMOEP
peOKAMBRQhKvdBjejtO5M9yGq9IQ1vDYMxz+svBD7F5SwgJANiVi2bw5jGCpAg3G
CJuyhjgjDb1Msx10h5x9umKg6f5dY+OLF2cUxFM+4wf15qy+ywM17HtqxVwJ4vIm
UcReO7gomBrdK1cebqirNjAOVTnm7O9CWQNflurFPmBpslk9r78JdS3paZFFYQnK
JyEo9sKXmBGAySlx7B7K3aNnysoRD+lkAzi2N/5EAsWu83sya9hxVQgCOlmNYvuu
EevtzNY1eklptHoCyleozhdJHXwRIbWgiw84RoaSVJr0rmvAdWcoD29YqjE4m6pf
2D4SseuWrE+Kw0jKTe8VO9lSl4MioeT2pW8LkHpF9KsI7kkExIaVG3Ei0hiKyuwz
fpa3PwlsKXSiK2wWpIQd8eMGza/kOIfH6wYbbeDBDVzp9qk1mh5BtPW4u9x7gV5X
LDiw+PH7+kHTCyifzBkh+tr56qpp27oQOUmqIPhcJQshCwQ7CBjgW0+n7KaNTAlf
Xny2HuLh7bGGs61dMWdOyigChnE9/Y5Sn2HqnWQRIWPzjv85aoDkvxwi7Xuzp2w1
UUzUkInZxegtrN4mjBgX+P3Rhr9DjWDy2YZqoOIsgeJdu5pc7og3dAsRM3cdoCkL
PsukkLxzgpOTX1pCfEIlCn4/ZWsKYtdVcEYhhDWizT0B4g6XevUp6AvD8qgNvea/
zeL2iqNwmUVENLn+KcyaCtpz5ak91IiD6J+TGBirrrHo0NrAnxF8LeAphNeQzxa+
+8y3aMPfW8mn6R2uyrd+Q8jjy2R5u3YdLX/aJhYe753hxVwch2b2d2kxwGBInbWA
ePkl4Abikdi+Lsqo7drSUL+oeblXh3gBvAeBnk9D3LTW6mIZ1eWJMvjFN/MvZUr2
+3BbzG1bJ9mxF2EM9l9Eccyxu+MX+bnpeLZV9/f28C3Heywp2gB5cQZmkzxCQEV6
lcuHa++q6nzsJxPt62EGJ2csfp/CdtHlzAQ3wpK+WhaUcLcHMyy00jQl2WvL24mA
3RAw/dZdiozwWs09ZSUkfoEyBAQIV7fcVo22RrjPEKEdChgxKGjc7N6N/+RF/eo/
US0mSv5c+8waBu7CklF+bVuKQy6dDyv8psUOUaHPIJ3WypUvJwmz+b0NArmcd0+d
PKfcCxXq+mdUZuFo8tC35R5Hwfge85NFtgPC3gutNzQISOjrPv0XrASF2DDyDVwO
LY1vV7PpCqK6ToxKwUIA72fPPoMwcrJD8Q66vOEz1T4KIqNRbWlMweQmM79MCzJ1
jES9NhHzhQwrvn/90wLSSTtTFhZ59vA7Q/xzI8yCK+huH/Qcq9K7tdmlPShitJ8q
c3Sm8bJ1tJo4UM4/8yZIQSRf1wGDhUgKuDj+DFZ/HBCvYJrbOdsbIwTjnxjcxR8t
xA2nQIwCIzm43sR/Rhbmv4pe4ChoddfoNUy3Jg9QVx0G42c5bFrkdQZZUlVX2pyo
hqp4twGWXduSDibhNYuMFd1hoh4Yi7VWL0QGkfh3bF6bUbwASPDPqTCUJbg9p7Mg
XO34rJbAfbFAjkNRnRCwHz2xoidtSjfbEcajFTyehFXALdgbhFcaBpBeRsgo23VX
D+w1iM47g6JX/tps22GfSPJ8n8D9/im8g7cQZLMPuuKAX4P33/isdrQIUmDUV1zT
eWrszaNWvij/EE6PVOaCW3m0Zd0NOxGZ3Xv4j/kldcJcR4PsgvgrRB7ejRp0YN9s
9Mw0OsxVAiu0IjocrAm1UC46QdwMGO/kwiPk0Vex0Z8adAJG0RX2AO95avhGmOqo
EZMnthXV/ZsbilWSo0vcVlCesJmND1PoonqVzn9Cdf3YisFmSFLa8oex2Yp/8M6s
3qUnAaI+E5E2gD/E15U2oCvRLnE9/nkzXSxloSFTQ53Usp6wfVhfUrXIzhWu9wPf
QQoMDKg/TPgqrGyx78Ck3ggq98ogMjlz4LuT5aw6JQ2dDWR3HqvjarV3fd0/e6tw
NeS3+6cZbAYkXFQiaR9z46sfZO9MVtVWnS/wRj4c5+DJv77FQ8z64APS9T6iebSB
0hfKpn26tOdZ6BZ+sET/lwiGU7+DWPIQm37kr3XhrqZoNewAt3vHP+YOm8/3AlAM
bvzldN8mwFdptFGy9wX63Te1N5yjYlBfgVPSKDt/4Z9fVa34JKKDf35gcQY5ZCv/
epCFzjG3mfgf9CulYl3ORl+VzptODSa74q2O74W7Aae/ZnY/MCPKCXJTCPDFMLYY
fUcrZ5FSDCBGj7/BmwUCR3bTtahOmfill7IRQ3ALkmm6hE2Iao1z8d+SPsqIaArW
1YYTb98N9R/cIs/8XxgJrpGgsm89Qyr9Ey1Z8E3bPGpt+CTN88ZNe06Q4nw9qfpI
9hO0RRE4YpWYSsJc/J7Szib4Sftb40uiBT3UUrs+tALQbg+1ioVkixUqfWb1dx/o
Lqs7mikXgfJMJM17imVWuC+XJNOL2Ass7XjK+nQ4l/HtgO8nwnn71GnKhHH7VGXb
b/cMc0ZFTds0Q5bXu3WiSOjFdiMGZg19Kn10JPCpLK5+3zygE9u1ykWycZaCKJDk
t8CGOh81Fp53Sitw3VmpzoNGW+1st0a+ZI8WqQdqdTwvLBl2gmGoc58T01Jhvltc
5tFsl6ploNaeVjgFvcfiUXpHBNB86kegZ+9EXYjnd2hDD2WXXCwfA0u9GVxj5njr
qiqLQkRqkaXASBfE0NMNchWG1XW5wYy10v1K6cStQi6Liv4CVux6SxdQyiMLtdtC
FFeBbXHOBSGLjRqHJHE08kr/nsOBEDxV+a6O0UKLTISIWar+rbCYc42EG/no3h31
oiCCbrlGe9hpSqbQLr+lTXKUciuqjBwQtSEbcwyzcfI7Se1ueJSnqvG4gM7nH+j9
LTNAOteAXz5+76NrcQVifH+LItY1/8TRzz2zTvwbpBj5VrqoRs7X82nQHWI5EB+W
L/BKqzS4ATDKCL2TVxerEzF1STSUYT7eJwbD+zP1Gr2XPPY6Zj/h9KeI3njU0w6t
lWzfMTq2r4Dq6ZAdwLX3owKs2RVyxwlL8jLf88Y37evP/NFzIojckNAtIpkT+/Ka
gHahhaH3AvRvQzq4HBdwV3L3rVXffL2f9ZfDx29UWrM6NO9mmNnh2tMPsATS419W
mQEOsNe36AkdUIwqugn64g8WnusXUg1HZqrFaqwGTMpQxkRP3GayFNrwIdTW1gD/
6JexHPTORSMM+JBD0IR+yjtguZ263AxMg+khowNaY+bc6uZUZdyrnIpTZcyuLZj5
BDmP2d2hj7SDjxgsO7YNc0PE8VNf4dBx4j/uWG6H5gde/qsJiq8MT/hECyCJ3wEs
jSrGFnFxURJHaTVb9TLLbTvAmE73BwH7yypCmNxbrW86NF3hZoExLRZeu3yszFNL
WAWZE+Yt4LGJlwrGOA4vF0AJ8/wssDXSTYE120WeHl+bApcPLPnWiQCJ3LRztSer
nI8o8IiZ59GB3bTdbOSY3kdD8lopg/iVCoKpCxjpKm4jYYYwR/l7d40zaya/Q8D8
gco0wkIW1P3NWkJbrojTLJigfESz36iPOp/FPQcqH2frZdFVHiTFc4/mrvL2s6oZ
PMeX6ZzoYquVr/jvziIzRJxN+artFVFYf65cMJA1f3g2X99c5habDQm2MfvO1oDp
ttkM7MtHUQWnvXcFvoWJoslCGzA8Hwp2SxvsraekIt3FG+F7fwrzCQNVvzNcy2YT
hCJvMq++Pvw7Qmbiv5mtPTlH6plq9KoiPZWmvYjMz+Fg5fqMZUl46bFjzjqtdyVa
/eB/ZBkbKFO4hZ/icaA3Jx0yFMNogwlmu155TzQbO0+cLixu201hVCmFuJZR2foL
hQJjNaQNZFoqwxzwt0Hgv0NyClkziaAuTmZ2EEFAMA4W0/lyUL87i7c84keVThmG
MFnlzdj0+3SDNoTVY8FUwNGqdT25I0NnvPpK3QwLTrYfL4pjFQ7ApO9TJPS8Hy1f
S5Qbjm8eQNQHD1zWU35wlBHuQ0dRbzxBSmPGm6Ll4JNwoHKinLpaYH4siSE5Xo/q
X5rhU/iTx8C3iMnSYurDBmhyAILcEO0XlvM8i4qjNMb05QqfO10TApil7IU+XjjE
SYPvLhg2ZgXr6panWSmQKbwBxHGJje/Mx993Sobg2MJ6ogvajm/kijCBPJC54kUT
MpAobijKPkdqkOhpdFyCzR8tV9fiF07IdO6sxbf7ChmkG6hcCEKcyuuyarUuwQwy
Evwvj7Ngl8k2+K79XIlWarGC0tnWLOf5VbdfCHzL3o1ERcLqmzad0W6w4SCf9r5G
s+sw57SImXoEa/Cs+YEoHzi4LwusEeUXr3qqhP+o+INKwIV8vvrs6I0lV+N2wQfu
QhoDrZMMfbUga9gQcmBdmlr9/oEwT0coL+S1f+sNcd/9MuYiyLCaRoS6XK/quHKJ
+yu6jk1ssLZL9xMPj2QcUxXXIz+XpCNHevGgdGGrZCJjahaBI0XyR/+HBy9GePJv
WCgqPh+le4orxB8TQizw49lLl8dS/o1l4hH52UeEaQuTSbOJ3hXe05KijNs4cahc
mK1vAnawLNLcI2xzKqmx9HTRskallAU1NQqv0WY4SRqwDLgMi1C4BvokAwlwnbzC
ycGluwxjB8NZwgGlR6n8VQRWi3lLwTms1c6qtM9T75iNkRtFyXg2q2Zu1Lhs7Tnx
M+dzTdUwn85Uk8rCpe3VEVevn6mvqsgz/YzACjMfiikgbe8ZJiBpHPNgbEDD5b6c
B4BgQ1pMSOfodQlXlwFhB186IaM6tT6fr90p35GnvNul1X1+7FiuLnMq9jrdgXFJ
MVGkfpUUciQX8zcKX4yNDcJ1gb/ANpCrTkY3PIlPASxZCuc8fCDHzeZj+Rpjrqca
aHJEoel+rMyAeI2F/xfqTcsMG7ty3bIZoO6cLUvKWIgH2A3u3+y96rXWFYRugzi6
80tGKWrFw+OlLA04GLzgXsuAbueAZ09adpkVeGpxMpoPzlyc3pT9Ab8OqWvMEchT
E72npXEJtxpqmPZl7/J7g154ycB+5vGZZCP2W3O6pqjr+q+JOPS91hD0HhFxhtg8
sy7kkLer0ZdJOERaMes0w7D6FEjEhGjgFzrnEpPeQIJZtq5kG+JJ7oPaQyfGz45U
Mv7LxNWRTMAjW56J4NodMDW/Kj0AXzcoQ8QyzeJxYmDofBw3iu+VhagX+kywrHQv
rBhA87tcujZubq+BOliAUTUeu0hD7jOSI6iu+jtZmcgIS2qvTtBCQJ13MUK39I7B
u++Foygl3zTwPxSUEBJw85b16qaAcQ9OS28wD8INyFWQuV555Zp8itUhZB5Frea4
WDtkwBJWcpx7AA5IwDogfX6aVAPSw4ijYx0SL4jM4GXNks0zeidN/i54x3AtbwpV
eBkHoG9TweeEZakNeKJKlfAOTbog1intKgLlOqsFadzzZnPN0zojGH0ARnBaLVXV
GnM7iwcJhvBuZ/HkS+X+Fqta1hcb3zXns0N381TqAwqri8Xa/oI9EEAuaEeiahRB
fJ3JknC15Ng/BBSIAdKTSH3yZiXkOHkK6G3OQNKr6EiDpxVSix5ZYqxXxuGnJuHd
DMM0L6xMXEq81Uz78IVWjFnYsuk8fMf3P4IDmWy5UsCytQmjGOulISAcXgkUpgQg
Mc/Qrdn8WIS2+U4hfgrasEz7GlIraEwZaNxdSli7OaumFd6em6QszTVHhDkuxRPf
X8ufaStNfTqbXowc403flE3M2bban75BqtNy9sNlOw36daWd32ap2htygbeg/9Jz
pZN2Cj4f/SwmuVGWvkdCW2z4PHHBN5KmCSMKZ8Kt+ieOB4/LwuqXSKYQ1+3PZca/
ZXCOAldB/eALfj8cid3TfTOpDvVMMKWbXWildTju3lquAgKAmQ88ikJduuwtK0X3
pFRpyUlZoA5TVL5jcXv7h12V6cFNmGiJ9Yq6zqOAa2bpSL7/uL5z8SQ4AbuUTILb
PoX8YRkl3rpKI8xnqHWG/sh8RZcMm1ONZzmjtuQg23b63FT2GBIskktUgVApagM1
hR71qoG2kdQNjW1XWZUxsMzbaD99jh2h0WCoxfCI3euE8OxrkmLmGmgzls8oqWxk
dKKQBPm9jOgAhYI1K1lBRZ6vYGyqI/sGHf5KabpPnEU4YmB7IQ8kg81cI4kdgNNr
K2KAkkSckJJBCkBn+CIMjw8n8V7QawkqEJr2Ec6JPtYF7zH5rXuZ0YNvMfXR9zn7
jL2qb+sIFRBTrPv96rE8/+tJwl+OAMk6A81f9yq+uM8ODtzZBeslCVZ03mp0dk9J
pq9u9S4VBZoZcrB4Af+1mWFMwy3bVhajI2or9tbmCycGsUIbz/nISfrN3dxZ9HdQ
sGiLjT8QcalUECwJvtPd+h1vFOcM5WaNVQhW1yF6iiq7wvxyGmRmnJzXCDTQnVdU
H7TC/1I78GyCHuCpoXG7VWldk2lBTutcMCQCtUkXkuvw6K4A8IUB8q4nDZeH2x0a
2leTW1Ybju9iV2R3gU0J3Ug9KbCsWWcm/em3gPjJ/tVoqjeFRTcVoCRUoVn3KQGa
No1WNqYoJiZMIXvSz3mDBysSIf3nfVj9tBx+353yUwTtEFX2j2/8cx4FodylTwpG
wYAuOMpY6J0YuY7qS5XS0fA6/2iLQlPmglxNcQLVR0Unq6adrP+xeDNLssvCqpK3
i9lwZJ92TQCpYi49GLGBb2TowjpoWi0cDDmt1b+PMLDM/rbQMMHZDudqsyNtJtdx
gvIeQt8TU5afpg4eTwhjdZZeC3NIHGGmxjfPlkPxiVOAGeC1KilcNHqeiiTSB1UG
2onUbLZmHe+A7S2iHebTSh/q3m+hjE1T+sX4Kzeh64bbD4RVecLHwk42iH6K15Ke
L8xB/P0y+wr3OF0CM5QoFJ20BQnTuWUuXZ/DzeH32ISTw3H/eJAzp4uHquq1Y9R1
T6AgCpPSrbIozhU7Thkt7Hoj2MYZ7S/6PvEXtx4zh24YthDEXlBMsC1+VKAJa6va
5ai4P+SoJsqw5edX8HdIPrtD3bMG9AzTTp66XpV3hEM9E+hcuRcv6LSzjeD7UUSS
cCgpekzNZjvMN8n9Lz82KiCekYr6jdEX0c0lhRg08Z6C4w7jlAShM9vfkNYgEl2P
62XhYVRJnDrzMw4roo82NhZ6g1x/wPKBzKaTwqbWikGslrax0dWLAlSQJanRJK+Z
1yzW/0VboPgmQ+YU/Y4/rtkLrxxy3Zq/n2OD3eLHbuSiDGqObhT9w+dJN2976PmX
cxEcFxpVIbw+6RlX5CHAiAyxRo1Sm2eHTlbrslyzuHJ76+tzgO9UV+StpckewC+6
i7U5yJtXTE+NS6bqbIMLW3a2FSkfoegO9MylEpC8uELfhkqcVcCiIG4n7/VuYbid
za24LFo+iJsGwIrb2eWxeEl50cJL6ekqsMXD7lQBZQfZ/tXIBnGzbr7KEKNXCNZQ
TEwlj5ZLeiwIKtXo7nS7BM0UaW0h8GofCKWItFHhyoaSjU0keJm5VNIYpRJhzK2p
WFBIH7U6goDWmOoo5syfDl9bBWssAxJ9n3NQavDP3HuAzQwek7zz972rajRwvpcd
9bRMHjo3JUuuXdPye4waiLmapuk3Q7+PAwS6KK40T8GYJVE1PL45ExD4aaJ5B38d
Rp+smPr1B4Lxq5FMrcYsVlnDdYTE4rCoEFfgiYrxO0qhaoWnNxuMK9m5ZSs8gU6T
PRClKpZTcgFhVMo14fv+cdAXNIEwzCYxuhnLNjg9vWv+ZpV7a4dhdVNyUXnaWOp4
bdCdW3/WGc7eAd0m5U30G2/7qhr9ITUyWf9ggVwQZQXkEQgLCgNvUjvLtHULU2xY
A/yHtCFzoXCjc3WZVf1OSWCguweUB4w4BbncGTgH4pvJa3XXb2afXOomZMw5h3CU
jnDB1csY/bJwVHYIuoKmrJTJJzSniAXqw9s/ZWwsAURfd4Sb8vZmeBpOpKmYYYht
QuRIpvzj16zcHEhX99OTJtAZOKQkcVYXwVWgEq4q6Z9nqSfvTM3GPcGLEXAZhC3/
Y92kjw0A7VkSBw+4n/dn96ZEFnMVllM+MW+h7stzHpVeE1g0c/4SBnBANe1zoWIi
gvgbgs/xM17dxdY1rYWKr1gFNI5sLMgobREjnuY8gt3rS7pjcYXb6U6JXVc/2QHR
MsDqJs89zPpZQS6yFliVqL7XhKcWr9e76SBlp+GEafy5Nm6CxzN9L/Fob/V/INxp
86Nn0J0IU0kONQaVkrnDXej9HLxvsyDar+zlh4Iiv2EYGWScgc3d9cGSkIB/5dtG
lS9bSt2nYjaMovEfd0xtrslHq3trlJcpmHCBRaCZYgIV+/Frt4F9wOB526NMjIkS
xgofdNStTwNyT8pgaUbHvNpP1YryKEOPze4QJDiAYFFv4sDqqk8u+jK0/+mycQBj
A/n9S9fp4yHBnE1BwnqRuqGxXb5b2J6FsUui++UTE6DHCut2b5d9AP1cCfHMcUwH
EMQKyakkdb5EAJihMoWXzUciopfyqZVRTqtI/INiwshIvcg1B9M0z6pSFe3hlqZq
n8yoe989mtgjiHvRHwZ/Yg4fngo+W7mkhjIHQOhRBUzVmdp2CdA5Y4O5Cgavfoc8
ucI5EukYBewmcymkPE+S3LIXkCyThJSaM01q4lBUZE9EBnDUPWnNPhvTYacjya8r
UqIStxSL1hLBa3BFUYqFw4l8WmqNzncZ30AfGqB8MNfcrcT7U1Zi0ULwtvjCHVW/
fVZPWSiqEPajwI6BOkDYJFL3wmWIuo/1SXlYcy7jr+JmkwuoDzW4MyScovsmoqmb
CDC6HcRhYT9sJK7gjn9eM7qYr7m5coXywAgd6GfYrLpn8YvDkoxZ6v8pPu90g/Ik
zzaOKJy+sxBVcEENkZxbEEp/y4vPLDBZaTOMAIFcbLzava8CuThQtGJ0MML2sYLm
2J5TjYIcNRzzq923XOzFIDz3htUECLHKFHCmqzXpxhGkiSzJwwIxhn7HRT31ajFR
MSSlh4wJkxfHTNe3yRFiAeiTZCHPdEE9tCCanHmK/Svy8r5LHl79ZEaRZzUK33n/
FXjKzKxRABfE7hxaHVNjmOJ59hDmBmEGoOTvD4JC0OcmPySlFMSbOoNV4qLCk6On
aUNbJk7x66LK1B2isjAOpdYbNexm7ifkWTdckhIBjQaMRtd/QJ2LiindQaO7LOr7
/P+K74Uj2n1pRWSjGdmsvlIYUB/DoJU35ULKBIjjInOxT1YAajPzVh9WgVS4gIQ1
PqHH+1mRDLRdlf2C4a7xBY67VRCoZ/V3ilJNJ+nu2MX52xMwuIE+lawnzh9ROL0j
UXGQg3zjz7Jd8/+2pa+USwwONp2wriAUrjoysaSG7nEd9nwZ8OFik0B4NQfZ3EfP
Mc4RZuxr13Sqbf7X5lqx/4Dr/hHK5NKGOoO4iCl+6oTA0axgblykMDXzZfywhzcs
h2F8wez/uhI2Gw186bjADHe2+4R9J+ox2daW2Ol40k63/nq3HoE6oByie0stT/Na
c4OqdscIfjzSmUBvXrx6BYWdz+nVmKJGgZUctHCM07qlP5TseyCzOlAQlrnrWJg4
LMABUnvi9R6N1TozM7HYl96Kv1II+VNcmK9F2yoF381apDS3vw+xd0iJF4K0pa/x
DuS9FIa9bOe3gZ90DgqQbVrSSegz4tD51gb7tvq+WvCWr9TvZRnPxTs61pW0NDWX
sP0uLx2r+lhGh0A2tv/VHNhNT9FxrSZtbIDJq1goGLTRUaTHVCIta8vRITEndNVH
QIvxkULxQUntdAWIaRr4ttupEkD+2J5rxTjbKmhVvfui8TKFFb8+M3ypuIlpdfix
VM8rB0DDMIv3PGAyiBZgdMCMja+1IsOYxL2pLGK5UCRIHEZjoQiWtuzCTWbkC1kB
CiZWSGJTutj2iI4xtedbZxbOfIo6JBBB0rkchGmxrAD3IvPpF7pmXbExJyHpy+Px
ckYTuyVRkx9UIrUyWdHg+Wc2lIKEKMFifB2iMkVX2dAtF2x1rpIzOH5cDFBm3S50
BtmuymY3eNChzQ4oBRDoeg/lEfzbazvYclUvs8DZ3wLkLzjiV0NPsIvQHnDeR3iI
QR9VkpAE3lgxTnngiMA3wsgoSgmnNAv/1uDk65vP1R2o9atYp2V0O1M+8Jydu4YK
8Q4bqjmx+V8WOhTrN/rQE9gGdwXgFuCVsj5zyg/uud3bhqKAUHgbdPwiUIOgZEKv
m8Fe9miSlvAigKpfP5HVinMQEUoLzh3URCUzHKyJ4vLYpTBneZaYfMUcpghSEPrS
29Fj9zrPR/1Skb9RBlv4pomGpv76I63mmTfHWFBkmHZOPHD4cJLVkXBIntwUKSWe
PCVhOQXGX/xs0yxYDpgx6iqjgQkdWEBvdStEkRmVLDBDQ3AZQ/2klbuc0kigabTG
XR5lyEjT+W5rDA7rbBRFMBQesRQiahwiCFdwSMPeq2X28TrCj4StbXML5kA92EbT
xGdgLUAfcCgI5v/rBZns+ZNXUo3QK0j+2Nxxe3/I6hH0andpIupTKPT8W9QRU2Xp
Db15pwHvuePzIkieT3mq1kOVOb08xxdf4oqYeX0XIJF3e/KB6XcRPdDzbUQo30z8
vdjjCj8Q4fl5y6LxK1ehiynU8MFstBfj/sFSEb1WVF3slm3we4BF3xTfgXkQYL3B
Pi7A0yrRwZxZCRh+ocwdwo9obO/dXEeO1tEovjzw2YkMOAcVRAQTmRYJ1zMKK5Gq
xuBpi6mK4okw2rzbTc3B18KSEJoI8APVHAylIu2shPs+OK73aeqzdg0Z8E80I7Jg
Zv/M12GDkXMNZhGXYiLF0b1PsQJaiQQENDqth0bs6tFfEAVNxVDYUDalFNl0BhBa
myRiHhIoeYEubzw3CLoKZ35v6nAN3swhk9KmNSlZ9m6P3mqlrU+siEuZ0QcvrYPH
gpMN2fjkEqoj3yJjAp4aAFManvyiq3z2mFevKTu70hyjSlB/xslETDYeb3RCX6ps
rxFTKyqJaFw33kFJsw217CvXkHRV6HCMm9QfZzEjXWMMDlsw+5JcS9vBVD9jioe2
AmVOWqQUimasCpHolLuy9pHY8vA1iNgGqYCzcpFeeVusOM3NlS2IIjKtVERNQG3V
bUrikwB6CwW7yys6UE+tcxUgb0Ai66Ivqfmk6vqOlFHFSNZvqCRvGLH0C+x2P9FN
ts0EeO9H6FrlI09Ep1dZZGcOoUx87SNpnFBJxNgONNxij9slsC16Wq3zo4FzJkbj
BZnKZwueWvJvc7pMTaEBelpZvTtdbt7q9WEMFykgrsRRsm4KPD8QN5618nerFQwv
VeHjECXO6QgTVpGt/YzqTnsx6lbNG5NN/qT+corkO/K7TvstCQU+sohgKFmPxz3N
MzKmY/NMYHvGw2J0SNWVnuWmLx6yqhxekJoI4sMHLkQGPjbY9QB28lG2Q/AbvPjR
xWcrL/ljJs52CXYcCqkiIU+BmKefjw7Wg0I1O+G9uZvbaJOcZJgNPx/ZXikTylzy
3Zg943wcwqik3886cKPCX7oxDhTKbgmztzXAW1gahY1Frb6ZsQfixdJKWXxwf/nH
kQDtUOABYjAmCC3vg7oPj+3GUUe6YpztyzmA6mMCxQjN7eMxE8R/+qadSUkrG+Rx
hM5blQJOaplK8+PzTn9tB3Lmx48E/uZiADM4tKm0ZVMbLZkaUTOzCcd1ZJRPyU1d
Bgj1c+Tii/Dp9b7qaXeL/x52tAUDOU0TijmjiBt8Q31YEFuFE6lQHq0GKBWtCNwV
KfCkfDpRy2o2zCF67Q7rsfxqdp5CKURdTlvnzVoIUjJO+m+Xl53Hn4on9XIiS7DA
wRj0S/5WgOJK7P1IxRNzlrW7iI1qfYz9/TzAdN7xN08dIWK5fM0nGfD6ZGIfcUlD
SzFiNTlUdClDJC4htjnGPRTv6ow2xKGSUthbtyT6f8JpxVpnrqMRU61WdndsickF
QnAKCqRRilt37RgbgCAHYo1fLMa/TBnDOCEGpz53luMlBW4CHP/xeVY9zXchEhdR
AoRICDlUM9AhtdKnXk6y48UBRgPfVk3qDqzaA5ysXp3W75KihHZOwKPLGUEnf7GR
wodkpb8+yXoxDM9zRr1100aN261HkAcHYcr64xGZy4DSYvcsWXXGspCuQmed0220
bCvtcD1TX698hDskNQP8ffwPr9y5fgkX86I2v0MLAjsnTEkEXZGTPBv0/N4qHWis
hmTXF9M3NIMWLbLKVN16DC7p/lJSLsCTkBqlI/iQVX3qt1rKE8U66hRCFx4lZj0t
0++VtAFHeEz7OM2omo2+FjZVKtV5mrAPCgtlcME2OgGMmk56twowtorPqlAijyns
mULe6K+IYa3W/G6WMa7I7EKgbEzQ/d++EQ3pRgTMN3RiiQxraWK0NsT+aBSRmKSx
ITKE17urD6jbN90Gkg9dKKCRug91xWmJppSpcjXAtMzSDKgAbNEm4uTpl7JeGukh
7UzN2NcZiaSsp0KMD+k/k7TTtGoQ92UaAMO5lvKV1aFqdCgpLAUBjdmYNcyx/g7q
i+ZyyIHp0p/y8RphAOG0KTKRToNqnWnhCztDHUW8K/YATjEcunu+uq1GT+NM8LNq
KwnJZmz3gzieYaT1buBvL7jIx987zTgaiPp8j9i0gGTCsFBjUSVeQkmAUZsntMVe
qBjSCynqcjs+Z+vv4mD/gSwpWGD+XVBM2pTHo1v5N8DPqhlXHbY/aTJfiuMBIboa
0slidCwIHQTSUtLm5BCMWSrmCN/BzcbqPH2Cr2IYVs6GgrOqijfgrh/n087sb+0i
z+MfhxVGna9mjP+h3G3cyNgruLvjxN2Ht9pM2Ooi/Mz1A46Rx1Rbm+m/8c9W3NUM
RxaCqhXY/qFy4v2nSRf0xA5xNVzCHucRjueNyrCVj/JnS20pIPdiCqpF3ULnoTkG
ugufPNfhe430fEDUdWUywNqnEurGnGgMoEWgdNHvgVZkPH4qib1OKfnf9zVEPfou
iRBL/OknBfL5xPghRl1+65tLAzO1qVAq60B+aG9X9sSzpI0DsZh7urMZlDbFktzu
OWT/HP5lLIAurzgDYHY9SlsDycmg9GbZKJRa5IjG76zjMpzxPnRD7qeQL3inoTMN
GSFj9Cm6wDC3AU9UaYbx/lPPQ3Egtx3T9JUX1vBXR0VwfiIGfpyVmMXRTC3fYg3r
T68p0w5eqHbpmVr7OSM7gX8pMckz4rRcVSXqwxFdZo1WceR+6MUJFSRu2vnXx1dc
5bPvFCQS9XC55jbGnZ0oZDZFonERsnHPrRcOvZqDvOGFU51hVsJXutRpTfJH+DSd
Ywa3XFnNN1k5ug+zl6TH4vEZk4ivQy4QiZlfhYTDa/OO++Cchn8ZOpTsS5dg5Pg0
BoNg1FFNjqT6Jz5UTDSk5mGLGlHrJEsn797YtnEHYAI0NfU6x4xwHTxgyPoRITjv
rCjJMkxuBM0jhPklhS418n8oRAHCx9bId3jkKgsPjq9tYd49cAd3JzurHL64rqdG
1CW7RnFKvcMf2zN1WnB0fUXwS0DE0r1AxC8N9x4Y8a90/boSqHFNIYw638/i6NHX
OEFAml8st9tyOvyK3iQpLcsn8A2wPw3Vlgeg1FEUmgIqS6zOcW//95NPmXiBYf8f
x9xQv+MrydCKHFrF9b1RCYHT9vtRUrir4AwOXPzi1DgqlD/s8NIBajO2o2VYraTE
Pdb2+HhNDCngMVBx+/LTIdI4ryT3nLktV4ETMiyURyRDWQuwxAM7Gxtrc5d1SkJ5
Ox0DCc9GZRyls7jRa1LmYYYgVcDczehmgB+6M96Gs2MdLV7JfPsM8en24dzCKYQT
N8/TRsqrpigZBQe3alHQ/JtSMX7jHgGIlhMj9bhk7PHytzzRObpRaFR9dhtwJAOU
ODr9O0e9KtMKtNox/zSzIbaihMrEL2+GydiZ21/mVf0X1GK2qDZMFtWyZ0T0J2vQ
shcNxcHIWuhf7CUQemp6ZlowREaQIhu18SMOkBWtT+F8zVAvzEAvvL5Lt3nK11bD
SP1ZLiPY4b4x5qYEDsTHW47I5OYL/PMYE50EKN+YQ6OG+THvKtQ0wBOLH2ccv0rT
GCKGXo0LSem68w1kVZ9xkD+UEKEGF0WWcGRT+sN0vqOcOXgpBuV/s6FU5JbGt+el
MtHGx9qcsTYhkEvBpDXJe+8tk7PjZFpEOTh13zvDgVTjvmknU+rEF3c7C+6xN5fz
1ND4ZlmO5gtg6xGA180AFc1+qGIK46JTTznZ1+uFOH9JDGRwlVpvr/mRkR+rovoD
7jwaIBX4ZM+cSLyBV3P7Uo3I2y0yS8FwwGJlQ6HuBXQiUKhFeAzB4SQx5GghtAYg
9D7mTICva+4/kH+Lqtg3hR6w1EGgRAvSmqDiEeYEq22E7P/I/1Zx6mpLgdfQo/O/
gLB0ZmHkXjgZZWxRQmTppyWpQpWD8dihEQ2W1TgHaRbnHRHRJWNEhlUlgEPdwC6/
8/pbVnuxa6P1jBvIWYRnsofBtgsfbrZghsY5PpSK47HgkcaHXsaDgu6dcujJETNy
tkeDzOEpUPVv/F5lKP5+h1vSMcKyzkwQoVEANk0qD9Ct5+ZleMvPNVxJk1bOuDYo
Ajv5eYKvFAIMaZaE7RjxI52yhJcIB4I5G3c1LJOFdC0xkiNhIyPkBG6/KDSHIwU1
7S+taUPuo02vudVO/8CY3lIg8XDiN2zxeK3AV+momIh44LQyP448TLY0slxWVzsx
+4T62/8+oxa3d3gB0eUHNkE/pe2vJnimjB9Wd7lEz70wqu5dg0u9lUrSAzvA8neJ
10CskHG3XAlCup8M3LOJhB0jE9AsvRJHVB6PtNzVasuWCCHOYoJz2Oyn71r9bwxO
DkhuWnearXgyUUqFdwJHYNiEb6h/0458s/7dM1EU8X4Hcj1lvzVBBih8tloBtIAO
BfwjBswC+AEX92cfjxtBuofJOT0Uk9jPHwvbiBdmbxiyaC2cuNKSKl8vuUeIRG+V
M4FW+XEvk68rj3VcksIadMnlvQwGnsY5HSlS90A5l4xvj8esLXG7va/uCy/KgYXR
P3Wob7DPyol6MwM6jdD2VYZUSlbsWf5JLNZJ9PE93/yliyq88FFF7T2Himvwxbcb
JYMR0CQR6WGzvs9kz60nfl7j5uCFDN+njR19dDekZQwfqmbt0uigFE3usi/qCKnI
UmE5+eBGXv1FyQBC5bbYnI8VEQIYyuIVLo73hUGn2jK6y8OC4rFZwjZY1Uey4Usi
ENR/oXH+CANUFSq4kHeV9ACxPSgJE60Nce4aWd8rWqmkvLssBQ12a7L/4mBA5YSl
CTSNgAmplcp7LI0Vwt1amljNw8rN9I02b0T9jpgzh/Hvd9lPZHnA/+fx4v5Bb9Ww
5wnoc3mLTfnacgcc1iAKgUHWXLI7+0+sLF8RdOmju9q7nu6mIF2HXuhO+UYUPbZu
Jl2VUXoBQ4bDyjWxwS2kipNF0pSOwBvHqOvOY9Wjsg9idYcFBsBUcMyRN7s8wOzi
C9sqiHi3FMcvqr85WkwtbdjuCF6zYy2iDoRoFGoPwcDt3ByyR2l1jSG/B1i90qtR
r7mIbBgC4pr7QImsYz3xIZkZeQJSzDRQMeQ2BlKJUDXs+Yi7cEOdjFeUUMzSpGSF
haY03KV+2DWN++EXy21H0qRcZeG88iT9JJtKA+EBu0CfMHeR3iJ5pSoMFi5BdGtA
kaqpYXWNKO+i0WHQFWkF2UE3+YiHBbRgxJhGCPqO2XsxH8nZT4QgyCGKu7ot698o
pKmbu8OoJOBAuevGxEhvjAOM52Tau0dDoc5IhEg615tlEeuvN0TUoZoG+3SrCyZ3
4FNMlylCq4DvE+01bpP9YuJZBBDoNajubtdRs+93DvBZaRs4hKvz5NGuBqV/yuOc
oSRjoxi/34mpA3NKgEsYzsXAjKuOt+NTKEa1gD70OD/oVK2ycHVzeApfTKSSDg5O
N1OPgBk8Hnb+WKIX6SYGXG0RR13+2+eWOAVE1vccVPjHS00Gu2C7n+cf9ps45CXE
r0TlQDxrd3oZY3LZsJiYEwUHJveXT697w0ibrmI0Ylff+4cAnhRJ9X74ygJ0xnJa
O7h/kTF/U9YTFv8eNars5GJ4KeIzUeF1RlasDbc+IW+2KBR4404O2ywZRuPg/mdf
8GnB5cZBAoeFzaMR8ZEru+UOE2nDDidojqS4Nmyq7FUiCDNjKKLy6ANpppgAw4Mi
rk7JKTDkxdQVsyKk34D2KW5PAlR3kpx5d2j6PQoXgEyJuqkfPDEOeV8Z+vqSMKIa
9VKmZoHNgTDQzG1DDhPo5h07RI34kZWZRE5qVxjKF5VWKSuGB03b2EE4DCp8EIYC
ETtS2G7LY9K56rPyEgOkj5mFNBlHHJFGmffK9O8177m61uNYQdEwjXORlj26F4qD
AtPd7rCZcF/kBuW09BWbkrQB0ghAYkPQ73RTSpQqVdaTm8b4c96qICzGlstHUm8Q
aSoBhdfwwXR24zg/0FLO1ZGkppNq54/6k0mi4xF9Odt4sr/DuNpVB9ByZhAJ4OYA
cm9QeIaOCl9yPMqZhA704MuVPyZ231Qdh8qM0LtJ6TOFXiuWYiaIE8rNWnuRmqkc
K+d8wFuBQC7cRSsB0iWFJpwWkkeDGXdTBh/YqOsB9aClsAd6Mqf8S243dVrVwKYm
ulKSuGEfXSyQrhixf/FViZ97JAioM4OhNEE6g1np+IeQmj8ziBRVWBnPygBPl7yz
Wd/G/cBeDu64LnAtFRpsbmCVjnJjhYhrT4UjjpDPLX5PsfIA16pYhEmvr/fBT0Ki
fjPrJib77J7mcQhqrgWz3NAfOu8vxZ9b7r4AhGjWa1UqKknZFfldaYNfbysX8Lua
PCjoVgwKVHZ1Np57QSAXerIa4GxV0n5HfjI4dkx6uvk15jeqtCIkbX0WaCN890Ut
IudC2YefMW5mbCSOlfIDFJWJK/73lDMQYAzkiAs1V5wkGBjeILSJOXkTa5v7dhDz
mO7z5B3FkRjGAZfeGfWFqZC7VI9dPvGo0RqfohQp8zNM4iEnHIjWT/Yj/2pwgakK
aR32e1PQte2GMoRDOjfoRmrXhS+m1RSr0g7xDQz8bOrO72NYJ2LFSlF2Ahz4zdyV
/SvxTH2lWFBXHJXdxt8LITUzCa1T9+LaA+ym/iVHAzHqPm6ct+aLAYh2Fj/G8PGX
gDwqGclL8v578Mq2Lmt+3a6ZT05D3HZz4NDGbp2A3iJo2CAz0oJ6eeaheIHsbejt
pAxVcobew1fz9NBnmYJDGP8d8Gtq442+EklMamv5xbnCNIhDALrCyGCa2iNvQ17r
z2Fx3QCiph4obNPJ6AmAYqg9QBykX4T2YZbNdbyEU+r4Fs6fPfRFzP66R8omuZC6
Qh/G6rbdLG4PfWuftmqzxB1pXa83U1JkOQwWn+0Uzop8HxGHTdx/WJrlaWUtHwA4
kN1XX3kBGL/FVeUtnEDgB3BT5N24EPRnW/wqVuqfAswojurTjqjGkn3qjw1mfztm
nYc1z4DJPxK6GdreUHQPnY0+QnjLfVIskyYqVg9tRLl+tNSWHxS/2YiTnmKiv371
hRWVT5gDzgHEtN3DRAN33p6QFodnWha8cBL1t/ibkmFD073WEC7CjcXy8oO23zmG
g3UhpL5mtRyio956xwpD8iSrsUz1i253pq8n2rhjRxoZptB7cnYhx9ElkOBvodCe
IFaXMrRrwhBvn2j/dfTrBgAuKc9yuBlFrMj7bxHyWZ6SEEV9uFqIY6hTm2tGisw8
MDXef67ClXKyj7cXhrxYmfPqjarR/6Ktp17JsLeqbPhw9N8di6O9fTzIdgYC5r7z
TEYYocCQE/yTxuiHKACSTGBfuMo85yrnhdYvVBSUN7emGf0HAzm15Jkn8+lACGw3
7peEDr5SNQ+FbDEjaYxGPKVr+HQl6LQyVuTu3Sis6GD5GL5hELIXnG/wXri6r1jZ
189+cQaHx91w9nkf8bs43oA33YQwJXqjw2jWU2uWKcMOeO19OuxvXK3q/zI9D+WL
9G8mpRitJbS0fVSuwkh2mdFOL/5M1XyL+9p9iY4XafIAKSmuUBsld9noqxRAwVfN
CXqA3qamM1woqGdXo2sY74Ii/46rwR0zKvFBS63uUcfXvOkAHssw1TXK0imeAy0F
H0H5nHyYWUY8PX2/dR5OkydmiSsqItPZ/228876cCm20WoUuUc5yPD/eP6AiE8Js
ZaIeq/xfoAEcdbnaSLgOH6egncSwKFRQep/6rpr8WVcGiLcVihIj6kmUL+vmAkAz
828iBVzg+v4+LkQiUey8p8in3WeStroiVxWJW2Z+Pm1K1xRmUiyLK/sIbkD/mjxh
/+VVNlbTyrzXmpS4G09BKUZ58lP/pB67B/3TJZW0+vIFAMwf9XlPNQfeFYrA0Hck
EYMcei5X2ADm9EAMVhBZeG39tBOh8XXGqZpvbiHaN+USuU3mmKpd9WbqJFg8edZf
TYCQnDq4Ra5b8tZjEA3px1whaPPPRKIdI/IPXjWJ0y5jegQn4mW/UTzgwagunPsU
unOYFBxb4Zp3qCzMSQkLPW3ya6RhAtt6wCrTtHsrcAkdzRbxPgiG+wvSn5mm9BKD
lyIFJ4PdK8XOsMq64tAhBFT4uRLmaSyAoyYHyuFfJJi9m1mLtjxiPOUKn8/Ro+ny
NgKVAurhwzbVU0o4ciu0s+NJXBWmTrxppk7Z0AsRuUdWjapF0SA/7KnT8qfBPy6e
N5RjWLuZiLGlE4fAv6xJPFkby9Dw+DGrf9w6gkAa/oBhg9f5VZ5V7R5rlFfSkb/k
anh7jSiclWrov1mhPU3PcxPOM0vVSFXUGs+yb+xCHpALvgGMCdameCPl47AYpi3O
4q+VGIPeBK2WXVt0xWdMd/FfJTJJcHSqZnjy9ThlJNe59cPDfoiWZOFnv0W0frNY
PdSV/ELgwtiOMFi1qVAlm4Ia4DP9u9n6AW4jAn/WnPibut1so2uHOI6tEaE0b65z
1KxeUN2uzdWgnxmPb7SXu5ElCK1XlALUtQmeZOQ3tRaD3Q6jt69m6yajXD7b7012
25GzgvcJ7aaWWCiCCXJ65qaDRwLiGpK1CFoFIo+pxN3Ffs3ITf6tve4yz/Gd360Y
JAHl8nG2h4xhfGN5LeJtCnAF4fZTP88gupLcYlrNm908KB3vrzstpfnt8NLuVE5h
RZiMfuD6ir4CGZ3S95mY0f15visPcdnTe/3M08PzJQr4CxNJm2gIQSv/F3AF8e04
ASGjta3b1YXTv/AhUCfRIpfZ0HuM+00ziyN+Dzj2X5qeWrNB5HqRpWqzu+AEhygX
Gbmqn7WbIXFJlDfJRIPDvM4sf8RGUIyIdMRLTzsPX5uwQg7R5qcYWwlIf3UhoLER
ZXLP17nGnys4/qBlKFNCuurSX96MPzYe86KBSh7zZ1jxM34Ujdoy/cHxrXbs0VRY
phPLGSN5mwYhot37xFqR6K8EoF//Wm8Lze3O2NNp3v1MNFZt0k2Y+B3nVCgjEbOv
ro5gbsiwzRByoeGN+qb6GqESqPgh6fN8cUuK9uzewEvRY8lrth9GTDKM4ORaYglH
7tXxwyeotqfj/20r1NHTAHGncQlzxfwPHQrTzsfe2DZl+etZ+/ueYGSWapXH9ad6
ypSablnLDzrkQ1Lm1qlWShFge28KZg1MJDbZSKpepxIgi0IBTWrSe1k1oIiE1DXN
B84qtxk6xoZ78A/ZrGoLsLvNH/4WtWzNiaqVsJoan3uv1axjKkNgjkIweXBFm5xV
9YOWUCi0L4E2q3t44eDQO0qOYcBIEkZsRtinJwofcGI+bcJHgicoV4gui5eJ3Rr8
y8TrV80saVH7o32lG7hQqnYAGx0KPDbKeOCINggq4YZVAxTD4Gl0GmyxfTtEeEae
0VNmAdSwXO3a2C7vmx+vxnQIBjtatyHrHqDeTfGjhRY/RvQUS8LS5TxZEFVCO8EI
uIxyJArMBm+YU1CLjOza/YKdiGFn/R+4opItCU6KWhXLRpm2fvtgjO3k68mQA7EG
D8OzsKoWoWihixjvfQoMNniiKzNmFHKCka1MbfS6Q2uU1cyPAFGkPtsWHQOAXH6Q
0pBeqKg/S1mFqGtQcGT2lf/ISadkySgtw01Vx2USA6LDxbyMtBeXTeXK30n1Z7r6
NSwiXoJ8nfuYhjPWzSVBG0FkuuxMFzPk4+e0UrNQmk/Itjs/40WD6atxV8kDGftY
vg5H4na/XV4jiO+fpyZb6YY/pAmRhhd0+ozVXXnhBKgC/cq/HxnmImvS0gpZv003
kZV4+nttlBWaJ6j8+UE192N/7sMib2oUSaI6d/fXw/A7h+ybYv+hcmQZrHzTQH6J
dvGHSWRy2W5s0JifuV6Zydl3gexuoi3tU8OYMg+JufbvweT4Mn1IoFaojvr9DLR1
R5DLlKVGGeXycdHAXCaU3aJh0n6u/j2650ZZ4S3wUzD2rUaH6Lao3/ejUxoYWSoq
B/LhWcQ8GrMZuJEPZfYSmDmhv76fyKwbSOnJsGnEaSGIDofXgdTr+zevXiPjt6gh
LjtoTzuGtrBpVtilVDfHxLPX21f48bI1xz2GMyYHd1DBZjX9OKML54F0Pj/N9Zyx
jifiOBlN8oN9OXgDE1PvHgZZ4SxK8PScUSzYI1YtiT7+G3hwdtiXv+HvonUteNXt
k9OtqUqBUSKDEc+qsMxRGoigbVtEuBYyNK446iJzFoENy3q8vTFU/MF+6TT/soxA
u8lGiAuAXmIFyi6QZRNkqfrAGgxioZq3nuOgerjbDCQOAldk8wJdCjBIoRoeYj19
nh+uksx+wzpTpRTZs+QOowzlebPD6UHgCM12Wr6LfjsqeqM4+DsifHm/YUDNN9ko
uJCc9oR1wVqfxhIWdaSniJabZoXNsC2kaeMIPhbkQ4yE431WWCBoErSzI6vIsYi3
FJkXsqAG+8Xu9u06fPLF2MLLvTeiDEundhLiwCOHm3GfCqMVaj0K0guKwt44HrIN
jNYM5CfEmlxhZWZJFHcpWWARC1wRJqMrkKd678mhcN79qJe2Oh213rwx7V5foAbj
DHxaiDAsAEiB6EDZNf7RVfLJuI6KudvJW8F3LXV2IonzVCIIW2QacsCdTKkD9P4J
O5u8td2uTODoOgvsj3ccznwqeNsK/W7U9Z+NdQMP3VOVjECHzsLwdhogRU1Loq2x
Z3FSijXwPmKO3di/ecL4brxLQmO/PbxlDPUZs09fLVL7jfX60eUGlgsuewnRpTHL
rMTjg8fygeUfGLFkwueQ+WeV4LBmI915NWGKECrnHbn8BmuoH0fh6+qDXNxhUJha
esPIsBlGdvMpAiUk2ld4D4eXS3fbVldwPEQiWd8Va2a5dhHNLJXdHGlI0zgnleFq
nRc4XcsUTO+MIvYy52WlIXgVEdPutP/OCre8o9sHyoVFbyEqiEOXy54tAjXLf/JO
2Vvj7p50DD/j/RgEdIf5RMd6WBrM/OPCSjZBM9a7PrbtzCOvdLOYAT0Fv7SPu1wz
8cjxZq6zyHWXCjL8CztqoKdUFrNmV/a8N6yWselWlS4B1u0o518dwE+CIcM/lo3k
I5A06soj6oAyD4yjj14Y8ZYzTMI66/iF6ySb5OjHTDtR3H5FEXL5D80Lzgk3Vl9t
2TP+rKhmEWiQtzM7DcuDYyLrpTsHdXCkBVZNH9G2qJBDTnL6TwVkTLGxDydT7cF3
5Rg+8BO5SDp8ZKn5uai023fNIJRQOBY0o7KXxtnsucT8/jIBiUP1hnbbGWcHH5Jx
YpnWleS+kofzlF6rG8C4Q+FQEoEf9qCLiJ7vubeIkuDE0be6FZG9ij/r6ltf7+Jm
T2qPM/tkc25OGf8CGnJP9Sbfo06vtB4NPvTH5GQSQtNlgQVtvmkXZQevHSk4hfxR
9hI8hHeoQNe2Oh9tuyQ0whXTqOcjE0mr4NbIPoJAAd6ppaCz4dAVZ06TYWNLtmTw
C1TtXmc0sjE4qEGMep61fXd7KQPI2Q3Pul6kK6FOGVre+uBQ9igNyxjj/GXjPMj4
Z+jdkUbEhTkqSg4uPZVvZjjKe5apEUcwKVje3hChh41QlyPc/v+6xjXG3bHkZ6bB
uJvtuhOw85L3GtilopUze3nnwgi4LdT8gTAzhPCR2pWLb6dP2eysppVVKvvg33il
hXlVnGThs8Rljma6HTt1AZMjljjtEbAPAos9dCbXEDVUFBGcXbtGCX6u//ruYcQT
vsUX7aPCjA/ssT4h69o0ge+NzTPUJFq4fFBs00iVVS2Xr4UyWlW4ULtwYM3ZK8iA
K1fr4wmRpapgdO2OgXy9ch2oTQGszOzBhummBgQC6OXjSLPxgVjdysQXHMj2kCXY
cC2FW3OekVUtuYRmLUaifsr+NAUzT2NgYS0vtZXi8gm5veLvsIy3g9o9PbJ+ofwE
fD4RF6mZCBadsHHksDB7iZRk8J7is3nKY/ByhA2qJEAekwRpKxJ52Pb95cKd6LPS
dVj1CxklWzvXaSBXAv0TsMxZkZHYtNzAA8vfM9dhyDQiqbVRhUb5l1NARY6jQ8vo
JRBLSL6XyLjvRZ0kMNHVAMT1Ztoxuevvm85UAMu6QDtps3NSQH2B8fbtB/noWjF/
RX/MLF/rsfo6m4KkweLKPVSDkbMwNqi+pmB1amNiBsceiBSkV3lk7VSCnh+8FkzL
120einSjL2QcnO1kzNNZpvxU7vGUO7L7FbviO4cOp7TARlGP7qeUFI9YOiyFxk2r
/SAcUFPGa+dy/tH6oNs3FzJd5VgsvxvuYK6lbCWp7E1pK1QyuiQ9psxYe2U2cqJ7
cWfEA/6uC19P7yP4+s3ptx3OzxlsGjsoxO9k8B5dEAwEX27iBaLIWmUN4l8PkgVf
y07HT6QO/YrYBCnMe1ae6S3E4qf/oM25TxjRtPjuThVsLToKEUENNA8G1l7G/qOM
xgNjOVklcnEji2WtdFCcYO+017HDcc11Cf+78E9fXm4ILefu2cdp+jNKGGGXSMm/
jGYrCOHwFFqDOkM1LI18bx9lHsaXQssyFWxKmjamGsj0sWbfL0OYUF0BqbEm62M/
29UIhvq2HcYuyiuMDHvTAgTjGAmvkZ50G9q97aWqaT17RBUbCb4GyrR9g31w/pd+
P9EeNQkFw8i5BELycFr631UqAWfSCZnHtJQuHjYHLIoJYCSQhwx/VTM0fr2dzWFi
ZnlFmxc7oxoc84LmvYqjM1/OuJLSVWYMVEF5SsuS+uIeIodyeJ/eeUjcnI7rSzMD
EQADcXCowwahSWJ/brZjYsKVEGxCqdZnx2adx0AtDOwerFHoIoCUVKH3OiKsXcTp
Do4ZkVyqXQsFoGgwjOa1cxzd7S0B2u3zApyFKaN7EUty8hYUSCvbUNj/PXWy8bKN
+zAiYQTu2pVyAkwyXB8wbah36ku5ScbtheFRZ8SQzNGW/hS9CpoyVcMk11TY6KFd
RehRNl/RjQvEW1Xcqobzibjl2fBDPqRu1TvC1u49WqTXgjKTeZOftcIGPkyZj+nN
GNGiFoP39JOc2rDc9C47TTjW/iuHw+UVYNBrlxTAQHqnbU3FrtSQ2lsrLtTp/c3B
dYY5Gxd7EntnO19i6zmOt6dYGDjkFrbqoTCwimNj4OkhLvQReqYErJ1sozIW9PhW
ZsS1NjkhS0scFfzvYGLwmLj62EZHqMlq4iha6xQSBxVTpRaUQe//8CvoxEul6RRU
qOOV7xY4FPRgWSkVQ4kBZzye0vQlrSS1eFORpI0eXVA/HVfscDsxiX3MQZePalYb
n3uH4hGrp18QXHXv+zoqMRjlhqATHqWU50Lpp/DT5HhUCinYHAbcZ4GSgaamZs1S
JtHuZs5PWaZVidZdocj2GaF9SDjlbdhSWbrI0znDDFKFg0vdk4sQJH54otDLog5j
Cg634WZ9HqjyzKxJ85p+YAmxg2eoKgx5ujBnD3ABRuH46WEnv92t/HCwBuKJe9kq
H7vKXzzC132Owwv1iAydVWxMpaToWw7lO1bu91P3swoRVW69nTLjzn4hkQQGFiMm
lplfx+yElbCs3BjbAlZzwipgM9VG08RdlaiE/WZUeVUYcXZeaAqTimWIQi8O+Hp7
sZMY5rbp7O4flVuEKrl736eV7mxq3pQcbZHDtxZ65La5uADbbTZXjB3eySzhldrr
9FjHrz8NBYXTAI0GQDgBfmSRIhXUKCeiNoH3L/3RBhwSjLWE7qmBOSToikGtxGJu
r3klj1IeNKsy5wRISCoryLQlaSgB5rpOdvaowllabuHO+SHXy8/y1eFz8sugOCMW
ugEtwvkdXKCcKxbubUdQ1u4l2NNA9rmkpMGKOskUbPgaUHvK+5WfFuBTSTtShen7
rOkE0S/u/ef/FWKjJb11TvsekggqteJF99Qwlbyi/HPMcOyJUpUOA1Vydismpro4
cTNybhvRrcJZ1SRDFNhaejAsu8mt2nrLRRGeOmqZrmFyX2TgXwYFhn1XhYuRrrjM
QD8W5SBYeR8/d0/K7EH+KbgiwXMxV6hAieY8bBqxJC5jd3equEVnWAz9YYByoz7N
pc3xwCM2qlZosqx/YeWt4M6P3/HcSDUmuw7eCOXIYv2OtDPIHfIk3Gw11m4M3Wg3
7prfgF/soMjr+GuZTRosGpysgSqWcjDvnRFkecQsDSPvXNqTy2v6OwwDWagjCeXA
xY1w14jm8ssg8wmqgTZGrhrxX7pRgws911fkHTw0Lq3dIo4hn0+ofBYM/H03gSIA
XL9VYSd75hrOtK2zvhNOqo3+paRj/w9AFl+exQeds6zqk8h3x1CrJTqqFonyfO27
28AwcwOLa5NvfiYLfrYaFXkW8Z0wsQ3lTaRuQjAhdjbPHrEMl4oiQTn8hDKOHeKx
teTTz80mDFNV5X+KJd3c/wFI/yjpknryNYc0gR0p8hu5GtTYwkVnhoRzwPuQ1kC4
ctQ6gLKbxcCEINXTiC5AUU2eKKd+AJOr0QyisXZlbKvd7g8cA76hBpt2iA11OXu4
s/FCtAXAq05PVM1NbTyfHy/qvJ0DWRyntUA/KjsV97jNgH/Ej9ssmKyiFPa0DJ//
MYhLHBLdjRiOOmkkrm8S71X8GtjZZfjYwRxvznKkhkeTx0GfioC1PDWLaQmkwySs
ecwAYTLoR2izPo9GnZbBskh06M6JRBxfjsYTb3qvS2L81hZFpMSDdtsv8WYeON2h
YIZZr5KFdYtivp42tlXI6jo6gMlsTde5kvMxKxuMlolKosM8PoISEukMcTYYG42u
VSGxGi0/nC9mr70o7rwn7hFiPQw96x2ht6YOX+9PK1wGZrapj+XOhvI72Uo1Ro5T
PN+BtzGTVhlNrhRlKpPvmvsK6zdxGrkhxGr1OWCEr4fP2KxKG+tt0wbb+hwduRk8
1L6nwcqABVDvrn5EV6iq78OoHWgdQxXQ00u7cZU6vuFUDzp7x453xNGiK9Amz6ck
QDkNaQtURXQrFl901wV6txqEK1zFUZkhALB6Y9jYu8Gq0uLhg8VOjdtjPXF/sDVr
B2rcjMIeSqf2QpMR0Fkq5XYkmM1Al8V4Lmu5llUUD28SKPQsAyPQJFe1NMrtppV+
tS8VTyu7GYPA8QKLjSFb+VQpy9N4rQqv16sM8AYFI2ZVB+Yb7jZSRgc+CJ77dz6c
KMOKhZP11KPwQ7HMApi4btPP2mjVA0tgJmiqCy5hPIIligvaBartfz850mVuvZys
xc9Y8F4yK+DsjQRqGwMz3vMCgrUYK7m517wHJAH0xpkXoUvIDFgYgsc1HQpjyKpq
Pu9TGoHelk5pPRWshndQgSH0HdtQmhXJod7EeBF15XIK8aUwQLBb85y8eHYpVG7z
FQiaFrWCp+Kh2kTv543okr8izE6+ynfQT1IH0h0gAasrTFpS53gnmX3ktnpSxesA
zqa6zGoQQNA0HQNCEpSVsPFWcFckvwo770exmwcHpTqgmOmXeWTOxJ6+K05PS5m/
i4LmuOR2GZrghfDBG2TIG2J2ScWHeOK4M7n4lMfDgVT2fkKBC9fEBuM5MXtrzuo+
xH+5b5pQa2OSjcdvMPp+SK+YIXMWM9qPoI9+FLKqyMHZypnuPpiEZTPftEnEDqTq
CeClotFBhBE5aVuF6lrEFA58pMIk340DR50mO0rVyA/lgcJQYICxcjuZ9wlpdIo+
GXxxMe+LGoUXMkiNDP7lvz4GXiSqktBRUDvvCUgi3DKrtFpsCZJ75rC3UMswvXqc
lMgk0GlTYJOPfrXDs3uE0LgZGTrMPBpbjpcdZPoinSgk8bZ3409DvHW9GA5Mv/4v
BTgwU+4kqcZJlSxEmw/9ofg79iFDwQGtYywhRJGR/Z5Cq6gA1ZR+r8BMGMuRj6LA
AME+5tR8S/bTSDE2FtoEqW8KNmywvnibq3w39YHX+n/qNS3n3sCBJTJWMp6w5T2+
eFdm+/l/O0mX90B4Q0k4YXoXPI9QvkIZgBj1ImS+b0GdR4u8QJmhAoTCoTyhenUh
tgbHbM3mngwDgN+QTFKeGau0Q5ll3CLCEpbSfOzXRzrxM7zUc+K+IWU3Ew8BgMx4
ERVSIYNQsBeqOWEU4lcq8xcW7znY1fBppH9MdQ5X6IncgZy2szUtDYROigzr6Rju
/naGIkG9EHPZf4WsbC51H1J048LY8+Ah8/aYk1G/3hdoRKPl21xiaAWLPvXaLSf3
vC/BDgJiLR/BvMf/el7gNIe3uWW6OjnJbewzkkLp7gW+z+1jcSl53gvP7kur/1Fq
KJQ2gCJWpFRCAm69/BBFyMju0jO1+DINsxqzBaV99ny6W7vfb/bcygVMUEQnxCYj
adQRn89bP4TC3meDOyS46sTrHEAcRQhK+shN/J7gVV6rdDZLEyTVXhqtUHuG9eXw
g2DHM1IuNed1z6oz7Dm2ITGpPCiMlLLnLtAS5gI3rXi45ncFb3xt2mGSLR+mii36
6N56SVBXliLUndzDYhjVS0JYM0XEGRua4jLHYK23IUZRkZphrczEct5MB6DTMLd9
6q505NANp48NN7tkk45hpXlFwBGSJRVaCsa7D/rZPD9/qEIUCJG4TCDJ8uNCjQfa
dx7QhFkbQ6FkYNg6gmk+zJNcHufmx3utvpBWkH9ZpnW1vqbcv8m8JxE481/hztXv
SbDeUkCezr0V3Xok3+E2KDYqkCA5boJz2Br+E9ZRAm4uGGRpmlozwdGtr1Bv3HCz
mp7QgVM0roZSy5iJVsaxvcbn6hL4bIXvSsG96Xmi4nwqCCmTVWsBlSl6sdnNiB9I
UA2ODrBrW1sdcq2UF4+OyCJB2tIdunDkj4gjnzhsA32sxlCRUJ4bul7E0MjOOoFz
CoBQ1qfqSDRLqqOPMzoYNwVqpK0LczvpuNcEXN4foe1k9z558EwFd+HVUAMH9t82
rGu1ig5Tg1vmgifH/UwsFdu5Sa4wje+7giOHUBRIwBYC18DbSSqa5Nv5zW3uM9EY
fGf0at437TW3AsPGKRJPQOcSeCwLhw2ZDVGd8GuNDmX33hINV49Vj2Qc+JdmH2w8
cD8g5C257KvQ2thbxnLgn/Jqdd6pPIkIZ9zVCxeKtA2PTOoXi2LKI4JyAg3/P44t
57JbJfvyoWaX2E2baxcGHj8RuynggnGGZHhUIQUXzGk/wEkpfn5wbTK06jdg7wNj
vOjPJUuI2+D1XELzdnQd4VGHgOppNW/T0dcZja1dDKx6MZw/vGEIxX7iKaLw3R8p
NmVr0rq6AtjQYQgU88Rrb6z2WQTXanLCSTs3jmkUAW7DOSHY8E0kO0LgiZLuKXcl
JYq24yj0FbdQFpIeaK+TjtxQb6eC31uCCQ29w7hsa8Ib4tJ6s7TPCf3tJf3tIx/T
qtOPVOJLJJiGgdkE3MszsYbIRBYMFH1mJWsyOasw70RasbjLcZJSE6ANDgsBMRiG
ldlRzQ70tfw+26YgevRRPQSV0KHHQgZLkQO4BKpJquL6lEgyrIOczWR3nrBm5NeN
9W3VrOTumYGWW0k1gyTjEbL2D/8z8mwB0rBfYCbfAqAAH56Vshd1BepZC2iq7dZl
ONoJC1uPVmC46uhuQX3WKZ0qNPgA0/WtURmKSb6RIs0aXX7j+n6C8rHA9vew84vo
s3Bfu8+huPCCHc5IxxTe5KQ+dizQkGnsMn7PRvwbV1WCCbCzt8S2gJKBna1Grr8Y
iPB6iY3B64RSfPS7W6XEs0RcIJoc1/hW9d7oo9asOBUwYNnr53d9/C5gLDp4eO8J
NBNMh/oqUmspTXCH9PnUmg9ffbIccEiVu3gPvPPa4IxJVBpFBd0UCqH2p0Q1g7IH
XXamQsVjhr6tbmd9VnjkQy+51+Bvl7iTRHlfrXzoxvBLWHMAbFCZ/bzVNMXrX8jI
sHtmrpN97RRLN95vEXBEFEqlRzzEQeg54z+6ezmUHup/wcOWYE/+uH04jkAKnSoU
IRa2l1VTQFrBWZ2NiMT7by1KfrZes/ewne1HetnGYp+XxBehb9VBpRVfIofQx61o
fFPNjDsHN9WZ37nSgbNIBSXpNAAyOfpUcxc8kq0UVpKBiQGdRzAH+wxJOl66hIJJ
t9U53V22Fes0dUWB40KUg76b6M2KkL0pQTWgk4ng4UKlJJgf1uZ9xAqTXvHmGmJX
9bNqzXoHc7Yuuouc7oCfLNcu3uFiSMKxI68HhTMIsx/h5Ses6beWwKMmgq5FO9MJ
NK2ZSTRDz8Sj6VjBs3oCkvUGzqFv8JNN+wLOK/6/tb90ONbH/gWggwgwikED6RHE
xrmJke5QtRXecsHZyh2OMh9nsQRGR+ehnBRc8VVHY02UJl4sgEnXk9a0Cwx0M+TM
9e7osCmJaQLuxcy6xSmU7cXqJ9z/S2O41ZngvRqSWQcylnM2E2GWsfkPqJF1qft6
0niWbXjJyoqMnn+hBuyJFioebNs95Vfk6DfsJ1glVSizEOERoXEoFuE7fOglFyJB
99PjbuIJvKImfxJUVap8PFUoNGMmefWyslWQFC0lDZrNwgQf9r4FN4SoaZ7yqIay
veRrQ7c+PWXKWa1G3f578eXsUUfSqGRuxAXFWwpIgLSScpB+2+cwLBK1oNuZd/uN
K+GjBHoI5IShDaz0tmoxMQG8db4RCNBGXqDtEFqwNz6jzKK5uXLo3nv7qB3V8DR1
Veby+MPTuVuap6A4s68A6TPsCM3ryQafNbBviQEo4d+imkqv/m5CAOjr2LR9DWl5
7CouhORojw58Tb5NdF8gB0EbblmC3l0ldWunbvGCRR5b6Ou8yARvN5pt5xQx0h3G
uoxrwlABeNHIveudf4+WhYADE5BIbtQyea1xkSeuOS/x/+tHKVqvirI9KEUNXoDX
+bVGBKQx8Xzfb8VeDUCQceRWHPaD+7PAFNUsA6qpT3e/3NY4uhH7zc7sx0S3wHxp
LhcAKM1cSZnqbVDyflbkAxwmMp4xo/1Am8XPgfVkOXcQCzOAFUqenKwqncqxanFx
WnX9KLecPsap4IDrt5Ak8Ido28ge56FdSsX68Dw5+LOXU7Te/GZm5HTVMRJjIPfo
jMD+A+3P1/u0TFyWfP+uh0JxOMUtP9nXq0qeJ/p/EXmced2QvUVGv1sVVjJMoPtZ
U+PR3yyGveT3OJ4s02ivoN3rWYngrpVOtV944pDifo5fKkxDuzFbXP793oS4nTFN
Ca7avWXmVoiWqGfumvTPTRBtG3CJXBCMcdrhtXkIe5nTSjwcf714yXZIiSVocpto
T2Bj2Y+dDLgJ6iquOK38loQlQMXNYTMKGLoC+aCCTTZ0lT5Cj6/PBiw2PZLJ04cA
XIYQ8yAJGzhL2FmyCQXkGq0wy/otmqzGyxR6TpgNANhmX5oN11SQRaGfaXCN3Omu
IEVaBEecfa92Eoy/dV9wl1EVe5GFwN+hcA5+99bJVkVNaohANO6ekA5m0GWLaW+G
3RJexrvZwf8HgWOVhknDvzo86qfM02O9biKh8fePpc9m2fhjWpupJzU641vz6vpO
SbYvPTwdDV6VfN/hC9AiRSAiSazFswRKS5Y+Vv8ArKdHnkemJ8UDEP/6CV55/1+C
tWCN9zAN4AHLsNFLjlSJ4RxBXjmgW2VGdrUfTrWbqxsKd3+z6JHhq/AiButciQor
UzU9j8cgO8HqwKkc6vTAVY3HcszaZ33c3gC8XQj+M6JdkUMwdZF6dKQE9x4wePCn
JdN6UPCJQZ1DhvhFIaCsj0PPxGbUTu67Oxkl9FeQKr8pC51SUR8HWPrFQAvIl7PI
dQTEdR1gxGXrHdchFLBeYpVAVRbtiDAQgQNUfHvdbQALh2USPSYx/VCsj0qFZ93S
k5a20sfuPYo6uzHBE6OthCr/VbHko7f7v09IeUYQH6NjxTiF2Iy0zYNnfS/6qxG4
toJBHBk3nl8TSUE2bNstStTn+nDSYn0ijZtq7kU9YWChN19zzKjP7nzBp2gDmUx8
O5XpPZw7UDMM11nr2e9X/O+vWHRUOkfQ03Lvissa1IoZ5OOpPQXoOz6TYRbtkcOV
0j1sKy6iTG1OvcYMvv9m4+jXqPM7+o9v+O8v4w6out6GGefeL5dtN7X2TUeelgkm
y/qpEz+uMJOl2eUPI6BwnCMvMLuuY8xGpsEGsgHLEUCcPbquaxfZo13UrLkmSBLx
NHeZWdj8cPW3C9cy5lhzmBYcW3J3cZCofBftDl8q1FWuBpaDTlQHE+tkhn/BBHsq
T9OzxAd6r2PHcCNOJ+zkekAhvuBPke4YrqJ2ExfimLLastBuS/aB8wwBxrCcB4Ht
ISzcBkGSDiZX9NSi3DSIj7aNxBEBaNYELjqs7XtavR3ugxz4s5bP1xXEFNwYDqaQ
CQSdq8yxyJR/5egRxwc8YiODojzfDag1V3xi9NSugZoa4UsLMnMoDfyeZEDqSt1+
PUA7CxnoiGlT/fKv3MwOYvpjEk5Ri8Jr/AsVoHlfEphJCG0xQ9xBdBYeaRfnCifB
V6Fxo6JaHv/4W23TRQw4LOXqsHnXfIyqx7xeR3h+UecjRk5wVTYzUpS5T6BW/YIc
39TFCny1xuIUKZPW+krcFXn9EaBSqmdoj2GnQ1fNWNHEqVj8xHEmWXwglGYZ9z5h
sTMu7Ffo8eDkeZDBuSerri8bJSEkBstHEjSA5qj7tLGwMl6b/hwC5jK2MHJzl/Se
1RHxFnM1lmHAlYzJuQxqhsS3lm4K1jMmi9S66VeodW+j2eQxErW6CaMO6piLJq3c
qpFXhpMFSXgR2CdYwJQJ9poo4Edy/W4cYgz4wpAXNGBIP7ehpAEFBtlimuPGfSZP
9tyVD9dIyfPhE8+qWOrYssIktrbBoKZt8FCaHMb7KE5uFt+f5KFqbHIU4h2Nyu1e
/GVsg4VrwaqpZ8ZWsQchHu9cIdjkrzlp8WMhw2O+22lUhvJ03CkM179VcXpURfOg
P7bOujjZazH4gUCOpERVr6jLmpEl1NlsKdljEyhNvqvBUnV8FhPAP/C3gHCbU1bm
6pZGfEWI3A/usCTR0dyjUijVqSWeoOigp5DPNW6jTCn2ZHLxSLCqwr68ONCF22JX
qEvDYUaXzOEG+nTsz/UV0sAJOw9d4GRv4tzOkzgJWq6p03CT3kJV5Aj3hROvrz4S
185k6wmInmcn746ShL3l7y7FyFYraGY8ByyvJhV9ohDb/uxJf7X/UK4q9NEkjYYY
F5Iz/6JKTTRDoBOReDZfWE8weKwtGV+dGJWl4Jj5uCmAojqu0H2NDXKIfyfBqXw4
h64isPgaEBb2UudQr7/oumAjV0XlU7IIM6uG+4CNVNknBsXR22CIWLLoZ1QZU+JD
ieBkRVBYISgciiaM1rW+vUq3LDyPtLAFc/dqm0el/Md5XaezngIsNjnB7lpuPRju
1eciNVTq/74/bt9PeZwwVuMPwUmNnNUJDq9lBX3dmQACF8BrfK7v+p4oDwidfXel
cCRdPgcNMwSgrrwbuisX5On/3Kg2w0Ily29XmVdoL8rJcOK4J1CT3j/gYwbFiIyc
7i72UZ9M10NIac1LTKrBkzovs5SRFosqBWkFAUBBTH0BrFP914X4TYWx1/aN5g45
OsoYZYKrOrnsm83EqtewTD6HZEI6Qg9Y1z1wK4EMxRXFLcukZ5QYJXT3OMJPaoUn
gNmgOMXzJNlkjkpWjZITr66BizkIHRYomBN5lve/YNgz2KlflOqzoiFRcM5wsnMy
/zpcDo5D4FmFZfMIMtYXshYxLZ8t91gePVSQ9LCVO1RQeYPQNuqs3T/1jqDoh7Lg
c9xxjWtMGwVMHv+8mw1bYX5YxWJOExOSxDWxEaFHUj/wKdZa8FnjyCDyirBkbtUy
Rpd6/tnHFXXVxcmZGqoknZ5WcNjVpmeoAbaoQ6+pVPFVROWNrccbUEA/tcu+t01j
7KO8FsL3cApNzXCBZHwF+dq3zeVx2Oc/tb3vcw1BuJXFAkwS4EJGuKY5Jc35bK6i
WBwCWQtm3iBXuBzc6kqULrg/0OJYmkOFwLgyVpKr0NkcvpGXrIR9Gipa1xZ6/RsS
lq6MWxa4yxYn+zjpsH5d+HEdOHcEfeXnaSvpbgGh5fnlgqPeQP6OExhgI1MrIQHw
oLqJ7sZOOtbZQ1lcGlg7aVLCXP3P3YY1sXKPBqdQOdIIefgcjCcW2u9zHUSAxLxS
r136JNWBuc3eRXsRo062+hzN4MbDiJv7MmHaEIY4boOp5JEY27ECPqC/goKoMAER
81B+0gpbTjfPgzM9il6N1oFMnwH+woDlmzsHVJFPAXngEeA4QOwkqhnzU5ftsdwM
0Gl1r3BXyHldzMPCY2ctscTLMWdllhapMBKgtl/pWet9PbQdFtqniKxzHLW5CrG+
RNNoXvpsH8Tm58a1gg8KuMyteg+T8oxgewj812JTegwJz60sch5vS18BJ0Vf6DdM
MXYMO9tGC8vk2GetOKpTaBQBdBN1eCF3WYd5E6sTwxGPy7Sx263FQvFLBgIJ2XNR
VajymxAty+RpWxdW3IlqIUS7N27z7H5DRgA1zgrtoDiCQZsgyTALpr0FOBVvX4gT
EwAXMXS14OEPcYWsUaPpJSrFcxx1NrWlcsxSTffmkEO77XynEqhu1dK5Kt7A0Pgz
VwxU9amdScGMnbu/3rxpNwSGuDXNOKyT0d1mDtxvOdMAnOYyoQFwXJQrkyk4Rpnc
XT/8xdMY/T1Vu7nihcfQPyfi1QaV3lWMF23v7JiDiGqFx5ozSBRqIKBE+eba4Ywk
vWabWjlj+l8Bzt8iEStYdpP2TECvq3FAYKGrq/TnUTaxJGffOzcgPQnzBMK5JG7U
zBif+PCewJMZGocPk67ZGZ6Ik7qbPVE0vLsswl9gTPeFEv3PJLGcXDkoDG1OsHi1
fpd/zAAluJiKwMHyhHGu4aiF/OYCkazG8Ybsq2Csf2MXd/45JbkkOFNWFZqT0TzT
5ksRQk2DJ6OZE0G03cXfv0fMmJyMCPzuo1Ojgv8KIXWmup9lcxaIPtiwWbiF4sxY
JoUqw4I6XVjK+Rqf/tVourFb17x8cj6mxjVFJbDFrp9EcuY1v0MnETrapse9Xbpv
cNcFKGB/gipTTTGJlIpDeLu60o8Qd+H5l0eIGDW9twPh29IHuvEA/vKBtE4S9l1f
n13I8RNDG1koHG1vB6S41rxwdVfJyMb9WJmqMyA4TmTVD0SOYM/HWwBILV47tFpw
Y3hmSHeFy5002lZaJDmqBUKF+3j+I48zD+44pqz6VdaZIqlSR22nbTlU2gPEeK1c
MVqW3ei2i+xqFs/kdklEKZHqigIwq3dsfKGky9lWKvQWLCh4h0Z6c/82qoMqdOj7
414aTyLa3voXCTDmf2ha4k2fVxwUSmLIhxZKEJYTYOnApcZzvKoKQ6aZ1Hp+ySzv
WoUB0dR+RMmmidMlK1BT2+9dE+07ZdZrj7mQWqqU43j+MB6SLh0MlTWwwbXulYs/
c8cO/d8txU1WcfzIw9iCczoCWYnE6wHHjgTqdlW7EdpmB8ywHEG0HI5TylsSo/PN
2gdlIssk0DSc0a0GnHziPI1Gql+6rMjcnwK8S5oua/c5nOnI66b3SCqVWHxqplVp
NJBMQnVZXPiRiyujSQecYtVNSERx4VSF97zpf2s1KyRP6YOKhRp/gZwTEeX1Umsc
jbhZaUkIsQ/yhBVP8DBify4LsVCCxgQuaYhF7nxOfkiTtKl6NBQHBVTTIyLg3uFt
7iHtIA2gtFhqsHJJB04u+/S94G97feqIZC9TRyP4ru3Qj/grt1RwIp4Ehf+8hAM4
4nPxWS3kDTvyQshz53pqyuxeYtdrNkft+tYj4Wwjr4HbQlYmz2fuH80iVfA0Evgs
+9KoCQVB/Y/Vd/ptu1Pj1o9mLJRmmv65msTuO/wlE1DvdaTLWVPoPM3RoyuLzE23
4ywnavJ8m7SzwPsTUwoI1fxvEGTsqrXCKQGyrv/AX1aUlLRWawoqkZYl6gA8gGYq
uUEjug3ZIswJOsOsbqlan2qbyawk4UeIMfpwY3yhEtw/p+8qwve3+OQyFJzzftYj
FwifK0JZntL4gYIkQ3NkJq8Sbj4IzZ+kQpv3neeBxd3s5neIgxpC6BxVbHZwKsY+
qX6J6DwEEQJAgYHXJLypbrCvs//otZ1EbgDi6tkl3CTuodziPcAZg6BheBh3mj6M
ALBnRHWUDW4Y3zAXMLSHGnqU2CDdTTqGoKF1CXW0dsiLh80ePuvKa25faPRMQeFX
b3fXkU239vZv16LCUT8t8vW1s9GgcnxIYQwiT/eu3WrWhzTP23vkntGfsjTkXciN
8nS9TiOBTRqJ4W+EH1oI44BUBuql8oxODpDT/OoyaJ9XmfLAYNAPyNXIQEQhg8oP
S9NQdEne+M5X/SC/2wuHREnZ+axI3pJQZls+75WPW8grANsjmrSsyYE/5Tkwdfww
ZAF2OgteStya7J9EEe3EhPA4vrgQ7syVLZyTlkSE74qE94huTS5XXQQNdz7w/uN+
VLEBR6BQqqxZIOSjARAGdxWhdnyZS3lAiFe55UymP8/laJ6RTL0QzlnIGUNMdWna
DrqDIwmruv6Evf4xwozoY8avmeB8jYwxfvKlOLTtajeBE9+VK89hOr6ZEvamRcje
R1eqGGec0pS5ELHb/grDz7OJpoZJKvO9E6MDQMqT673gCMzkOo5OhfxciuuCJSN4
DGDGDfdhMiYX6Mz/aA+GC/Ij85J1NH5eyyjlqPnkfxXA1C5fuQ4+EKMfY36L3SVV
GsBVqBPAxYdbxbd6npK+Y84MUSJyjWK3w79oIJ7Ms/PJZbUNXFRQmTFThzaVRnBF
M2FtM1r6ufZzIdKu7byuGwaaFf/dARfkYYJXOV7nqPmdCOl5qlyIQNHD9OaAS4CH
cc3BL4zctabihNZQjHip0M6yZFxLyEMawpnOVdwUsFV0W46y2zf5KnClqDwmHQmJ
f8D3NAUyWj1PudkpT1nXCZ1Cbgzc6YmoJ0nvjZJqfHOGDVNNSkk2wfFQPpugdtEP
iYABK3wXjIc4R8Hd0rqDL6UU+vaeQjGMExfBX4AN+4YNSQeZmAUJKjPqo7CeHYcI
iyMtwWHXOu7Sd4RqtSt/vuuRhvkRNotyitmuVxyTrH1cKRrL4xXGZ6ocghFic8Nq
7i/XWGcEppn/3DNMJaWuxB7bTboHI3Kqmscd8QXJXDgkZuV5ELnkHyy7IOrhMuMf
C31VML+fWU0I4MBHmpmTbF9ahJ5HzWNlFwAD/R4NexbPtWIzyT9xW158zlK77N17
bF50XT3UdbnwEQjeo9fKQAcB/Qrt/zTN6sWGyIVQOR5NCTspMmeDvh7rs7ifDm8w
LCqETMab9msaZb6IjcsmcXzIoJTMMN0/2dJhKKNsjkD55s5HltBVvreDhSLGr7l5
FFjtDXiXXgriDPq0KqNG/GCkN3/9Dni5/tgXVDk5yRsAkUlfzUMHhyQpCTCuY4Zj
v+nbJQtvLUJkb/h8epc2lz5ybjkKBRPNNeCLqGGTyAGGyEQEpMu+RTo7H1T/RSG3
PuFnVVunNrAJvXIBjJLE9ULZoywA5mk6tPbVumMgziHkt+gv3e5JJn2+VV4vqgeb
nFCKmJGab+pENqYjGR+b0iZiKOSxOQekp+psS7z1vN9zo6oSWpdilXU4LVCPPwpk
ealnphtw36Q6Ifcv4Stk2T+ouddCJAPokJWhdudpA/g7G4tJm4FhsCk6yk/wWjSY
re0e7jDkZs1lA0UToAV3eSU/acGm7pLNYlBtWeS8ubdGkLmltFhHuWK+H0mKq0Q3
cjPdItyCmw1Vu2Od4izN9sP01oG7ElVgr6mQ0Pw9q3bKnwedv/kPmhipohy6vmFD
4GERw7pMH+OS13hokKwpCoi1PBmzpXBWmyMm//eOp8TKqe6ieLnmV8jGJbYQeIx5
DahCfoqfYY+kMNhw8RU4q5rNwwHABTtyjhpvEqgnTSBGwxrVJVEEobE8ztPrc72S
ZvyKvwhisipg6EkNXWuJm4x2kXycBmYBzAFH/IpsAfkRvWJPX6ToMdhQi/vy0803
LnZysej1V9Uw/3kjSCK+1WveVaNmEkl4gXDmNoHsx/f5ASbiaN8HzK5mHKbnXpMM
Fz745CiMEaPVYu2FrP51sn/P6BOlDZD+UTuHuRCgjpCJbEv6jDHr9wqw5uLftWTM
EFj3Nkwb5kYbQXjb4WwXPg5kSFT/JiekiW8snfuw6aJ4cChBIqG+QM4EbwsKWlhG
y0WYVg6ezu74AvhTyCoKm0CeheGWajQK4E52/M2ot3mrBCDPz4YBNGDFjRFlrdRE
bA0WV+cRKIW7Pg09D8Cw3aKVMT3uLiS2Q0M4ibREDfFhfa9kgmjj1QzlGqTxPQ0U
tMcAgQ5EDOPBJJd/5OEw9DLFgf8y2ljftQDNbyITn8xcWuwkApUgYNwQsrPFbA6H
RIdVPnnY6yPNG7IM3pX6k49+bPUZE1fmYc1RCBG7rolplBRgaRu8lvlZvt785uCM
tmK4OnPoQoNPy30eoT84kDNJ9POoYSpFrJw0xwmq1JaOJ0mbXlPnlWvxFIe1nEZF
SwTGXGBg0zmBoWNYkTUWugP0FrrT241mxKoJPVzL2RjVwPkqJFcpGgkjp3WEddD8
RuazYm0SW1NmGvoDqUfEPg7kVeaPVvpbh2X5FGohDHidTj0raP9DN/XJBtlLql2v
CBYY86N0DuEFhwhSbkHhF2kvWOKqEp+vi2EA1psnm3JBzDM3gmmvcUpHbGNsXZg3
VPXXDgoSTbagKtTqEocPbFtX3gAPziVN6JwrTMTAd/2P7zrk9P0ex/zc2X93OZYa
LZe/xYBfKqR+6IsD3TCh5nMYvL/62Yh9xVSLsLz9UyUoJI+U6ANmlrk84dG6ntJ3
lx/jEb0nCcwgxgMYxXH2acg1brDl8qJ5A+ocVvlRHpJkLEsYPwrTNgt+Hd0372tR
70d+JezZDIisCTvQ9WntjX5e05SMTrhU679hLE08yueSyO4W2rGs6XS7Li5VIL8w
YN/IVUUCjS6rnIhlfyxJhJ4b/eeoRn4e23HCHCEMNNfRx802wPvMcr2uJZd41aul
dky2ZdEPtegdKNRHEOakXwAmRY5SqdjKdMJm/DEWjoc0lljMeWfJlHjIYkfNMGAX
xKNR4LIu8EZsCyNFoylIHInFjhMTIO/9IDJQbsQ4eDPJTmKCLvg/u9gUyypqPSel
R9iw7iN2fUiIbNOoLZBDV/McPrWbs4DeXmMtFq2zclz4oj2Oa9ZnMcLggbaDo3yI
J9DhxC+Q8NxFvV7cntC/Jdm/9begI15k26pKSvfpFL0FbulhW18l+x5a0ajgJ6xr
PmAcOotpoACDgDRpXIUcVG85S0IoYyv4xGGwq90Cd5l6Ll3/ePXX5enn+BH3FOTR
cBMspbbxisBgj2Xwq0f+OHVV0q+aomWN2oBn6HalHZIahYD1E8THwces4LIMPdGE
8yCF2yB2o5xdld4uhtu1eXndbnso8ckxkMpE2P1OUNIJU87ygw8mUR4CQUE2FfmU
2+UPZ1ntDC+Xa7qM5PHkg1p8y6lJ0Ahew7VXm0aMUHHx7BnKhqCH6y7NdfPRDBDf
ypbmVcAp9QSIeEAGk205UEASzpd4zJGuBMuUUjyktf9HjnWHxKl2jHqj4MprYoDu
R8ZeA8C6j7ZRB+OZotFSIjfA2k55utRlUeBPaOd96sfggP4zfF5W9NV/6PRoOKh/
g7je3S5XCqdKUhZ7UKqlgjOnvfLjC6c+OTbvaCuizJa+svTCN1fhQDksNyWmRuIA
3CEba4HjoNTgnyRM4zcjis/HHkUDimPsR50uLyteiYI8+2sCmniVTus5CmvD5iBV
/dZtnLVvIGUsZBkp0kIR/L1RSVJ3RGWU6TJEOWCf7kjrLxCSWt/2PeLkll1INbXp
Z3cdvIHbRLKtC1jXG9MvUyLJLX8spGL1F/1vb7EcNZUhJpb27q/rqducUd8svhe8
u6+W6aC8iin0sJd+4PX52Sty+s/8/kRWGpM0na3LFLAEgyV7kza80/Y9mo3DVQxF
i/VliUATYt1irqZD6laFKKf+BhLx8pcTHIOTR56fQaDTBWNLAnFBDVa0IkDA5UeC
bNSjKR9VaRjFeYO2KekyVShj4ujI8Hz8ezZHnX4QceMQ38l5rCBCBvRHg39MzviY
DFZicVUKKqU2nuxofpBWL01Vn8P4ksJSbghStgwTL8kmKSNbqSqoJgj8sED+eM5g
aaoE2gg4OtDeCVQqlrXvAna+wdC2j/Gqv1oDKCQ6AmMx8sbKZ693Z5PUwrzdoTXU
UiiwpskaScQp/IWTuQFNuUTFv6MZwzTbuLc89fw251E3s67xcBvxXk0qqLoI2lgW
653idpgyFL0DQgiZqaerGfLXdX/s4XV1Pd1yiSFbpG+s/bE8u3SaSOmGlpgaZHyR
eUGF1xYEsmjzAj7+gxzSVDXtVm0EiXwKjihg9r6VgOVP4lIhBsq/gtp9atA98tvN
Ryr/0vXaSDcwPrwsRisldGcKbLK8FWOgmZWHgE9ZtNJjs170nc0mjBBIi7qUJeq4
71ePnWRLxmkDtYVSPR+nK/F1p6j/QL2pHvz0E01xjs4FJYeRM88iLLTveb4DuEOn
0HoI69WFQY54KFEebxxX+PdmUL5Q0gGxHgFzRyXjzYfD2wNVxQBx/dyPUDEbCGjt
edVCh2UtBonOxoZ8jzeLHKJPhc7lckH/YdFAa4/V8imSEEC2OWgxi/6mk1T60yBt
xQyAovduU/TYol5cv4XpB0HNqYaF9uE/dWcbRzv0VVezLVItj0TJrHl7XUH/yPhi
YJtmDxoFjVkoqcKa4zeCREL4g9A9qaYM91MARmx1agrontA/Pkzg67ophg4BpcBS
eXNj861kTHt71yAFNrrDypV3Yez32DX9rg7L6cBhaRtLAGeUS9RLZabPpqPLCUjH
viYRoEUYvX9LtiVgjNir4/XJYFIjSU8lkan3jkU6eCIdKAHvzirD6u8xzi6MnqIT
fTw8raeBO99ZB724V4tpW16k9caPBwMEltmr0eECxg+Mykm23awUdcsu4NbpbC2j
xsbZWtlRSP3Mm5sbB+L66yWWnLCeox8nN009rVWajhGgoGqtUZFFr2J+nXKenFMQ
YulVfrPNPHnY0vrSmj1WnLwwlX6nEaOziL1FPzdlqfseAvdYNvK+KslaARIylXAx
53gVzsyEh15RLVG6m+mP2VwgkHITkdBOgNIOfY6lA0JSCMaFt3+bM2xoXfvY4X1E
rZQXDQYt78LiD1zmNb+qZP7EkypuvyE7RW2oDwXa7KCKKAut3UahTF1jlMJoMCRx
chMkBLbEjAqL/XBayI9+fEuyC4Cnnom7dTLXdP0A7RQ4nlg578d9WZvCnnIHtZ7X
dS9d237zvZyEwUkLP3GQqX04t6tCXPBTcv2o6139MOGuNsGyK6xLROVBxpKoF+fv
S+sIhd4F85NNPJjYLy9/MdNvQ432xi5ZOuBcu+f3WJZ9aW10OwdAdQmJI4bEZuOf
rYli5zeU5kxS6oSYhsL1N4ybWNtOL8eca03mzJNf2PWkrIuXLwqIyXw7aMtNPrt/
95yaZwzd9tcVELOmoPrrU/6D+WmcsDLfCT6zzqMxN3ZEwoyLK1qEoTH11rUBR65A
q7zj7v1lnoA2VmMujtOyjya3GbW4QSvyhf8wCYVyrwAb7h4aaQqb4RiOtW1hKK0p
IIJ+bsBZBP1XlxQ1dhIAOf7mUReVW5IeYbgYU2Ol3BXgRpbLyuSoqg+tE2zvQWMi
7rZb+lbIZrVkbmscQ608DotAFRZppdjXElr190czv4tPiGBO7hUXVFw9CAyubqYz
m6h25F7yuiFfo304wqfgdfHOu9DRuettjR+HrjIZrufoY0LL/SvIRhOFUxh87Je+
sgpA55Y2wFmM6801sbcSizRiBvvuQ0Ryla7L46YF9JLdq4lgGHylCkHhnZHyJDBA
UX50JvqU+3q2Ouq3x7nZjpJcJHEqqo5nT1I1QSQD1XqpM9o8TDaZrI7iryYqPLCi
c9kVkUlcF9RocbBy1qm5gINdZNpo1L/cumzwMls13xXKZw8Y8vBQJG6KwzRXbKEX
2mHHN/tEmCTsBAdhqXqSf1+wmr93ZBdom0NGb/0jy1Ve4Fp3Rin3lRZPCh9M7Y+P
xLQrHckLlqP0CgZqwZKfx4LjLHX7qq+Cdqslf6V2IDYpzUZiueuO1djKdjCZn6j8
EVUaJtA0zUgB0JBhHJ1E+8umvR9HVh5XfZ2mbWPt/7YvF6k+pMFpBM39iTmdesV3
JK07/otIGlT+PANQuPakuqKItw1SLsR2EB2mY9gFrob1EvuL0nJp83uAgO4MHcCU
7Tl1gKeS8WZzUVa1FRWOR7MX5akTKI+OpA2BszEp5xF6lAIkXvw3yLuN+6Ocf63Y
DrNbN9wMKYk8b0fHNMt1vkiuhFCyfyAUrcHo5PdyxZyQbvEz/Hyh4JrMYWf2101C
u+x/MCSK3V/iRPeBLNg1k5MTL/N3E2w8SuC1d9IDsHD1A5vtPejazhk54lcMDI1b
qd4/iJZrnVGK1HN3DVGkqVEavQmFj6sixWIhgIwimLkUEH9PxpxmEXvHikWYybi7
ZciWjIuZ0BA5Ix5APEIlAdGyacEb5oWfZjKMKDAxSsOn8G1lryLCrab3q7y3VNvw
vfB3NkVXb3rqeUSYljsHDO+pdgisGEjUwzsKIaNCXbD+Plt2KuJxnnAGqcwkoVeV
yM9F4CYuHRhBZhxPf2/FsKQObmPXBsQsGlJV80vUbu3/vC2ysnbI6FZtzQ+2EbE6
3yWEmyiScvjH2qDbWcI2X6OFPpn7I476O4t5u5NJhm9PP3X7LwLrxm84Tk5txD/5
6j3kseL4rczQ1urHhK5GFZoGggPjIfsGxgVts1f6rl0cZbKGA/GPViRsaQitQZON
OkAq1bTH+ZxGHAwiJoVF4HbXVq6Ow0ImMCU0H76pVKzYs6MeZ5/oIOgc9ru5ktI6
NQC1EY+QtjlKFnglVxc87I1QqvUh07bqc3CiryVlcIwnJwIOTpilgjsGN0ASgh11
5A0qTXMarbeLPsu+G05ZOYGS7w4jhkbWEoMaZjoQmrXOvFFiRpMvObFjiyHvBGVT
OaJsBQZtbz3Y3xw3hGqhtH/zL6NEUGcdiwSq0b9FmuurOOXUKjmRSogOytI0uafs
YGWV4oaYJgcraSsLo4umD0ys9S/p5KN+kNBWHAWr7XmPNZHFn0zWMjYPj9MjXrLw
b5jTV3UB/rCJ7z1zuyTIE2VlGg6BE/MKKaEw1fmQx1pzUapNevSlcUXbiY020oKu
0uJ+Q98NGtTTnAVycIS+eb0MmkkOZptSP0plBTcmUVVFtBQqI9TiDNPnULeuyZUy
9ADpr5cN+mSqIPoZordBuezWof6NL/Hpm6srYjlbvi0HeTQC2eaMu6XctwgueeBx
bOMpQhtPFe8gZ4jlxpFcfZhTaEjgNg6vMjU9UD/bIPPl5Vy2W18vl8EMGRHjfrK+
40cUOYgzJLaXEXW1ukvehaGn8nM6x6l8hlRrp1jqImZyPzRa0heccro8/CgACGVJ
UCZJ0/A6fW9UVhDsKLTTz5LmD8gH/ZqY8eShHY0lhs8wbwXqCOpBuNURq9IJEl1K
n6tO+xw4YHNesj4eIS0nobdwTT4hfzVvlOYD+XmBjgJbgbTh+vav3jzJJ6CwnhIt
s1pocyVQU3ALw0x4Ofo5crLIHycbROsswVUapJHeyd5+Xvofj9igtFPF7JqMc0n4
V3iA63JRgWesyav9ycMbT6KJI0LcuIeD8T8T49WVzSaEMNaiCCPjzaAMyVMOv7Tf
snj4bH/yKyTzTRptFSdUjUZo5mh7jM1Ghs3/8wjQsHw1MUJFbkQWKJUCnc/shCe0
NWJlpZhnP9qLS1gD1BwAzLlBckX9dsm1L5M/nUNUB+lEIGGBZ9R+2gjv3LisRaDr
93mpQ466JwPbaZEa87fFmW+9DgzjYqWHRZrvS4oVy939ZPJbmK64Xv/BPoojiM4Q
cngL0lxcnPbmQMlP7zIR1pPpHIbztLcW1p7Ux79FhCtT5kWaveMWwtiMElxd7bs3
si1fNuCzaeWc6jIkyf/1CjjFUTVkHPaPwskz1yScLjUTUst8DJBobl9n4cj6glXY
glrVRuC4n1KDvJrxcgVY5ej46zc+SWFF40gssh7CElXUeRzhJZBbRPEjBrvTWBJO
K7Q7LF1XqcIGnZHM/uMOCsQlhn7dOAbE2nmF3I7voCK2/Blwuz8w0HHF2KrGbkYL
KzylnYBVY3AjIBH1O6aSfR8IXbfkAzyHRFYz7jrENAZEwfF1b7iPenR13e3Xianu
WqMbn7x6j31b/R5s5FpEtale0Lu7FG4cOhtAAyoUivd76k4CwiwuKogROx7uOyLz
vndRwu9P4Nsfcd3EEGedHSHG0y7YECnQB7RJiHEQOjaZAuSKv8TUbd4I5mfeqdll
7XTqmUk/AcspFT7YM2pb+l40zzHLWwWtVVxBmD+MqeMYODA4hLS/dH1Rifetcb2W
QGtcsoY9JDuRydqlNCY2jtsnhV5EPgXoCxJ3Fs2g0uI6A5CkNzCf9ukudE1HoGh4
DUU82Mw1WZ+/NLzXz8CfCxkkl9VkSNKWjDhl4Eh0PfvDgiuAKn6zB7tMd2YjSuCY
BD1uSTdUtXYhJ/wQwg3E6TVIuYDMKfvewuFuJq7eQD25djgmRCMONJX/dXjr818A
qh17eFHyCFSGlAcM/DWWDmSOIPZ9D/LP2opxPCW/qsx3DKiZ/aRaFoO3KfAomz+v
2Bo7lVZdOIxZp1eiPjxzTTFfwkde2BcuaWBhLN70H1NHRHjW+vXgvKUnGJyWQAS2
sCkzrp7C44TQNEeXbEN7sCrHv1RaFqUHteNouW6eXoUTjLs5ONdZQERDFllQ7YXa
Zte1OhHZriF+rP6lwwCj7kRH++l53+P46LY4eJd62Uv/cL0pRCwyadReOUrM3xLQ
+wO+9twIdM+o0wzMTA8DSmI8gtuJrrD5M/8kBXrOWF9qMilXLkOib3kd9P5woEHi
xjw8z8it2Lw/eHgNcjJsVTaLCF1d1L5gWVK+yyOBV2W1oNAQ9fxG8oxaQKcSIfJR
WocsodNkWvkXYa3cjVmrEeLRs0yWRaJ5fjRWsXrpAkyle7gyezs14bwQYewco1j+
SWQp/K44On0Plo9BpTq9qvHCjF5oEGXMJFrp2uFteJsTQpVoZu0AN8MQdO7MSnh0
ZCjL9CeHsgefAD9tn/MPl6Z2BrC3l1m6+ypPi6NKUNKVX4sDBfUcZ/UKddXiIJbg
6etbwLFq8GWe5BSkQTA6cpV4GS88U+0iMKVqVHlUfrw16n1v0Aw94ge2pBc8Aq5c
UATpRr5B8QW9el6fdW+TESBVlUKb2uwLS1PVitRP9hL6eh+Dy9C+WNL77VNvuLj+
KRzWXfPtU+cPD0CAbBAastEIgRp9vha66L/MZKrs245M+hTWeAhlk3JvuRYGv6YF
f8pu3ms3Sl5rIgbuafOHV1THUzpbjuZTkT44VO/9tdY7lShydj3hY5kKQv1vxKjk
ubNLWXCAjqsZEJQ8q4aTwazevPyoXhK1GCvDXk2gp55HPiHxkdabH3mrx887j191
tjXvOV9CofeligiGVUgtnG74TyXiAUzmNrHIAy3R0z7h9T5PsNZ1GxmMpuLrRF/N
rUMrPIQ3GRCGvY5n/vOvTVV0xQFqlDbDg09pIpbWlYGibyU2ZY0Uyc3gwgslGGSt
TXtZGFbJVfwmQT+9R7VE+9D8i0yWfvCnBoEgcxFZMxk6rni4g76FMcigzFczKCWm
zpjideJ8QoGH76e6zX6zW67GtaHHonbbfnJT0k3IDEoRrO6tf4lmXp3My5oeaWUm
07MWvA/4Z/D/FfFUXxtKkU1mBaVIY7imgmsqfrYijt4zQs1Ram6gK5BOKp9huQTD
1s0bPloaA6NVm2x6yJ/uPW/15WLs67SvHtpZkWB2dhNqDhnu6w9XX/pjFlT31kHG
JE83Iv3CePmOuX7TSF+TMi6oiPJXa/EvTolk/+NJU7neKWrcWt72s9OH+FkzEtWg
iIn7u9QdOdWFIhymBIa3pEmKwL0JNAu7vZ/1KC+1khMb0YYr2NPgvmz/EG+UkBVQ
xrc+DQOSY5rwJwvXVlwisyHgILCXhSDXDhldVhJQJ8Dta8wWX4g+I2fKItBl6tXh
DAI8PNh4Zh3sERB4sQZgkxx1MCbCHbLsFql0F/D98CdLUYGl+6NjjyuTQ8dss5Ku
IJGnhmpsiXblMZmvD9HLwOGf6Mw3kuU9gvlfH7fAplXAi19eAZBXZaBCm1AVY+TT
GCeEKQZhxpksNBxOOOE4D1LlPcWBUPNvbaOFJf8/5lW5FLAcGg+lGMuC8UWNPSEA
EU9MA5sgIMR9HMzTZeaDayyZAQQ5e4VKA8B1aPgKFV+njjKHaRtYccLBN/6nimJ7
+58DZYmzgP7a3bGppjB+Wuz4BhkVrh7sHrM9jlIhNZpjJNhgB8mejvNb+JYkKAAL
rgaklNfznpSBmzHqL1Nd4azMGdKG9GbA5HZs+W92P9B4C/bt+K9TIUVGqc2fz0Ay
Dkn5ay1iDutIoCDWoV5IiV+Y/Eqvs7oqWykMCunNB1V1KAJQZGASqWg2oCOZx1oc
xqVcpVjvi/wLtq8xA/rqqagN49fewQuBjckzc4BfE4f0oJkqWuCg++axhv/KugB0
UF9Mb7BHH4XsrKeACQeLoIMf3XirI3TpLHmJPcBQIKJxJ+eM+aPfGG5Cr2+5RqCC
wyC8exCq/FphTXdfPf+Gn5MkORcGOk42mxWKheG0MaAGgpBt6D+k4Pb6vytAfYzZ
A1kxKvnOqtYTaC+0VEFI7pWllHevgElj2e2Qi05jfKOl8qkhFOFZyWf7lFRIxR9h
oe9EIgSbgx4rHWAZ8BIgYo0wCi+stY5umT/brGH3TO+h5brsTtk8vN27/ugyyhCB
WZL35GGDL9o3wgyXaMQc2V65l/1t0PdlW5EhnfaRFcTLGt+DQhb9GuShfkdmod3C
363zRrAZeGCs609BVNWF94kDFAclQY3nkAeymxMKEERGO+/QqvBmLRlpdZZ4cslD
r2p9a0ac0L/EL+PrxfP7ylvLSQ7Y3l55R2buQOJxvPRQVUCwYhlnxsHqgeEh6vkv
sQAUZkNRlJHpi9FUgOQFDAd0CBWXgS7iSx6JMCq7WAw1mbnh0SLuhgACb5dUmTsi
UXmdrvB69n0el97MTrUEfTSK5XKiwi5n6c7cqjVx52/4DdRxT2mQ6in/lcpS1dWv
I1ps7HpKvk8WAbkrtByvJko4mfgAhe53lHMCdpry06LzZ1ZZRCKA713LhWf+cnCR
4q0kwydylavQ3F4EodX00J9JX3j0vKAHmBFoZjD3AVwHDtDbDsTlan4L0a5GYbcv
htbt8REGIHE5iXLvm4DPd51gwR2xk59b0TgyEveGjwkgJXyZGe6bwSMhBG5XYjXT
TaDoDRggljqIXFSPaVT63hyN57/t5SZKAsxLVEYosSNUB40vMvN0quOvEBhNYdex
Kk0lGom1SYGWbK2LOmnjFbjDGHEYguP1ovTPEn6vFpJiZZ7FC3L2w/i/2nulw1bD
qAmKsTzM9jK4AAivUPUDPsxLeUkjb24cmk64f5Twx4M13IV4fcio3lJO1WzSoOmd
PsbFIcGa7Htzk8OPNeEUvAy4P3gJgsKCBMNSy69s7BU8k+JInRY/VBOrPfL9X5Fn
bw/cnc5sRQjd10ux6zCvsDN+Vx1lWnyPByIAc4yQWJGuyfkqRyc/q96vdy6K0KTV
RROnPbm8ZyKUXrd+0PrENq1KRtvyBbxqb2VfDKdIiTiBaLm5wqWsDk2wBf7wt07/
OiFOysgcZndtyDJUL0+8dr9MMsTYAddBDE4cJGSLj/dOwkqa5pmwSI0FjH9TeDOo
1rq5aVcsjX0IDh4kGB0tDh4o41ioDYr+WhIlEH1v+qVRJJ4OMjhXZJ9ZN+jTifdW
wvkaJ9lPfE1Lu4BXeDZ08ULoUg9AyVdfU6VbpNh/nerM/mtyOhk2YPOj74eP+EOX
6LZpD5N2S9003IBBTTN9v80zJp+2KHLGbqxrENEDz1/UHAFGfquXaroz8yNeBcV0
0Zo0bz17yyq1fTRv6DPkraObn128ygphAnWSn+WgFYdZZvokpxfse5rgUWG9FlbT
FXfpty6u+mdsu8wKFsvb77i9zG28ta3N2RatVctMchr5ikP2Fy4YRmV00nGxSkyo
E9+R6v6ELv1sphvnpGgf9f+3ULpz3xXysVLjqWlmoyn3U85oZPUODTUbTUF0MvpA
MYQpL/nqlyJKY9CwtlkuscgOOV0tnouJxoACau+9pIXfI+QKyKGsa6stpngOFQVf
ITny8F/xeQdcY4yyg48RZeAp03t8h1+s65J0ylAsn49rZjAREtkkdjVQMyyn/4xi
FpQaicyjgZCGLDOb/uRj5cJBL3G2QK5c8WtU1jidibXedm1NJXB3w1q3WIkoq76g
a00RkIaUFteD7FOwbKmZi7AkKPFbO3Yvw/CBsNZ5AS0I0q65iSVDN5KE8EOGZ21R
sDZsio6gqJEv7tumEWFjJbmHKjIFtuzceSIraroXmqnSZUmpqRSJTKqEcEAYd0ws
vRR3Fwve26CGfNyYnioKBsMS/tuwtvUWxmI23a65IjB1vUpACoygvF+g9DqhsnTu
DOW8avwm791q82f2Bjc6cOGfIuT5rwRf5ByoX/Rim4CfMHXl804ViZMlG2fXrPtp
CwE8/r9sk/XWhbNuap/imVP/doQN4DPIVzMSctkiGVei9bixD9ZQ76c2Q4N0WFSi
dJgcixZodmd0j5Wtm6IhF6bDCr1buE3XKZieB0OXRtB15gBGm7JziIlzCMS0Xhm6
40YAUO3SJ9XAmIMfJW4ODy30RsXHV8nf25jt/StNlkLDINch/PAJ3L2nQk0Iv3LD
kCjMBCeRdrkgeoWcqKwj7++alc8SOkxxD+NnZMGkRd/4Iqetf/pZvIZXKK5wV2zA
XYpt6UR8BS+1scRy7FVRXDAwnZdkTDgGGYPWJ6IUdcg/ECp3XcFjhbft2Ph18WoS
F3mSp1B0A8A6oEcx12r51ljX0S7zTd6IWgOo1LopJWMOX5UpUI67m3eq8UbaLh/j
0a4goZHxMgBEROB2rgt1ngBES3DMA66BoEbsnFn+0Wd2wtDS6kZuhCV/GnzjAzuJ
Bxo0gTOPfWA+y0c86R+6YPDByyt4VxOjhco7y1p7+a/pqfNtK++uXqvCOCa6jB9Z
JCnRlybYBrOMQe8B10ZEKDPFh92DOb6Uk4aBTfKPbdrx8yzAt0iGhFegNKlWAwGZ
iRqCX1qeivwCRo7cWKK/ktmGhCwI7rpfdoDvRo5JDuyrpZQ43PxNGERBAZ+uBM8T
37NOVxrbueFCZ8JOzZl/9Nrvk72+02D66tDKLdLhmVlTGxPFxsIje+ZS8dHKPpDx
6LTICSMseejwSA0SqMysT4eynjgRUGzIuCaBWcbx5PpdAMRahOQ2DF9LEAQdG61M
sz2ang9C8AXnwK9LCdkhY4A3QENylVsPQhE8UoEoDrCPQHDAWi6/G9Yu/y9wF086
PL+ejRCZbZjaXiH9/gjMVw4O4/GGDaRxFimk7XKvoo4rBXsZ7f9vY9L0qQElRcrk
MStlQtj5UpMYGSAafeZDtLkejjVvhV2ONY8chgYWulDi+RwkB6Ths9+Sv1wFcXZb
QHayY90cr114aGpEirhl2o/TVEvfGsOnMAQoOICLqzOidXa9qx/EZ/WjBuD+NuZc
9edp50qSroKE2tTraP73fUJEIJ/9pSqOq8Tragxbsk1VzPwEHqz1reupV+TCnvjK
8U9Ay7cX1cw73VET2Vx29mFyjHxnhnatl4f+z5pguuFs5J5/FPjvIxyCWzt4wogv
SkgEXiYqTpVoIEG2v/5dkiCdT97bqYRRz7ttW7BaXb2fRmax3vQwqp5n2o+KaZCK
7JQ5ZG3MPuOCGBIeP2YxOv8qQWZo6zkLCBLvZHRGa//EyVF3Xx61sZZ3c3iaKugX
7Ui04C3vIuQiOdgm692HQzKp3p1OZL9R2ZtFme0/4MO3qy6O0+T0Y7SLhwkn1eJP
xlPUKjUHf/FhzcjRzkDum6EZ3Anw+scvPyWWfukqn/hj2CmQtoO41MB/lJKcciOw
hxBsu24fCSWBiiD6HPfrF6IyG2MJjNmT7Ib5p39b5o10hhy17BW3lG0Wv7FOVA/U
ECJslP+H0I/1Zn/NrQtlRKmNFtJM9ErVhlW6CZ5xI03gboYuUBTaAILF3XW5oFSv
aQi/LvRyyLc+46mZLxq6P4GpPPyo4LglACJXLHp5SZ+t7R0wpq7wxAL3GCWAl+Y+
wguoOjn50jVYdW1NV5zg5HpQtpYgvvsOr9aiNl0mm/PTg2WyJ57AN4wC764mWM0v
PjWu3jCNCPq2Y/9JfjdA+J/irLWNEw3VXnX3lQQ/Y5AHx01KFND4EsH7WKkzIIsz
eVswwLkj3hfhIqK6665XBjJirRR1xjmegBhIAQzRw7IGJjEHZxaPjg5eb7lVkgFt
hEdbokU9YiFCvGDBr+oTr8YecUBV+uB1SQCWgabmUuor8QeY19lUuY1QFk4ewG9U
YaWoNzctsfiJVj+4ForMbf0IaKeCkYaJNhmy46aIsE7xqqQO3IaO0+rUOCF+r1rn
EY2yOCkCjxi/djZANn7IbvtFfUDTadZnPF8QaKsMGCq+i8wLF1m4i3X+e5WVhLUD
p5S4eabPtMf8sWuaZloqMVF8BbrNvbkmsMDeRRDk5xVL3GxVsW/leOyHrRjmzv/n
vdqiklZDL9S9HLcwEgHyvwQO7AaZkZfH3ZGEwS9JlKxN8KlE6GV/YdatY6IJ9PxJ
DDsllVBZXzaYNzpFYQepyZQQtKFr/DnGMiI+l/JqOb0+phjGZX1hH4B8hSAB5+eZ
V5cdAZ3ommQeXsh9MGIYpGBt/1yEYricWSkYaSCUwgEhOl4yVG/WFoGz8oGnLJuJ
iwnD2gGTwgZLZb7coNS60V8XlGda4RIh4jfRk6timCZyIbURP081MY++jCnjcPzd
mbMz/uXi6L9gaGFXjUpg2YV3XwFOvzcC57rBKv7co8D3Il32jv3iLQY4Sj28+wbs
TSg96HY33dtXZodnF1wno1M4P/JzAmnIAa7EqXFZgN7ggUzBLmAwZziI8XuJ0F4V
GlRg0RCazE1Ri172FGOpue2UfCMtPwvpYFQ+HfDeoEUyjzOIrodsYmfzDd7CXFtX
zA+BShB861crxQNgq8E3m9r9eXk0iuWdT7AGuz6FXzTupzzzy/3N6mjx2huECdTq
LWfbGiShFF6DtTszh7zRks1g9UBK9uIv6B3bYQn3ocvVQvWH/zmEF/8DmrXLlsYV
rVIv+XgOEFn6Mv6zr7XXeHR+F/IEQ8UWNtDiCEnz1zMChik/1HqyavsMq5apky2Z
cTuBBKIrqn07/npm79VYrcaUYOMAKnjRk8kSPC71jM+KAWoAr5gwul3IvEFhYGUt
jPnr9NeGWIqE406VHG4/hVhAag5817U9BfHybVcbcN6H2cXahP0c1J+jOr6isa4F
IJ2asZ3TovjIUEbXPuglShueEZ1w2AaEkunoCEdeJJISQo6QvelzKriGWOpvlKRQ
dlxIksW4EtppyKqwW+i5DvynU6/mmJjY8DZM0+JjoUZeHr6f2qecfeiEGxywHZna
vlMd9236fcruEIvLBLFLDC6fr2xXVGOiNp18NoIZrQIWiKNCzGp+oAAprfWe7Y+6
85B6euqCyLkKVX7ilhgC9s09KQ7OKWGsgZd4zJlm16b38VJJTw5bc0lDtN8AGULe
TJTYHXhBKF5EPNt+jW0/Lu3ASGxFWfXUxGtpsPE5GpUjPXcoQdAG8vyZDzKekgXB
aNIIYNxI87IxM9BMFl6qpeBT0asVBS/axW9q5W8/cs5gPa/WPsRCPt4tMWmGsk2s
JkbvB1YSJ8om+Gu+ymJXHJHFZhwWURQVnd8LYAwsIjsA90s2KqTNHjDpL+bMAW6G
FGjNsHhfbwJNbxbRNfvNZezqhLKwTKB3vVs5Ru1inbfKeSNBdRuGP9v/RcKyfsyY
IwZi08NoUKCF4j8mjWM3SBK7GCdvU2P9EcDP1z9GfqrsPFtQOLVKO+1iLvTwdLEt
QBcsMQ9Pr/O80aYpSTkqZl/Evxdw0tPq0dhOwyDwpwdqWGB0XXspzOZCnisNqAiz
lU0I5vMkfSykjdru+8/+Z2QXTgZC4+tdK5m1H+qM1q28f30bFdXT4U6TwR4/Al4W
fIHvKDynjaQVN+832E97MRZ6AN46h/XdTRypk+128VUnXr3yRK86Lrk9UCOvniL2
VStNi9WHtigoqsZeialrdZ/6JEEy7nkQBmf9GSPLo4uAjK0k5vtRFibcvCic7H5M
RL+u6YUjjOuarE47bsV9lRDp3cF9nWnTX4/9OH4ekEJOiJjwHBalCGJHQJd1ocnk
iUC6PdlH1e18QazSl+SXr1Mzz6GzmIFwfnhIjpcASiMc2EyoeqoKksQpHrKOKTb7
lltHZ5RgasN8HHPKxPewD1OxdNyRUA6GTEFYn67deKDqyryUiTVERb95LYBtZVqn
u+mViJXKT+TbzNWVDYRVasL0qw5UIZqdDo8VX5jsQ9QLK7+PWpH6wyz+0YaUSrpZ
5iLX07CE8V6lcKzpiwDtNGq3vdPIbLRnwSeD98W9FmRhy9gNIMlqYfI039Gr4bz+
eyk1PlijfFzkaF6zaRvacjxNZzpK9SsQsjxhCoDtoSvELKQ8npVFzBOsSfQeuj7P
s74a8qhNMx/KYaB2qljg3xolL2BffDA3NjMyFIBIb6bnTZxPrKdPdxet/LEn+3+h
UnRe7uF3z2OFkBvkmHpRrEQqJnoS4EDVz5QX6azgHcF7eQO+axxStqH0kCDhzPMx
YzNazjk9kch2Pb/JvRXupaJgAkAwB1PRmAuWwuvxy2GOktE2Tyux8UH91p2uev2W
zfdM/NxkMiD+Mo/4Intxi7tURHimDAC2/vLsSUZf6/oQ2fLigkwjsU70iFVncZZ1
Jwjuk0K1M/BdVij1teiJaQdQae/8oVAxHVW3QsxOJ9Rl3/aE0XL5YuM7JMnZdrlc
b5MHIXWKpjYRvVQq1CpXbpNgHyUfsricHa/Nh9s73NLi6k6LzOdaNCFKNkohfHpT
Elsr/KQwJ2u6DMvvqjfL6wR2aRX0tpgimix3ySLwxV14m5i91bPfeUJnxCi90v9I
j/2OstnC/bVnwLs+1F1cD8arsNIQ4FA9s4WqN24t0cktj3qegX6FSPQlAlH/7WYA
uLWYTp4ZT204k8uQH8zQPg/dxqud6C4/d+zsSPdcm6UynDEFkghzfLw7MC0BRctO
lQQmFTkLELflDNrwq9gMpgfiZ/9MmnHldZVPedxCweubD1C19S3K7oZPldzv+1YS
DjsW540GotiJUNwWL4ftNq6rp9/UjyNG3niXhmlawy7TuIZ5EoR7G8seP+IRXd76
tjA9UCb54Pj1X45938WwKcsxIKNscKGtRx5CiZd3NnPtfE25n2Vo+NtitbcWSFqx
S5q6OI09BJTYBbwvAE70gGBq39/ht0vzntVDv2K9XYpXQ7O0bdfArC6XKc37TCmE
dk7I+/F0UOWCKdOKELnBrDQLmofuKq+1Bq3+Suwl/e2MFZiGgbjAxLPEpzw5x7Ym
Ker+lc4VmqSYy71uj1wUoqtjT8AL3BhK4KqUIxvdUjiOFRNhJtM7OOrOhvIoljjl
zOueTkWcToSZk084/fZ6pKMCVGZAhiL9tfj5vzsM6nYsUDAkqKHN/wMdkS2Tir1M
HiZCMOb5i2pOfSaM1Wjep63tyUvZJ9+ATs64A0RYi9qb0gI3BqJ5UPymTLw3ARN0
Azi8C2vQFN1tT3D45qo6GD3l97EziiJ0C78dCKa35FlpHp/pmXuaq1U5qtaLEqAL
6FUjJ7If30x7uDA0zKPj+Zn8I1Cg4FQhpbgyh2CatlLO2L6LYPX0nSiZqTOb1v8N
fap+sOkoXqE6oXMssVZvOvsdku9c/FphTinJV7+L8Qpp8O2obdV3bEWV6/vSAyUo
Z5wGnlGkRd3QpeAEoyH2AKwLf9DezBBVo237rQMQCJgZR2a/QAsuVYTrhO7zW4Xr
naGxG3DGnwX53TN7ABmvIs5DyNs8Cd9IF0oxAjVqFQ4mKq/hJGV7j2W8b+QY3mz1
ilHOOm91aY9ECfry/72TuaMotF98t946LzrGNrigw4gWRf1I9hAmUzdrWMmeB3Lf
BpnMc7s5U+/ZK004flvxeAgUu1zE4DkDJGTik6NLszzblQkl9h6YNvUrt/MAk28R
qWOrdZz43zYWCs0sMSjaaOn9eE38Tt/uXrpK3ISEUGQ/i6KQzmHtNYfnBKCrM7iQ
JMma5bTHTuk11iWSYhLAc0JKPYTxj3WjJ9rNEwHbeZCG106Br/ygepdXOE+NS6RY
502pD2KKmm7CEKzll5WseUObHRHOvzA9gX0fyzQ4qlKpAiJev0GFkx6qPMZZzUDn
swyfJcSQw9A6Dsfr6jU7aSDRS5JxD+fsRFbJ3vXyz/j/vGnqBgX++zkf7VPXTSCQ
XNcinWakpklSU5+Rux3T+qNRKV3q6BUjGaN3Z58kS9r+wX95NtDWHJkmbr+Vb/8e
PdFYF5R9IyT4yeLejBTyMTFaZc1IDlklew9e2FTffrt0lWVAeYH9v/hwtirzEplj
la2oZhfVZurrc+gCzJrgTDFHADQlTE6o1P5loOeB9jY8kDQ9oW7UCxE0CzT0NKCc
B8QrN2Ow8gPDzZDjsEwbYckzAO2/l/7jPncbR3qMpB3dm/BAf79QdFHxBO1Mr7lo
HOOGLiDoHJA0pUO8yZVRz8o+u4b5YrsV2S6lt3omVOgS3Cduo3Eyvtnkufw9yyYi
mJ6MhoyLyG2MghkBcV8mu5PN9VbCJufGYhtIvU1aIN0aJUOPqRPf/eDoaypjSkQT
W44FO0znY/JrcyDvPvzPoepG6kMnQ/0K6D9+3vNPD7qBQ2HUTdeJ9JybsFd8lJJw
03/3k10qd5AsMVL7klIUEiYiNOKOV76Tgyqdee9SCZboOuk1Ylt+Su44fiDlvyHW
BXoDzwYG2XhwRZ5xKMWEaCyV2z79R8N3BDYX31wtI+y46ZHLVkfylSNY49ImKZKw
xBz1KyAAcFGTl9wEfB+MRUK3Yaw45MURiU8Skbbl7IfhA9e2nyHTwYHwDXjEv9uf
luo3omZ1S8zIzWSD2tV6pf1sO6Ak9AHUclpLCHPv9qaNYmB3sF+LF9A97X0bwo6o
/IVwCaPtOukCw4ZesXbQHzJGH4MCWy1m2FlOEmYyNU5+7N1MWAYjSxX/rmO8rfPI
nCct+eKFXogj4j7x8P64YybDRYG+eInudMWbyi69p4SD3qkuEicWO0iZ0R8AySzV
+Gx+vBhKlC1vbyYvT+Ir/hMVgrMq9ASK77bzVb040RiDyqui2SvhjDc7SdIIio+D
lxxmE/6NR9x2E0nW6YLfxZ1KJbhRMox7Ax9Qj146CZ0FWzy0aqRsKHNpXUf1MqIZ
XL10WWNJu1X11ALjKIP5CtOPbEGfgssRSEmx6vH0JdWtcTR1gPbbKvfQCoNK6mRV
7yiQwFlsqH19y1R+Y7rGIuR2AtVsjsf82ra2V0BVm8EzpYqub7bXCyyQEJ1PJdMQ
G07JhNQrGyqjhwZu3eE3OPhUT10O9/Bcj7g9lVw9h9rINovAmHyhKnBsWeRhQz6V
iEF+9BvMuUz4WYi6rz4uQ/8JqgcqJWUy4Gxjoi0hKwlvsLPhxxh1l5wTT92XMee8
P/kTZE7D0PbzKgFEjDMVkonmreE9LjC1b96U7O1wTzbf+fsCjFpZ/Q4oMRKX10tB
/MMaS0oWIb+GHmDVrdoPWkxP1TvcErauDWG+KEs667zVZzPNgaTDy1T8IoPtQ4Ql
dO5BNcJ8rUx/CBJLh5Gwqyu9jtN0aqcGNbvWo6OK6eGPIzQAe27/mJhvTg1M4BTJ
9gmPRhHxa4wsspD91MuAH55tJVbBdW7DpfI5CCfwWBfwPYxJRMqN/dUyR5yFh4iL
SYPeoeiQwgeCCmg+EEwk89iTo7HbeOV22rta4FabM57C0HCbhqLapME0u2clfP0y
8fmG6FIR4RVkHPZACyMrqrszjWdMV+nGiuqYK/gHPbDQ0ZDSzXjHLYGq9qqNrL3l
g2NVD7uzIK7TAsBxabAh7fRYnJ9V5MDA64cg2tCLeQ7uPNxWo+P5lyFWdOoCbBN2
TJqHfuJ2yfMeFwtLqOPhoMGWYK+BGT35f5SDSsEJChOZTv776i0WKNW1elgqHqIS
gz7N4dMk1XG56uDz2s3lNcgmFVUkCHptekXXN+H/k3L98Orhh+xLV2DRmVQLzR9Y
2hE7+IDRz4VuNzOcF87lXmQ2tZ96fxiJYx847hvKsALka9RGcriVz81XKOkwrPCU
toc/6aA8AJd66Sifibu+iNdZl3sKEfpdH2R8o8uOdBCLN32V7EX1BYU2xjUT0PcT
RgkjiSplNeqNytsLKx5CtA6BJIld8cKPrKxTiLttsyTcbK0P8/1WEpsOtw/CaAxM
ozHV5dKO1xTGgCVzOFjLsl7Cv3/QLL2wQ/bv6OUJM6Rbha3ep9susKNDWQPovuOR
VoItxGq1oQWITjVs0Xk5hv/f7OCM/la8b8Vc4j005JTxBAlnqYb1cP6BWYlnMkkM
45tW/BEaQC6iUsA/2+FPS9IW/OGjLR3h1p1P8LR45FRo0Do3WOV9FMSkBqqhybtF
Cc6ZG1eniX2CcoMp2NkrHmv9bEYRqag2YYsrx7c69YI0JZFtDR1TXaIbtcnzeeav
IljMAgJ3jH4MkPAImApjwpHzIzkcS07JpG8fF8xWqxNRVK1ylHN4crWncHArjeJz
EUKbb0cpZanbgiewgbX2Pbdwm6c+9hiCvttzs6eCAwMYgXW0U7aeJ2GBoRD3OQxk
s9MN9dmh28mJqZtJZ/ykpaviKz+demiDRdz+GV/Qh/2DnN8haTPrsxP5PxZWLZU7
P0J7riooFJNUzZV6ETOTsEu68vM0H0hprUHaGQQqvnlAqmuRI+GQiblEs4dJcXmz
4fOVh7zKohlRpOilVverQty3Bnh0WViRUguyx9QHngWbyoguIit/rqoOvJOqtsPd
Lud39M+ch5C/rBz5QmuglCXIGlb0ayValcSzRNHUXeyj3SxP3uDM4oa0Xc++rAm/
KrDDGQ7K1VYVedPA5J8JRmdPO6XQ4QCxnwuuqEe0KweWcSP1aQ1KL8eguqKfJ0mx
PrQcFOJRozHl6/6eFD52fKJvic/GgZwbLoB/e7eogI0hqnW2jrwir87w2SxkVhgJ
M9NQGC5PPFnpgfkV++7C1QjwlDmPH9R3mFGX2i236Hc4Xz+qbz59toP89FI+cKDL
WNp6xC/NevTQRbPgr4ilxhdXKYdii3TtKaGi/iVywLL9JexQyqPxRTZMbYWZrPKk
o6iJDwBQ5xlwM7tbI2S+DD9eMWjF88tPysrAPZK0DkCkyXlmPxhLFJ3WJugiAiwm
y9PJ3HuIu8SsldZ0jX029IoVikK2YMTvZIYQ88W7HkP8FvEqToD5EjVD5K2egsfd
vFR4gxru6qM25S0XQATJcQpQkhsWFGbGG+he7EY9dUiKK4qFB83JtAfH3XWlVms0
Xy88EpICPnUxsWA+69ogW/8AU4CwSJW4koQ8IMEh6RYnS+z1TVS/Vwx8hbFmvEjW
4MF13cynSzV2nXnhymQzU+t9YtLVfayv3ZZGts28wYv02bOLdGcnN7ETIl/wUV07
gcUAVFLLophizE5YoPJY+kDn+eUMXcVGnN89JbaUBJx5E5vN6CtHBKAsAR1Qtv+Q
nqBt8T8CZ8WuxcNYJblS11rD3qmdwlWHa9W2OdX+lge06KkpxSVBPF5fFMS3l/wi
rNSoFdMig4rD9rBLuIYGp3h4qsyAqNVLiFjBU+jJTpyLFjhlfboyIBtHQ/jKkuD8
Aw8EOyMKQ7BCq5jxbpA8dlTvncmbv0RYNu9dIL7ROuzh4pQcUJVZfRLnIXhegDW+
pR2JbyGGpJ+IAJ6fxBJ9buoBfiUDBq+GR/It8Ma/VcDQENw5KVwpc/20c4jbuQs/
IJyY9PIqAafNu6p/1so1Gv/YUKLccVarEXCjQ7o1azBntn4OnONJgLgaDd9tXe9w
sL8A/3cNRaqH+/FDyxSVmDGu8jjFwwHQARVTSW8wAS7fe4sXpoI7vqY6NxpYuzpg
4wRo2XmeVFKMrfE59TQmIP9lH6KneOXPBh0ZuTFpXzuqKY7OCzYjmR5PmGhTPhmG
dJvDUZfDDohPCFWmNza5xK9nv5S19YQuKHwd3Q5TshBwciqyuauDFIXbjl1glm9u
6vip+mFeAr8w1EHsbHCcNngjiVFtnjNbZZ2WSFMmGve1w7ffI+mYU/u8A9rVrhZo
QVb/m+17LETJ2s17EuiY7+JPf0OMcHfNHiBaugxJ8NYafFcsgFPBjuiStfusI1GQ
cZBMOa/iNk23MPs8k/I0cfyB0j/Ky3r2Z85VOg1xJPp1XStCOaaXyop5LhaYj0Am
MzcFGeDVSKezSVloj+vlT24k3i55pd6YowqpAcpwhciGASPDVluyNUrv5U2j7Gyk
NSWKYqFco6arzHRyWU645mtkElP6ABlMG2yVISrk5mwDLSwQzu4vroPlS0IUmF0N
BtyNCmEXKAUhPakXcwEh7OSsubSn82TBBRBLkgLJjgKlYxEsA02+NqcT2RkfxmS0
q7sBCCYXFAO4VB+Pwr/akvr9aUdO+adk00yxKzmqf2PTlLWkK3W40ZnGzRoji41P
3EKCf1N1Afz3cNPc5ivxp2B6kQN3/sdPQnMx/+4vNyYTib1XU72rrUXb/Aak834v
3JyQhSCNBA1FBgKoiJHqFxHQ6vtT6aeQteaSJuZtlzJkLPvClNiFpTBjtBIIU5Kg
qthB2XGH/rFgbhjZfOnzUNmAJPAbM2pYiDz1jxeSszy7R1oT9EyGyDmXGTo7/Gj6
04GNus/VLG1c4/rLPD9+fWCHm3Yjx1fNVZejYQVtCfShoFIOJ08pz1vfk86idfNo
ujr1yip57fMycDCEpizxRvT8LUrhfE5YH+uliAfNUpCakAq2OBmhd23vCIWPglv0
ZHwcROMFBegmNVSMK6koopYpV0oZJepQn0WC0wGOji17n9l8vnSBnFxHYQGx8JUk
3cOu+SkUp9XXvH4ckbWqFe1EkD9Wi3odgsALJuEL8xEGH/Pl+jSF6yhkV8ddjjY8
aystcz7/nK0FhSnLHus++qAkOoYm5rKReCiRKQ9Qc0PWjhBGBEdPmf0hqF2yFzKr
kdvfEG8PXfgK8OLF2gyowB13D59dw6khcl526gGuyEvL4hvx6W3C/GJHfUv7sLwQ
WAkhfFWNKLvXFbsVpTe1DosAKjTDB9aWrOqlT1ipw147bAWzHbaP70YlslUzM5Pu
SfWUFENn2U/rpOUF0qw+q4NG9b33aGxOiRLdVA/jjqLuf0wwVXkGk/d6KJnTyRLq
7D1q1XicsrZVyIPOn4Nd0SLP0MZ6Fto+MYuDCuI2RA9ltwWo808VIzMFJkQwM4Y4
VhsXF93lcYKME7eeicqnO5UhOzvVbr4w4RXAWCcWC3QKZDrdzWMLOOTow+/1jc0R
gEPGmgmeu9UdA8K3jcAjRa2A2vOg5VPBKIa7cCKTRnO7KLPgpmv2XL4nrnKIzhbw
CxqhuxHNzipwc563eQ9zlW26PWa0ssKN8e1DlsX2e12hJ5on1L5O7RqEM33Jf2c4
Oj1WDYtav59lyND1EA+1Wy8hk/iHJ10cNx40xDjzWxgAFu8P331Ge5p6ckcVaKx+
QJoUja3WhNmn0MsCgWEgHqjAHaWcjjs7Oy2l3RA8BYdG5CIobBjLtmfn+IraX4a7
VF3d1hPG2fDtjmQmXuIPrSVJO4kGKP7IuQryNDfuzKtBtgHcksuRBrmy4O1++eE8
+6xxnNuUKyYH7EVv7RwH6R1MbrazqcYhYRZa3X2ka5m5qZML/j2YUxg8VBFFoOYd
AMRuyhAILmbOc6/49LN6zsN+4QpxY84xl7b1JlDBK0zKNqHCQv1cU6tsAFsaq7Dq
izJ909RqGEP6uoLn1qj5TJwKNZ3bN/NvYE+8IzCAT7yZQxpUVzqFAbB9IBLXiELO
y5kQVjK6RjHAQOzRUegS1v8RCVZD2rGqvMupMAfN6Olv1BzQmmIykPoVqB36QbAT
9iYmis0cybXCpTsGAvQ0NGR3QUC7llYA1uZEBjwz1FPQT2ULbV9nLC11OyT6V8qF
SziOJ8b/ezzpPS/68jsFxj7jagwBdWiqvig9uDSJ9BLUVKkaEsd6g+wFxAujKzJ+
zCqYeZ0RHkMjTCoZJ4K5a9I3dHPr2iw+BGCMHpVFQQJX2YYQ6V9sX3nmqCK3oLVg
gOakCkvj5WXKu17uzLVDyU0tBIfzu8L6xhnYjqQMxeAXe+S5wxU5aF/DKgiL2pBv
gSRaLPV7hWTg9ijBG4WoCI0wGL8z4dbZQVcBBn/rqymbuLUbpSiz4sBp2d9RqZXc
encSNMAjDvE6/trGGHMTr736jVhUeX5wjko7x7z+MCyVH0JGmJRxIseOG9aDIchi
pir1nKnDaaymx9nejAPV8EIbfojwIzM/gB2JBHMwPxfC/j78bPhr8PpXhcWY8ILZ
Kos767HZsu4OLCouM/G8QSmkQfI374xmB3OqpxIL2/dJLcH6tNq3KlXaXz/aaDvu
TCvA5p7LqQhe8WNAcGd2Z6nr6LYnM3jJmtFWvQzaFMCnWA037YcnRszayGQ3+EZ8
D86bd7TbQ/d0yTNMJ0c6Qa1/VSzU5L9u5y6b8EOQhfEE4arKxUueeTPT6ZZs3D0Q
JWN8/vPI2J/b0R91xHOscrFk4mTljyM1+KsHCOFXl+AXBcoywnTigjKxyxWnqyax
4GUv155w8k7WIk/aOdYb29LW1f27R1UNLiKxtERYbENW0VXQkPBat3x/ht0q14pO
j7WYWuSQCj6lUeRHFnsPfyrlNoIag3prFl+fS0pygccErxdDnwpAB7LOq9iAij3i
fufQXP7KLO3Z69yUfMqFXGa2fV+AF39wSyuQBKZjMvZYqDUTU3dECoiX2fpt39qk
IfwB1tn6WulqlHK1SS5jN/25aw+Kd9vZHCa+LeSv0sc79onRo0P+NKRJMmmW6H09
n7IprLk5AOu9YPW0FcWUyoZSP1TlKJadfNPcWVWGukvx09dL3ict7NrUY5sMYwSI
J5HClps3Yii+xi8hLMAZbX4HIKQABH74cmDVtVb8AH0/cz5Pr1PZVKxWWuBDl8Bn
3SmVAKwdWmVfm4G++BwCLqoGrJKyc5QTU7wBDhUnj73uWnPggFRxU7oFMWFjacI5
yZIO5K2zCv442RG76ulli57HEdwmwlXZE+3g1JBxGGo/WHKWJ8iZqo+vkqgYFYqz
5crw34cGqyL5HXerlBE6Lyj08qYJn4Z0jAT5Y69FV99UdU9qjrKlGvJzoegrEycn
jBsxTJZK4MmYcvEWQ7LFb4+V4U1PkDRt/UIM2OIh9hcRkZstJX6SIOV4egBptwx8
r2IWLqK4sJxtd+M594joLR6gCj9R7CGclWJhZ3dKDs0bnUjIwm9My7PXVV5aDKIw
kvcb6GKlB9pBCayksydcRV5f7TwqDdpPck2e1zGN3U6v3Xvp9svhViwlq+h6UnNQ
1PYG9sJ7e58V6NSpmqgRbrArZUcuRBtR3Ona2LcuMwJcZfW9wI/SLqFRHNVrY0RX
Yr9K0QivBKc9R4uDsZvLfPVFb9LFRKoz20Oha6jPSbhaZqvUV/8jmzZcr8skYNP6
3BDi0X5O6OKGlOoqyERLV7JLUqiVrAiqzcShTygIbLjNNVu+F+YHNnDAruLa02t0
0B6/S61Br1mx8oi1XwKlQE7z7Y8bazXuDWLKBL0VCsPPhuBlcMcdF5uDPIp/XCSZ
yJlcW3qAp1uP6KI8bBefMfsfrdsEV2AMGNLUQCMJjeMxA8GS4GXrYOXaUAqNTluA
EAU2A05Pa5c8oL13cypoR/5jJZf/dsyFo6f34rFlDjmp9VRiMrWGXjZyHl6KeRUI
dcwGu2d/TX1faAL50gMv/8PZ95Unh/CSUzFS5UBQv0pQlYkKsBQdDwUBQKEEwMNF
+f4H0fr7CjXrg5LT7SDT/DvOseA40xOsPQj/Nu7sSvJSjwOL116Sz/DzxSVg/meD
RPqLY42Ah8EZl9t8bwPaiR2opXSx8tqUaYh53Z5wN9g7cCoMrhE3in4M0kw2EoBf
d1UM6UYail0L7qpshV+QVbMvLMxP11luTUohpxSFYR91ew+BEV5gJ52kLptSU5lQ
rTl9yHB55T6f4QoSkHHldOxuNHhAmlPTJgRUgm65p0ExO/46tgCFtNzHWIRKPIKg
VHCwXJ+yrHf3GTSg2D602hEykf6vrLfgUGqUHnkwpcny9UvzyV/dmq4vu0+qIo4b
ATFyaHwziforCZTNDUw3wMGnutgGtlRc8dlubW11CbEZfY4WS5+/4mGIl0CA/Wf+
S0vjEHhbMTE6HoRPEqAr8/s8nhJldR7t3w32p6WUYWhY2EGZSi1WEeSuu5ZbNxFY
olE01l3gMOoIwtXXCocqmXG9feIxT0vFxf/x4QrY6ZFAc79Md1vdX3hMbN+cqdMR
+ZlprG4vkCWgzUUxL3wMAqReqywyyhm8Q17QwHt3Q/hWARSROlDaBQeRNw6gbRYl
qlOuks/wQtWmxAf77/SD9+FV/UF6lriR5go0Rip60Ra/wTzhXmMGq3zq6CdSkqfa
ryEMJXqPEJDx6i4mOCLWznQCA+1/xpgpEDbH+44TNHbxvSwih3tn8NZW+s1N9eki
PibzEcMBX7NVKPbeFki3wRqLn9NiFG2INsYs3upLqN5cEwtNHrHjoJgut+gfOK5w
HBCMIgXQJfkysdpp0udAQ3Avq4BGAVumaveg7gDkGTZY7eb6Ahy2gkWbmYZfwb63
VLDD/Hq2MjszDkcHef2JRaBFh9FeEw0FHZy0UrxQwsyexFPjEQjZO2GMA5Ybyj7f
WeVfVMe93xN+dQXdT3EODAdA6PkgJG8TsCx+SUZU3u9etgr1yEHjhQrvXV9Uj/UT
5HLRnDX9/a2Fb0FYnH2qEAasRNsVO5IKN8soUwN0AmkwNYGg1dxQ9Z5l3t4vDn8v
b07gL5G9hTdkORhxiOIzNIKnF5vZHlMmjUo2O0+hEcRjOjIrNiuUsCTfEQq4W0Hw
0ViG1h2nUqd61chhPy1AD9GWygYssUDc3WXz7ws+bwBFN5zxbmJrktr3hb8OHx58
0Xv5fE0mkJ3qurQefqkSHuc4TGcGIHfykQZZ9ZBHaL6RQr+odSG1ogXQ4iGrjGYv
nI4b7nhpKOM4dApqvtOCr4S3sE9T4HufhLTSMV8Ubr1H6e/Az5wORHD5g+G0w9c0
V7MKBa916mfX6v98rrBuYgBmB+kruQsoMIaEl83HY9pDi6KBK/xkEs2qA1M30I49
s8fHwAaFgZv06OhiIDmVrB7xUz0d4rrhLHZvCt6/Hy5IH0+8jmhZjj89ZS90odIu
XGT2bdBcWnaO5hrQ/2Ga1I4QSSRYHlMZoApUWFUYbbOR6m2Q6egYlS6A4Z1DsNLM
TUKKGolrR0xoVJkNgT8DI3yWKDDKen9axrS3LSaWfNhj6q74Ofwqnw2XHPAK9V8g
vEi17ZtWU1eIAfKWC/qzR7fXeOejCMv/nrDxm8mb/9ctvD1cDQD+3rEtdsRey4yX
q6d7o0yG+eP173J6giYD2ee7l/jS5toHd1lP/wz9MLssLuk+mLaLhPMNxU1VuuAs
tjwm4wJDo0KWHwUaCO4MG8dwz+NN5TX5SixMaeKPkNygrNcEfmesFdmWKlst1Qqa
/M/QV9e/x+xUtwrYzluhJDLuCoL8KDB3Hq2qkFN/ZtuYtHE68pY308aHIL8uo2tE
u0vbKbK8H9/t8VgmVEhZsLZ82EfKhqazyENZbdYG8ROxmw0e+OMmI4ndcNPuDp1C
B68gv278wpWyn8inKoWUb419i0QBdTHOmInQR2DA0Cfoq2MlsaxEP4HOWbWFyTuP
+QJE8P8Kw22gMouEt3vzxkx0PfySnLxA/oyRMu6Z0UlvguyJQ2FJwX4KJl3RE9RE
P9LlisJdUUIUJI+VcmhTPdBkG4d9fep/DCYCca3ka5SE9/8hBng6hEDC2BQzdUv2
+pWVRt9+BYloPr5QnlnvsHOEJgspEw6hqMuonu3E+x/YL6a79wuLi4M+2ZLsV89B
5euW8X4Du4pcVvH19GC3NJP0AavZmvJJavL80q8j7m918slHodo6uYMotKHEqWZ4
rcSmrf0VM3A7PbtCImUBxyUXH3RdV3XChVurhrSLHz/r7ZiPYNj/plBj8sqZRl+X
O7eKy0yVhMt3nu7hjCDG/nGYjP37y56t+8jSCYJwPbpxtNMp70fh/TYwB+K3pVWl
zZruqswAJ90fIGknh5M7urN2qm5fOBS5gLQmhynh93wytu8dO5Fx5glI6RHf9EtT
K2yudsL6Jj6QjSRPhzHDXe9e9xj2s+sOvvgljpa6mwQ5Q9E06d46i/0kLKw9aEsl
6XzIhY2TLdyGeX1Rg24S+b9HIzFdxzVzJ7u5kRvnr1mt2TFcU/1Wt50MtUEEVimV
7CwL5MztDJ2eSvNC0yTLveeHFKQBmfZn9ZJ/NiEPwZcRXdza+rfbKypp0u/PKO0K
O8FQUN5Z2XG2HOwwSFzePcB2VdsZyrFmLIoa0juVOastzunvIwF5vVScGwbMWMcn
NfuaN7cNzMj4PFP5zwpG6vFgbEqlBIgIwYY/ZsU9IG8FUoQT1xpRYGeAYCOlFN/i
hSFDxywiiD0LWaRoLcfXATn2zeQg99j70usMbdHlc5TINeiKZ9jC+J17YAU5hOZI
LB0stDJypQx7yGL5b7C/kYmIHr43QdPVKuSW2zuG7G9dAZLi/gE+VwtdENv9wvi1
QI7s/pn95kx0wZ1o2aOq5tiVgrCZDQgMlZs6N69Til48nPeSSPf7zoqVEUy/8dhE
a1t4jwlUAMHc0B8i0pxiSRk7fwy0hgUVDyc2SrTZS9BVGPZqjb9etirsp1nDS+p3
y9WuOp5q+uAI4Lf8bRsbEasj8RBUQtEyWxoFOAhHdDMQEFgpSqKiVtXjh8T/3B05
k2tGIRtrLiKeSGJhClrq9lfOWWM7LBexQdOUeHeqXJ+jzBOJN5ur8rcyP8Y0iKJ4
WRjjGbot2KGj+bWLZGa9SZLZFvsDd/TwaYLJqsom0tPUZqqHb4Z7UIGlSFqkI+ko
8ePKTE+iKZoeCens/YuKJC4VsRcamhYrAwBpA6KxLXmgNM1taHX4GDkpxBwz8Ahx
8S/pFT1GGHkaKPj/sCpv/o0WwSukAAR2e8gGDAx/BQht6k6tWB8BC1auyAQMeCt+
hl4O6My51oucIjDMJLNK4ZzY9TcsDy6SU5tWoXmYqd3eqcA0/6bXI875LN6GhUrK
xg1IPDLzDhX19UqW4z+XAADNngG93inOT21v9HvofIUH0EaJCumiUStX9Fq1DTPW
4doME8aSFePWeNl1H4IEuExlq9ZktE4hdIXLKK1WZfB7LcqCW4X2sy9B0pqetw87
zLCJfaPln2awyE1G9ngkryODBCpg4FfFf0mQSyTtP5t5lMtxLZ1U/QNy11/cPHB1
nCj4E0nm8nn7xnJEWUlaaOMOYku0jew+vloM6XeBCGWbxAe5XDR+3Po0x4qNmY66
U1RcB05JWWUCrksJHkdluKaWJV597G+4+8qS5i0DnYhu7fAZ80G6GmkAux0xfyQg
fUqA4xux76J1Ah7VR6uRHIY8bVTc6+5qPfMUVoX8C4WGzWVmNh2Zr5BuRQtzJcHU
E6GcViZ6wQi7/h9b71o4Zspbg6QyOTN8MkDTIMohg5zOuwomVcon1qxLwUIgomkK
F5fWPh/S0s5+Ci9rG6uSsJ1KkbarsD4Ac4iWs6z9AhxGPAuKnBGh+E4SQkPvVTUb
EJ6KB8i/PvUuX4mOHTrzUkcQLijdWy5Nh0XIQa7bjftDE7/mayt5xo/BsRJ2bxKc
dtRhRPMtZOLhqsJFRnNyBR5K/6UJo/FLypln/rbYUEInQyxsfr0LsVuIKwy0snK7
DZTO0DYc4fVp0Ofned3GUfXdmjk70isFDP2DM1HOZlN6a22rc52zKJpOHEskffpb
pqH/8/gnTlSfvQT8pEybEJoxG3SHtEwm+wnDKAz3XVqgxKFdqTG5IlrLI1p5aFVz
xCvdnQUz5v20zT7ImkJlv/+F/ydiQi7euwdZWEc6IUYYO2t26TVgf1+/KR+xy4f4
ePPVrjqtakxN4CThyRSBwAIjzXOvoW3z9OlJGMP6bsAKKVS3OQkwhdFxNUewursD
DU9ZAD200FCJWDT8A4cWe1mMO/UxjDGzfue7XeZFb5rKRiJqhINh5PUcO9dhmqZo
w8HEgq0AyDb4/p9ZdaV4eP8WwjCEL/F/lB46oXW0axlOT2UhkKBU96UmQqL8FazJ
WcRwRPFMtVwwC3jsPhfpv0MUplgVI+A6qjweMNTu+8prGSA0rBbPltzVk5HabmLQ
mACsdUX7qKvvTjcttJNQnll8+e07O7+iX4Ci05tvq/WFfc19dfU1DzWDLXe6YkZx
kwhiTMjpFNtpPJqnAnrSyWzD2ztBxHGO2A4dGzm+uRUYVdrmKCrFg/kSTAfN8Xtl
JVCxQMR++DUuNSHDQ58e/fTVSRHgFCkTnCYgxwj7E0v+Jbdg/K3/Ha4fy2X3vK3M
7MvzaP2ns1Nq9Q4UpTNMsKriIBpRvUHrSzHSRnQ9M3BbCTPbQDtafeDT2U9/aCs0
q6kHjVf08exNVu4ugI10KBvGBQqVeC7+sk/R8f0MyyU60YNxTBwd0Kx3LJoi8WuM
z//g6FVS9/EDrv9RJ2UQi2Vnz+jnnb+5pjunTCRxngKjj72rv/gWeCiWDzWhZ3Wb
PdacuLIyTuW7vsUpRmK/gFhg65TLL0d6fqZI0iPq7APcU4I2YRZT0q7qXmAySt6d
tVIm7Q8YE9MDQxz1eNerayKzYSarmmbmTrO+bDCtCa/ST82lEpmT1JyBxl/7TKMG
tlIhNL8Pzw38DqMg84uIXLZUJM9OKroRUqakmY2wIaIPjJljrTwCG3O3Jc3tBh34
8D9aQ7SNBuFu8HTAbpFWHm3OHeSwbT+Tuk103pT/PTVwn64d5PwfqVtKgH+1X9yB
lfHBWYcuQmCSjhArVQQ85A0+T4iq117+1ANy49AKb7L7GtqWz4DRKIlcYH97C96K
jglP+KrqYF1T9APvkZrnc5FkGDqafFeHDEvUxmlpZTqvGgnXErQej2EptJnqm7bT
/ru408FiWk0SG+39U1MSJEI0LGgOYyl47nAk8g+pOdFWn3ILJOKRThFTVFtt0n4P
h7JBwI/C4unOw1qnM3GcOnZZfFU1toqXUKRNjsTuBVMoxOxZ9bgPhxSadSeIKzlE
TDSw95PMtMu3tTVNm/eYmDE7qyCzbGSJlr8eAuZ2doLYEoRdrcsjco/bnF/zcUcD
67QQHemzqS5bZBtJ4MROOd/mmvVftoqn8CR0PwyyhWOA2bBqTPSgML4CYa6y9h7S
CbDn1ZH65JybzaEuYPObMh4t7U+GeASLIW8FfUinVFPQa43NR1BULri6FICKqlUe
ggbjBpoyutGtFmPfQJ73NuUXNJuDpwLYoCqgMbvXtUKXBREHrNmaibN/zW1LRjcZ
n5MfbDKCiAEaKOfz465ecqgw3IMhR20FoMDJMbJr79O10zoUbr4pGChUns73Z4Im
sMP8+Faq6qlhZKvk5mRtRnEAThGrv2HRa4tRRnobQjCMGOXIj7ngEl/Mv3B/j9JF
iy7Qgao+n3KWRaQRtQ1AjcgoamF3RoYT3TAzRV8QswgavbPQEto0vzH5vQmp+FGI
4O+C0rVN17Wvq6gzofGEdsE4pwun8KZf9BumHimxQJJNQx3jBHuKWhknClflWXyT
bOopBm5OPUp/j61yigO2bQwhYXVe0sDmJOtWuZdeO2bWaFeHpUASL0UVYe1Bz06G
bqbzNxssdwyalYACJJidHEkfUjLQIQdnMg75KxWVvAdFbd1IPC1Zxd0U6GyueR5r
XZqxM9d7v98QXlMC8kn2zlxbBqc9e6P2TuU/ra1cRGSQirkavaixHJTrZwmaKQDQ
ULaLBRGuQ62azxXQOYsomA8MeUhJM3PXYVjj5CQQk3AZZ4ME+yzE9Ye6mQMoYO5O
4n+820GWUFKw7LK9kGkZUKXkEcrfBwMPiYz2bw80CYHH/7FjtYkguQyeNUQ37z2C
4Bd6ZRcVRM8bEhH7YvlCCV3XmLWPPXic+fqRaq+XYJc41saBEmOlGtusg3z1gyuE
Eo6EXPvRi+jIqQbuc903oPH9CJ48XtsFwiiA++z6yyCDHqZ8yHo5bCRyUOdGJtIH
iil3NLJLuGjJRQffOa4SIS/q1cZlaS6GuFpLB/OR9aaLx+N3NZpnn6fHAuSeiA0S
lfmFP7wJ/wH/QIxsemB1GBT01/DdpCcIWFuuNz9E/IXSclav1tzJ+KES4/7TwzPm
fkSHn/c1UFn9p/xq9U27vf3Tb/gOu/lu1yM0LXzPgKwTckp5Hxxlx6ufmIYWOlya
xzj/P8xL01W/CfawgfBpo4sUFlUxvx9OVBXpEexXDBi5CTsAl8fpfL4eaWZZaKRp
F5Ql4N6AAaOJdupL+LWR3VSrXWnqZTyN68kUXMsbL6PnW1XZxIGI83u5my1SNXhX
a0zZCH+bsi7dz81xa3O780vFn9YPh5AY0UxxC8nWI4twpUEJ9RxDXIy3lkX42T/q
gb2g4EA5QF+UCvF5xVSgmOe9yzERHkgfl5DlS5Zh6qHeCaWBTgTkpn5umEUCDwoG
MlFRPITqSB+j3/3uyxVhSK/MHMY5Ap+mrZQgDskj2pPBNBv541M6tw/s3UUFGnOF
fRt5b4qbq6yqxdLd7NVN+g8mKPsQCgrMO4/NNXwBcFEsJl8wcP9cEAaN3aFWor3B
yuuyeYWmtCTCM4s+C7r1L1/3r7xrIfiH1/QHqSczOwn3M3v8sdU5nqNDO4yQrFY3
R2jfOLpUE8MIibW4L9k0eoyz+V9JAyOwLKrsQXGfQ+GMlYtUDgn9vB32jUbtVQ8m
ZB7D3dw3D2Wzo9hnIUMG8N0Bd2D3nZN9cB1cUALZGLqCCyduIbDy8hD1pGNaNCyu
vDTzIxTOLz/EERS2oBEW3Qx2SI0mbi5AJ5GiRZEx2Bp8pKmkoYKwqgbErhhoEGHa
ROxptJPQ8mppHK+70NREWv3BDbdMStLtOJo/E6o9x4D1odxuT4c7Of4nI0gwXKVr
qV1XkOexi+Kfp2vuQgu78TASeQGFtwSDHVjaY5F+4UBNw65b4d+7rKtAn51CCk39
wz0lQScxldgOEKhNf7ppP/4cLiq/6DzuZXbz910A2x1v7Jo1gXlysKg6YIaldEZG
5F3r9SCIpIHxnOiN4O+Q9vl1IW0pZzrPoe9ORM73+UZl0RGERWpGlQhIY/i0bB6j
JhyDiE7kjGKkBvYWFRT4Zeaw86DH3Mqo+ADsTlxD5d4yt1Ispc+rnkYRW6YmOJ3J
s10G8gd6bEZIKLSa4SplrzNh8KO2UOnHQJj3oWJeeF6mpu23OsL5YERal321jngn
13zka3YPJOtUgA/pZGC6+SuvDbpF4Ol9HxJivIckLnG7e8mlmaiJfRrgHPprXvc9
Y0fVMTDaZfmwX2gNYsCfIdvd+1FgaI18vRjjJ/9VWoVOEeQdPmYuj9Z67NnTjJaC
6pLr8SQ8YypwKq/cPp2JajxpaZ6DtJGTWAeeZx/4LHKzZfxNTDqD1ePY+Hs5GvCK
t3cgdHTol+3Xtn5ZcNyKal4UJB4JfQh4gAgOS35WJ2R8sRCZ8ecxGfY/FrY73hqu
dDVxPqxAAx9eNWCCvbMn8GdDSwRAChJqlC4yb8TQ9ArdV5lt02bTy2gnBd//I/1L
TX4dhN7Rdgp9uaKO0u54rLDPFaEb8uRwXp+7+u+2hc9BUwB91J4sa+8RVdYCS6uI
C1irMOg92mG5uuWf0LO8lBBogApCpiSbnXHd7NYUeM81SzpYph2Wxr7Tbk8cQ/aJ
cqJN4WF1pYQruzneRYaIVPIRAaruPCXX7Z9iWTpCQWQlVIW2X2icbitVfAeq1HAQ
1Ir5y3Y0Se6T5yK7sfhPfE6D5HrFfgmPPFxvfuOArb9cAR6A1PBLFSdAYaATtiCX
HxYcDniRsNGDQA3RG9GJ66Xc0k7V3jtotbZr9lIqNJeqLjuNQQXdHtfm4r6h+ul3
1I4fYSiVxu8BU59JYOFvYaNJSwF4icDIKyvII1bdpeBk9gedCqeWjDj8MBjOEFe5
aHPiviX6wTDCK24P4qaBGb9K59CNcH8fyNhApVBJl3vJrr6f4gvxfiInh+S3EWOb
QYEvbHg77N1vQ6jcr5VRbF1H2dDrMcQHs4gDY6ExJhO+At3H7ZdQRrewEdKrIle4
HHIV41HtMeHn42vKt4UrJIsTcnuzNJuv+q1k4eK2Thy58JIJ8MpyiHJ4mIJ5FK3o
cxaq9L8iQCrc/qc+8e12VZ5QiROvnRnTb+eng3QWQwts1mCBM+GX3dlV0TJfd1KE
PlFAGc1/vLvZ9v5oy1hCfUp/nnDnG2mgkuL8CKhP4OcPNfyjE+WZMzRicjPdi5nm
m0sEa0VyCs0NohgB3UT/mXts/Uh7j9ZXb+hT4HgbHutrTISQqIgNcrvYU3pm+6mT
6YKTurXoDmF20cJd4XjWx9C1i6jgdGMwyN2ltIU3p//o3KbFl0vDw+pUkzg6ScSZ
2tMLXUWGhi1jU8QRsChTlFAafXPKBBdOZTB9Abz/Ey/va2OD2X95USGV323sM4BK
P4p+ZHa0STYtYyeCsHiKIEyR6q5hgNfO14GAL8zba9byaCjzcjKoUKJuFg42lxVR
kwQaRx9x5dbQYRCXqIVFV9FvGWw/EadOTvmF37K80xdmdu8HUogJRlUewzfopRHp
ZYAL0kKYWOtARQH6T7UtlM33hDjmUDLS7ro94N/Mus0jThexHD7kMw+rZri0/1TJ
GRm9dHJgvRBVDuVt/n05aCZgsmSLnecUyC0XWhgCbSHtoDaxmBgnLPzmzmBnz2p/
wFhnQweePfKwacRGepFuw+J/VczAJKkTlIOs+SXY2GstR1wsV4AXH9/ss8YwP3tq
8zM8v6p1g6dOaS/R//cupdYJ0pRJ6VU8f/4EPNXviNNqr1lpTeVgxG0KwtcJykWt
Uqs29CGL8gd3plQaKhWMbjbv3S62LtiLewylr9pqJDn3bUbn6+ytb0LqkOxCcTB8
98kH7almW9p8CQnNzt/9+J7BtnejWey1obVh0f5Lj4SXQklkp/bzizckeGomj6wU
FlRencznbl+20vb0RGwS/7R0M75E1C79yTNpBJTWS99871zveb7Ey+cmIfahDcmd
QQ/bdWSukADwdGrAgj8wAVuRfZPvmFDibaGzN3AkVInF0mZlzwMC/iuo0HK2cKWx
EL9Qz9W0Ox1c49xFMb9ZUs30O8zLUq5TZ4kSYUomQAg8IXeHCz4LYzfEry2Cfy0o
7pB57M5PeAuigqzNwrKJlJR/uEsSg0wco4vrAK7s1D/HgHwmVPyjeiLeME+iePxj
iCA4cEZtnfSkXyplAZllGiCLKwdCzdTGZNoXdNGm6eZ4HdS8sfrg1h0YBM7AIgmc
aSp24fj2gIPQnEGApYqoK76ld5/z1DJ4pQlIm2lXqXCBAntWWAogRvfcjwdICxwZ
5d0LYMHMEXY5496cJm73qT26FIV3eMtS1Am04zJzYRFlee/E2Nx4PrHv3N2ePQP2
x5ITYtAKU7lYaS4tFSI2aT5MD1JZ6XQw+c1ibIKgRf5hCFqsrvDIgR43tBvLdaTe
kGlxlmgpQZszp7HWgY0cgzkG3P6493es50dEhhdWjU2kcTdLeR9rTcTEHkaYClW3
SN1j6PK3Bk+k+S/3BnHm54w0bYllXj86sBuaZUHMS7wS3lp7u0HeQGMioin5DeR7
12utvT9UHGYVu+D1B2pzsBR7qP8gRbx8hz7vcAo86UE2YQpEle3fMCNJm32SilYe
J27ITfoQsjwutNJkcElYK3eAzOS2YOcgNQOyK4iSRm9c7ExTGZ5+iuO0+JAHo5tr
kDt8K0cXdQ670cfD/m/6grYB2e9/zzwOxekK7n5XcEzlHXfEDKLrL8wGGPxspvBQ
JuCDLM6qWVkAUp9pZvSNC1lk/TEnlpvcXd3J8Q9Zjo3X8u6/kA56SHSylk/giqFG
KWswZtYf3QpW7/fMzrhPSdZfG896SHmXbQ1lF5FLGxHNRcnifOeyEqYYdeAuW9BJ
JCVF/gUCJl4PtFHeUIWimbP15Os3NzC9IPmeX06T59vfnaRtrgCvldvEb8Mm73bD
bUXoVAms9ukc3qkzK1kXRw8/SoJKXJVbisEZ3Q2YMTkXBmzrCM97sx1Y8odCEvuK
UVlTolMQhiHKrrOQ9gj7vWShyuPYp5NOneCy09dkLogJo//uzGk9Zo+zU1XbL7et
ATm4K/2mdQPLdW1MmhMWwoYdt+VvxLlWtE+49mMJqr4EBZcr7StF/G7d4uX8WluA
SNqJjPHYBQtwA/EkzemuZw7gzCpFCSrGE70y4oB20qPRemu2x+flu7eSsnCuoiDZ
Cb7qBiSOb2UVptj5bNNZX3jXAQmhxBV8i2CQepIuTWBul9Madqn+lEN0JMGyTleB
ux3N4ob3tIkEaniLtKDDSwTnN6VDzCf9mEuv4XZokkphFlMLF2gEAqWnA2rqH32I
cYpBaK462WOK/FH7K/Fubx1TXBhpNAclr5QyXOOrTveTofVIXJh5IzPR9VP4BKMS
OXVzbdHWAI0YXNYgqdqbBYM+rpuMxvm8hfCvB7F1GkJ4AZlaQ+TnINyfCOT/2m8w
35so4mlo7Z29isTUN1Aa2gXc6NTZt/kDF56rirnkGwHUtGtHsfXtLsX8FiN35NmT
eGMSARrQsdfQ4pXgSteW3/pUdNfnXldEgs0VAe43fK+Bd+/ciZiyjNbOwiHMW/18
HMGrrTIj9ElgUTb+QWeOA1fYt0zjEvh0G6hoRO6kvxYk4kGpMh0ONKdJt3D0TCC4
Mqa+rEj8dDmZg3Xlh7e853D9ySUlUUjIGrFV+Hv+278YynXANpc2loC/EQhqZRuU
T79u9bTXrceWbhU7NmOa063/426/rj5xT+d/cKPaN02GufGUy8wNl0o7E/rrevlV
iDQS97LTgvhIjUuVg3HvsVCOgoeHuUb/5hWi39cOkmMk4y9XuOZAKnV0jK0pwD4G
6qd7fYTQN71U9hL0R3EnVTtnkR0vZx+rQthM66uck5hP1ivN/+HKIgyeCNvFstbD
krhEinYQpMpIRpVL1EYMKt1vUcLj8udfbsOUQuozqi8TMA2L7syJhlGA/ouC05Uz
kh+uMNJOsvtlNUeTPPfQw9JB9WqAUNYmT6QiK7aU1D5SXUAs0wWgPdu+x9x6Ljkk
eFuy2ubbvMf4N+T4Ay5uyJ+zIPztoSnHrYk+e2RIEHZIkYtvZPGAxPIWdyqx34+I
8KTwflKWMEQYXnCbchqXGM4m6iK0DQmOWGxk/MXHhxnO4HLv0iz9qJVBfPXennnq
cf2KlQg7HKWFjGUWfYUWJT0I6CFVNO1DHAnIuplZmUr9LzjWv6lzO1sRDcD87fr7
sKcx1MzpdrwMIzfLIfBOl01SMMFJT1cBntF7umj87G4URZVFyBgTOXbhBl5tI9H4
ZoZC05OFFZGnAtuc+3h3XWs3MOBMGAFB8hIoeHZbcqPOJoWLvvANtSttJeUeOwix
9zJpNgNymoSVfNCYHWCtBuigtaJk4Z84MX57Zn/1lfw2IaVZcnuGs8cYm4TRnWDk
io3Ne4tkgMyZyQcLVJPA8kL0LOxKOWTvWSgZsVAA72j6PgG7YyaLmVQKdJCOi5Ig
V50Y5T1nYP8CoxLJCVta6Wg42VCaAUq8tBoYN9ci5jHWXenIYopLJgcA29f0l7cJ
JK2l0nsz7y4zEQUQ7M33zNlARAWQ24OFy5jHcRuUnWXTrSSHEGoevd22Q2dWBWg1
T268UGq21OItRDjRZJS1R0+WIIkUL+7ls+Ue9NsjYm3gfgcB8wD5GWg3dSkVa+W/
natqIlUV7Ytp/CyqBMEj2HyIT3p6N5TaFvODSP4BOGBmhklvlsjZUg4vkDb6mo7r
rsm960h2bD70gzl2KAlDT4kcec1dlf67CMZoLymD3LtCtRLawbl7zPdeFDkhEQV7
4vZVsxYY2raPPd8kLJcBDfoSjbuVb7i3aF9UKXZSrmIfhRLFsmnuyJYudeo9Lifd
o96AVry6gNVbQmzxnBwmDgV2IVbJYNznE/Zdx7q+sAJr4Brwv7Gaujm/Plk5cw1E
CFWblqXclvRSXepHs4NsIBmvpR8tVchYMIIO84kBq1u4alEQSRkaluOTJXb++/g5
qYQCAKoGFar44idG51k3g7PTS+lqDlXhRlDInJMBAQ56J4UW6OGqG9L4Lb1YF9wR
yp6ZNft8Kmsiu0CZzQ2k/lSKuoO7LxVeaCyAJkjNZCmlq857DMXTfK8i5uozsKbc
/47YZ/SJSc89WBI8KxzsXulvKVFoJV0c/HML5ltZYiPTNwYwnD5NXXdr9B2a80SW
pXRR9Glx1L37ObDUYNiEeSw4gBw1BEqvb3y41QD/gNTtLIAQI5vK/Y1HTlNudfMt
wIfGPZGGpQccKDIr3Mu1t2BcifHA879wY8nADbnKFoR1VC24QEY0OSBCTbXMm4bn
gViS/DoBDHYRQ8660+owiqEMxJ13nzAFinlNOoQJTpdFCSKqui5ToUJCjN2Bmpgo
piAJvVlemZ7Y5s8AXDVsUWGgaI8j1opA5wY8mNeWiG4FgrnUGJ5hAeYFHAbmuxA8
VxTnPySYf4ElibwgWDvORdsqN1OXClidKuFYVBnOXgowWJHigW5f0YGU4tRusoit
stpZ8aZfYb1uLEA+YnICkyasoXIwIj50AyOWpviLll3Gz3c1fRXIQhnVF/PcT0PH
GsvIQf4y742SzYGfCfElL8pXpRRXfEIpEZTGTwz7nXglOjZYlTyhvnuhG+t+gkZL
145c7zunSk9meAIJVkIsLWTXtIa4gzWBN4EWeqWATEKqyn3OUwbUZYLDuH3D3a/T
RksV7XVhR4Cm2To4y7xH5IiGj/EKKqIfROo16aDEtyWfw2HP2SVS+cqrGemcDxQQ
3vTVmClJ/dSryiBsmZ1q8B2RyeqoELNCPuLF3g5DIk+gfZGnAfmfwDXv7RDqwlbU
Khg3dP16ugUSKMfh+QniYYc8VqLJmwDlLndl2c90XpDjZKF4viriUL4pbeqdu4ui
0WpkPzMkXoAZ3+NCsbKZAq+iTNzPHKT7kUXjnHZlOQuQdXmP/6j+7O1aZWXw+jm0
ByZH0bFdoDjNlW5SjBdWmxOwcVCQO4dWnp6W7Qq3lMAGvrs4TEhL6EbzM4xgcGf4
8SvkkyRPL/6m7huc0R0Epa+A4esVVm+3Wtb0PWz0pGceHyth2gupY71gjs/GEPk8
fdHSSeuA9JPEphQcJfNxRX/g4U+dHbeOF9kYu8wxsxbo/g9CRfPkLuJ+8CfU4jGx
ZfrCFenCAjW9oCGCmTLx7rlNUmOerSittidJwnRoOjpJd2h/TWJLvb2VP6srP7YD
KgpTlYgTUZL9X0KnI1NaeDSoKdgot6jTYACAs/OswyKSJWQgbjeE4a5slh83xTiQ
ZL/RQAVEOOpyZqqWzPkzxSEuRKbYL2d8HY3oxsPbw6TpArMB7NW3nv678W6lUV8B
oXlW/Uw/LOdp0j90fhwV/7PPUJrkHQ0JKt9j6uJJGQV7kGBKnbnvhvS729rs3cn4
pdp2yS/v4nWMjajzU8lM6P7z69t8/oXXQnxDNKEPeiTSQVDWf6WZl9BSbwp1NoB/
npMT6yCbpJPk/AtHQA8qSeKxCSz+gQyq87KXaCDpTSmgDdoAprRtdC5PMixQHbOK
DtXW+mAKNS+rw/oUhRItnv3txGjF1DBiQL5kVpWE0esLHldhAbmv8z8Mk9U1VzT7
GpUQBddWHxbfs4MsKTAf11TpEWYu48nw5C2IVA/Z2aKCDOE1Gphfiff6IfMioK5L
YToIZjKJNdTwza1ZzcrdjG15wJ03rrFpY13hDS02xxWKHnOF/uV9Ck2qNJy2VNzZ
GZ+sGJ2jUKRjBaLwOasKvnb6ege82xK0ChZsvywTXTf1hyk5H0jC/fbPWn3Lf3Ny
11rPdscSYXvSxswFv/ZTiNQNddOSNnUpH403cJVLl7WcQjgwsK5+AGiyBFwdJjL2
KlyEiKVsDTlyHM3SnHw2XdHsp1rmXduq9jWOoJHt5lcK1d1RK6H69PhsbVahN+96
7BOWOyNLiX7eBDO+8YhygG2AtxusbtNtjJgg44xxcwoD9jw1QysRM2WcX4lNSMJk
1R75dVu5THkmv8u6g1Bz2i1uvYo6+9+sXiwlqZNaOo8FEv/D+BCE75q3xJySyNv6
+7JWOgJSA4b/Gn25f1/H9AUOV1GSTZSVoBBAmvJiSGVZF5lP6vDU57JNcK7WqsmO
Ug8ztWAnt1jqL7b0og0vQo0Ip/PxcNcL3+w0qWAtDFcR1Jll1fVpQgsPg5ISSsrt
nhbdcw3pkAqae129HeUwxKILZDrts+Ax91sK7pl97UDjL8E0g+sXbm9tmWACvv2H
N3+8bVG3YKfGpx0v/TJg1duUWeVAgNitCYiWEhXddBI+39zB9QKzW9j0X/ZmmigW
IuNDBQHhXiz18cxIwSGneYmWTICDUl5yH0R3ietxr2NiLX2Md2bcjly4D4QypyQf
geJou+hzQh7XZjBdNy0B0x492c4ZZZxH7JTtRCM8Eg7ACLTIp7oNR8ZMYsIVv/ai
b0vSdGA3lGk/nL05K/6aNNdqyhPPmEzCv8PJa7nKtpGFXMjIVu1cC6cGcNnXB3UY
pQTyOBE5sKJ5LRjQ/TuS89aIcU0hZDf26C1IaDZ4CAn+go0CCqBDTxu7qa7gkIwA
gK8J1c0YnIwduLd6MonPAYTx5cAVbHNJx+Jzj2OzeuHdByEsKnU1gdH3IpdM5hzX
tN8Hcg6NEqiPvIq34xogViHDEeNuDCH9Q1nwu8PLS2mFaj7NAPTnikDfyV4tmggL
YJOfnkPc/jenOMX0SLQpt85Zja4pnIO2SergCpPNs1PeQ5P0Dx/RUWqgz5cjzN/x
rd9mBTnlYeMp+YOo29q5tCj+1wR1k+sd5C+PoRtj3DncTevo81A8VoYn0O9nxP//
QATP9kpU1Xmb/ExTjcauVgz6Pl2wdcUr81PjCImqO5QA6n2fX1Uevnb1EP3e8uCc
hViCs886vKRV6m9PLkoc4nrZQfrhvUgkgPtS4SCyIix5y0/ZvujAW9w5rd56HRNI
fLFZ0lEXTiL6qwATFtTsgiWqCThSe8lCY0wk0JgmDFuYQii5vwmnsAPgl5D8kh4n
gOUDPp300Oha76M5JDorSzTWlbSwdEtgaFV1RDKhWbZgfMPqZy0LMqRaeViy4wsL
41VktDSmmbXGht+3YyleFwgvrNzjMTv3o7XVaYVAPc+Gz3h2MZd3Dz2fRa/Y6PzS
OzLxsc44AX2a6Cs4XGJrWlMnI/RW+na6NuyyxWflBDW2jDehu0cos3GrQQK7iAE2
lzRQGU3pAinCw+DRqwMbVdB8Yft/QG/QNwCGwTrrMLfvFxoYUpdxvaj3obf7bGG2
KxVtPcJBxC4mRqzWgBvVj67bX8q8YonRG/3pxwbQApEV4laox0I+PsQA7nUT92Wv
U1g2B5PvPduzVgw6L69QGKGynfBzEcuWYieIclGP3JEKLcrTuBZMoKHP7L7M2z24
jnpZjppXfFaF4G7Vg5XLaS/7+i0ePebZ5Gnf6nwxto2ecc0YoIBBhT16qG0IP/r8
r2crADDKHbUzfi39S5S5lzJYkEmgM+OPH8aEVk7Y8tLeYNtVh/3U6+TafVMq3Ci7
bZFFVIlVfTtepxXkdoWq2+xZeuzvMJelftDCTkun5Ph5WaLiFLBU4uNNZXCAC+rr
NTAkmx066FM+xWYm+tQwqsXnuXqGwxCNhhJ/JF2TT9giLc3uH0qePxJDFPcuxqF2
pnFVxdYJYdLvz5wNv1IeI8Dc8JIMKiXHDGcdD6LVeHCfZXx/6htLw2yFAWylZ4Bl
Wat9dcuQ+CxaMt7qcWMhsJBW47hZC/TNBSdM6p1BtFjFKvRd49O/JFgBurYyEIya
To/gX2SG005He5Nanjf9DHHR5is6pYPFDQzR7Y9I8yibIO68pps9/yv9W/s28o/e
An5WrB2CjoQMsQ2OC8r/A6zNkaeDTN2qT4h/jTecWZu9uFS5NPGS4tKpnIkd4Obt
zRM6luizbLQJWBumFZldirInKaE5xU0UEdjGJos9F8RKumQoAOjZCQ7W/erhd2Gq
jyAANI9pEdJh6cqLABBHFA7PiPBkA0Q9bM3XOvoJHFmzKFFstcH/6MBQM7kyvLxb
SIjmmnzWA+8Oy0SPYA17Z/BI1BZoNyayrAs+FNFWoDrvZ4gpGLnWuIkQEAo/+rF9
J5tEwnt2MeRZ/DweNlKBmjm5aom2ods4jtg8HZLN63YiEy1Q0+Cbj890FZdg1iIO
lNqsoF/aefT+LH49Dat4cgQNIvQf7/kumLP/HdOR6CYAcvvAh8llfMw/nCEYltW3
5NKotQ2S/rmvqBvRwExP9jkOPf885leaxKDro1saSwuC4OXIZmf4OFmJUmeMregZ
poTZwysLiG8ScDrGqJRhoUCXvY8ILU2mMc5xOtCSPZxR5Ln4bYoiG1rH5SDThn7s
HtYzexv14eyQJaGBJbDzT7z59IPMsUIm1TCQRYeDKzy3lnzATHSe8JkgwOGCJZ1v
juhZnPmctp/2XrVugfEcbjNazgF512jpKfMAVMgQUYjA+JCD1xc5EFHAS1W/03r1
XnHWLYo5Rvy5gwtCtHOZiEgYDLM/xNGEAW1q2WkN9bNQ6chtQ9OGOek1ia5kEZO8
C7gDnJqY323TKtbsp8umvONOggsBhemOQfK14MQj5GuixLXgUbb8MZGTHkbitH/v
r21Dubch5lTrhN7XBAEjeMhSJyvSJWu/4YteTP3ZNtBPuEpGVmEn63HBf9Z79DD4
R1wuUcggdS8FHKRDU+gbkWNxZw/rCkyHOXw/njOALd0W/7WRRcjgr2Vb66nSNxpi
P4/1NnJ/To8XdHH3GuUj+QO7gr0qtjlVixE9M1x2Q0uU3iJoHzCNScWyyHTRqSoM
l95PrtycLjK6zgcwpi5/x8toRs/NbtjdEwgSZKRmlPtxwsUfJwtz1D1fiBwuS3rm
CpvQ4UM1v7tADmINZ6EzRQXDN8iHULfb5GzHNCVtbhAPoPmp+XDm9tXD4Cqx9A1M
TVS0WGiYbl8WATmvdHB9bjqICK4X566sXlVjVkg/7i/tJo0xWDsj7cszRGS1InH3
6I/+O/pHjvvK6tCQQUsi04oehcRMBJIvQAEq7DcbGfWuLTmjpX9597I/opwTvncx
yu5zF+v6VKE6djHZnTi2tg4P6auaKBRl82dDBT3ONATgSe4+XVnf26NanRsGwpbe
fJmf4XUrNzI79Ofek5lvWBBWfB/O9Pptte41AZS6i5D+8x63IkIHCPX2cVPikxsX
xIU15lhFzl6HA2L2a44ibF/q7alGJWU/NH4zl8iMUvU1sqyMhaC6SPoI1ZfPwcQO
cMlk7f6IHYCa47jFWxsyCeGnXUf4Q3WGb3EHhNVohB7yr9K3Kbx78ESv2d8ZNdq3
ssFood0WwWSRu59U3GeBF1Ixexn0tgTpumiykgJ3dQ+iPirCXEQXHW68siyEyyrF
md970x8hZRghGYncUdv10GO9XhX+ZPwTiyGNEUhlLY8DNUDnKFJfD7r2oLC8unmY
Eot8fjGP7ZxsIwtapIBihPj6gf+JbcAfdnxz15tPGcydVU3g9vTc2ekn67d8lHCC
4mUQcx6l3tTqTbQF6JCW7GfAY1Hhaa719YCtnlc26ZHxgZBRGm+ddvnZp501zDwe
wus/0oFlzPuDA95vXMq9j2px0l1Q+YNhYf6AZhJcxdPl9jYCOGwx4ZA3emRpXgqh
r6AzH3dKigR8HQUlfazC/tIyo+h7plBizkLbNU3hEF0GBChifDkwL3/6NtMPXylA
dJOHFRORxZLNeNLy71H1Ura3+EWm8fLQmqg3ZRSMhDt8nWzfBzE0CvqxtrU4parW
7BpHJd/7CkW0is7/RGLMufnGbmlGw+hr4zMv+loGUs4Tyx05GGYix7dXMjlxExCT
kFLBRUt43lldNAgJLqXEqlFzFSJqQfTmdL5jWGz5qhD2IQujWmynNv5rez50PMTb
Ozboin3geabBspX9H0xJIGnmtpQ5hUFP/RRoFyDvNUiW6XY17Wb9J+XtnVHpzK/O
DpRYPbe9Z4/WibDObyFesdBdLxnrKkJ6VD8IpPNEig1OUEtjQ2EDucPaQV2tBzUG
SGj+Yx7EPAlijFbnT5TDzRoklZ3tJhi62gYiiaRS78zAt/Ts8y5euHQ75PwoimQc
NbbAjLxHHhCR+hp02u0PXJ+GdfXXXbeJ78wYNjiz1XErQTpyu+GfvPhdrPQLCm9M
jikOGnuNPFqDvk4tkV3f5WCsSNCxKO5YeUcYlaTn0ctrUEhXyPsAcq8tRj6xeWa/
GU6fAw6EEaKCmxL8N8XF84l2Qj1/niN/God8op51xEnnmj4qall1HfhYwkZN6B2z
mNUS9tTwR1hEr+PgWtNhX5KBldcD9FznXiDOkuLrPM4WBTrDGIKAVPj902I9hOFA
ieMZ/Ht4WW3Yp3ivh2cfkNGx/mlw2AMkoB8tnXUYtzPI8VciV/VcE9e/wt41+L+l
NV6F4TnJUgiw7PWOXyH8XjpAqyyACEhjlUGWZBgOCLm6JPtF3b/C8LxJgeI8vCia
lUtT45C18VAwVcTbBsWB/QJARP1+eKdoeFlaBKC9+dexgxh6PO1fJMRSCpNYi6L8
W0FxWhKNVmCt9qzzgbapmUDt4MkOBhliYIkPpHg6wKGeh9wgIhR2WhFpNcZLDpnJ
jjwQjgM+qxoJQUSdeoP+2nu3QIYbhgO5WA94yISQbQpiBF7DBuIIPryW1IW0ky7g
BllaYdoCY62wnI3YBXYk/wWe3QoWoCrYEjX2/REssijcWJaITUqg6RQi0UKvWhPS
YTn0AKnOV4Hc/uZ+4H2T2qqkZRrR9Heo7BiefVTTb6VdXXkOngI8VaNsDkdr/qKe
MKbMFWnuoKwpOsKgJ6VrTJ215bw7j59HjPmjyBibznqAt75jposH03Y7u+Q4Xlea
Rbu/E/dnR5ZryzO4fBYNMFBNdS7kIc4jU4Eli+eObWvy2FFV8hRyh2LWYHH2LUgJ
0bB02ijLYXp6o37BySotsXd9DEcuNxSEkUs6EYLIhSFFY947lC+lcIME/tVO5cEt
c2WMa8SmTHm6Z9gDslw73c8j+uJCSSX7m7Rnc7xpxCIy14DKDrf5E10e+sfTTruE
iqFRpUHp7hdr5mXHbcRe9v8R4sLc7EyuYHq9ooDjK5YvOpqbAphcbeBs/Y9piYRv
NCDLTiMStrPyC3TA0zNqN6P+op6hmTICLAs6UgtDBBw1rXFAeqsOcNAQhzkwJxLJ
mqUt34oCxeF27BFH1BKSzEngcwHQPKlGWMp6AjUjvGwHrGJUrAzNv+5K/sKEJo8q
z1QFx8eN1ULSTEvFhPBgWcFCNn2XUB9/2JlSeAcVfLZVk1K9wO6njt80/ylQTllW
gQzi+dvQ/4gP9Dw6liyx7aNh8vy3WoT1ehALfT0GgVkcaVVYINuOAlUhVz/VZ4Y4
byEdf2tkr2iA4FPFpNr29PYl89gYlY3G4trbUb6DW36cmvXlFEEOjAYJ8fbioSPc
vSeBaE9J5WoV7d3+PGzH47HfUMZJZZ1QhUV+SNUDoMHyYAG7kPDaPL4T4xdn6blq
+37tjMLRQ8CCrTqrCxxUscMr/bJgRob+pZJWdsY6iZ9ceYW/+1Zt2oif64B/VEIn
6vDPxXpPpqFhwzNQjUzt7c+HBntEJay//wafCdgG8x5PsgmPO0skWubhjeyAnUmU
O9HgtVYKHQuXUcfRCZzuXGx8G9x+HtztTXvsEOWvmf1JUGqAFIdRHAKUUfFSUFZC
AQF7tfHCY3vLGvSi75w121OnWM/2rj4jgpYNZu+Mw9zOnDTqPYA/GFIw+OILy+BY
7hNTqrC+mjBxEhX2eCFo7/hbhgJnmtJHu9OtqbQR/pAF+RdK9YSLroar0B3mKTcF
ryE/9yPskYjOwYfZJ1H7FPd2om5gzsRo6xIaIX3vYIM3jHo1Rgog6FhHKU/5l5Zp
BY3aU7MoR43yeO3NS3NzXG6myD+DkI/cbOdxKx3/QhN8sYwrzshIIapRN1mtWS/f
ZyKYJ7mp+bbrFV6d6ehkNqV45v1CPd6UniaNKhnpzw2Sl8ABhO+Sb5cvFkVe1Ejs
Aghd09Z15Il6N4P+0yF0bYXvFuLpXSkHr8q04XDA3izoXx2/Surbk6PTV36TfRwj
VTShioY9hZQZV40s6rmEc18O7Hn+yx7TDG/lO4paFma+A0QXzAtAXG6hzr6Cy9LE
30mCrZwuNdxce1nlxRQl2fXra30JqQ5ed6VQ9NuLpvZgQMjOZ3Pq4MeQwuYCUrZr
kGbi7bR3Pl4q2m7+gPkUMz2RoM7CbIrUnMz8V6SRq05xi9YJpB+xdJEkwXzDxKdE
XmLT/7c/z6r0z0p4sUfEV+q52GDRlu0SYf801h09SmDOzpmA4/SqLxDPWgR7oI2H
fjvf2v19AxJzYD5Ffgz8VfOZdC6NIZJ9doRoPk1Lk/O2vyKllwTeS861TeGIvY5q
EhRllB8iEwmUJ/URTjww8UCyWl/phuOTtkeBMu+nzlewd1IjEcOqm2bLnzHHOnyq
JFNiFB4NWty5k4fYCXaEfcj+P65LpIfmKfWEqVZ63jBHnQCrwUpFg4PaYdQZv9gV
fAjazpecgxgaZhGvLrlaJbWplKqoqjYvkRZiANB1Tt8ktvh4aSLoZk6MwU5jbviR
TM4oVqR4GOvFUpWUAQfQ7nanCp2lDng3UoIh5NRzEHHPZmufeuTTQsHD3JTixYny
sYtH6ZcVjaSkIKFlHiS9sLC+s0Ekq21W+onpzK3jbGFBeuQhy1ddWLacbCOzCbsk
V/wgPUCPwqu44YraUeZ5pw2Zn4gk72kVS3WgiwRvxa02YRl4gEwZ384Smz5h/41H
FlfSNP3CrmBCamkeBxJUC+U3GNZtWfNWVAiNnNww3lwSu4t1+RTdrc2NIAQWfqqL
x0iIgws226jsTHBGYc/rTvqbMsx2/RSxfx+/Y7gPCDEu6cxpcbfCES6N6IW5PXng
mUNDyW04NHR/5mfLmnlWGT+8PTU5gx8iET1qDbw3wThtuZ+I8jqOzsPBkev6JzBS
k5bRkK39rP1pL4P0u7i9n1YsGA2UEpi1P87uKrJBc3LBzDVhNlCzeSBE5SPy1xbb
ByMecthCxgJBZ6LcrEFvZwCBTD7apVnYPBCj9HompDFVPpj2Qjl43KV7Y37LZdnN
GchQeKv9rxPPihTF1dq/FLQ8YV+RZCNUa7YS4X0kF4ebrYjJQ/IfOXw6Hp77mmE0
s3HfRuFNOdlGmMs4VX2y9Pgx8XiXUXuw6ikEvrp8jX0nZGaQDXPuEf/E5xr7Wu/i
ksb9bVv9+oMUmKby4JRGnYuN4CnS5IRJsvJGm+MGlWaFiylGxEnRDEbEfa0rKA0R
iH7O2gT0mspK7tZaPESUrrZQFyAwhcIV+jzyfKmbSFythh6IBFV/ARr99sVCinGc
XPGI8D0kTQNfMt/YPZEVm8sNuzKvHuA6MBLVPSylGSEyENFSFxSr9LyMWn6sa0tF
VxxaK4hNRDnDS8Za+rIMGR46nBGOak9V+0iYt/QZvYD8TR3KC/ow7PGcD04bMqZt
xRi4bKyjhXzkoRMVzE26v8ieBW+kWpbHfq+TMlx88ypAyH9ba8BnKNeMVHGwxB5q
vOknt0a0Epbse6xkdKAa8RQT/ekNAVhn6p2lPosIRtScJew37BQzP06nNMPZiKH9
W1T/UBIa79FqFWthfdOvOaK8v1hVCsnMjisQ4LoenEmM49ei6xp3ZhenkVZTCwHk
j1n1Z3VS+7Bdzl20FAwjSVneaP5YS1lGV4GTpxNOmcdCI37x25LZOCGM0avtPi7U
pd8SJUpD8TKMu3Z/GFcYmWNwoEXfjfdYfWf0Hhek7mzsdUmVT79zcvW7p2y1cT4z
ztx+53uiHigyoSY/SOvt+LRTDTDrUeBDker7atyIkRmgiym5EkGMjDGTjVl3xh1S
hizTHsbW6hRl2zP2hEvdr4D5GMjn39sGe/faykFZYBETx+T5JU1AXgpHLk5U0QK3
cf5YbrJcqbGwtGJuwd0WRmQJNF+YhmR/2C5pffGaboeDb9pGMnU0cZMgSLat3YCu
xdwCe/L6riTxaI4sTy3q/rNm+hnN3t/kobpmhmFY/nfrOX3ZRhXG+USzvSq28Lrv
1M0G9d+G5zA6T52iO2cd1ck0bAL5jnbSnVClSe6PbzZVCgdE0xO/WRuDKhcpYb4L
k5a2gRM3PhwF4gG3B5N8FHICsnsBxr1+TvWZI2VhFx6ELCNUZ7K31Rimv+OH9k6g
5B0LQUrP9aSoLvI5CKM5nrCSv5byVuhvV55L7LUx0+UAmu+CeS+CNmsqKyXpZpCx
/Aq/k22NZah+u8VnEs33wexTuCX8gVXY6v8q+kLEYG5/MOY9yFdm52EJnEP4VopY
AwjFjpz1yHRxSSNgPoWKAWnOMg1gynFoshOZLLpC+fsTgy4yA6xe/SI1nfO/UxEL
0+coPI8wOJymsbv58/ip+qendYM45S/6t0Uy6U2G3RoXqkchKalWrQ9ywhRhESvh
WIGoHQgm0+FUUBY1K1Qhn2gLPUHvmDt0qczuiZfGOupg6T+ciIXc+g7IaEYyPC5i
4k2TkzvN4UQdCO8Qb8C2srHTsgOyX/n77M3pGOjc+OL24W1PA9viUSlFjhfHxAW/
IgcjU3v3lWXLkZ98a34puCpgV7jRjmY3o3Z4bjCVK4I6VG9ut0keh4tRb2qRytpG
pKpd9N1xzusMCdZkHEAYZefIUBLSAzprP5NVDH0bjXbp/G2x+V0hxo9aYkKWgm6R
Mr+d1LjwYuD/SY950GdzcJMuJ1V4GUcyzUj36Hce4gUNief2mhCIK6nvnMT5Wk+J
lNAJKHPdhKHVWUprxkD2gQVXT1nRW43Xv7D3pz25QjDExaYOIyuWF5JZMYjtPPyX
uv/B+VRf/x8hgQu3s0U1J2IghFstGd64qijUwaSE/KBvU4pJG+1OmL6ZpbtO8ncy
ebM9QkkwvquUxOHDjzHMY0SXu48Khfg/Pb/60fkRXhdY09/SqpTSLCxTIbh0/7aI
JBivoE1Trz6sPbSD4xqjd2YiImGyBdg9vALCE9JmjGpQQ8CP5okp4oxOaxXbaobm
7IFKf+ffEWG8sKnpo5VBEnanE6aKrv2FdcOJ1jyyv4fgD6iIuPYnMzVfEczsOGs1
n1ftcsEEPkJlo8/gJWbGmNL69KB7vuqtryb4HgUFOZjB4nj0hVoxPoTy8P42exSO
xdYjQ3gRbuiybeekB6HLwcnPRn9s2tfONaCMdgXyOc+9KXldvBzk4nhn89ANgCrW
9FWgpX8qkfB6tjyDXz2sdRdlcRkruPbeuRNngpMPAVRzUO+VJ6AYTsTT4SquLNNb
ZWA2tbEc65+m+tIs+N6uW7hfeHaTYa6ui3ybUjIdmH5MbQWlj4t7eJLKnP1DU+Bt
1emVNQFT+PH3c3vtg6WaQ99a5vD9NQFfSndYgiDgptGMcst/++I4r/QaWyxMs6WI
a+kn3reXqw1d9EvarIKkI906Qu1tezdoMDp/aefLUu9pHl33KvR31bgPZ3XE5gZE
BUusMh1fZnwA7OUh6Z6exHfFVzJmnqT4E3aYhxg3AuzaFd3pV9Blro58M0YJIiiy
d/su19siClSsPftzWRdH4FLl/eULW/bDdWOHRKbZwbXd48JG4KDDCJPnmIrU5C2e
e5CpPwmF2Q9Mt+F2exv79oTZKUaIxWpH3nYBPmn6QnZczCkq9nIYtblaHsl8gO5D
YOd7ooMWTBX4EvT8HMDkvcCMTRgaMj4JBnK38Eqx/HgjslfcQmldRmsPcZiEBPvb
JYY2+AFz7+gbBqhBPb0SsCqVh60rrkZ35BplE9h6QpfxMh4Q6tpZn2HFHn1j0WkI
m36keHxrY7I5gtX3tuWxKlHQuxySYo8qsQg21EopHhD2WKt0iz8c7x+a+ALRcKX4
pPrik55Im1DRH4VjBr0ahd/+oiq7gexlPDlKlivo/HiJlpdKQmhlIHFqrkMJB2qx
sWw+5aezX28g8+7XOWXOW0RyDnZp8xpemFmGzseu8DNSl5eZlL6fHroLDqNhbPfg
pX8DiW5F8KmbzhHT5Q4ypLFH9SIs9GJQbQ182gs3NOUEsmxPTIlbJcXZWmMXh0OV
DVhi/6VxjK0oK13JHcSF3PaynwbtJ0di7UxGxmuBYL2P1nWYsz+xrcC0C/j7ttIs
DGzdPEN21J4oDzJ8Jbc0IJRrNIpypoM6MkMpk5BqrK7ETmDceEi6DHovE7ultKQp
9MgtApo3PgwfpcYY1GAHOPZkPiNPvKVvrv9gHJDRlkcc0gLom8FKDPWyct/3UIDp
+3KlbJJShvbP7CvpzsgYu8zaeIQbNjMdbR8njKsT+M/bQWETQrTDqPvxDNWszSSa
c/b/TaVXlzaar6TsQoHe+xRdvxlqlZSzRBUh/aq9Jm+y2U8bXlHUgiSEdI7O9ySQ
5PLVawLNxMcZPByQdi79BqbltUzR3LmnomU01vs1ksRIo2hXHDPe8b6ZrwrWOrRN
E+NmZPLXEzSsrJ4TOmya3OeSQwUne3E0wCgUHyUdxwyGzSwynrghLw7JxHYqd4oJ
nBimE3E1SpckxxgBDxYKP/HlhXeXXXesCnJww/P9dFuOOEa23+tMp/1visJ6ERZA
x1CR6xGDZ0Vi1uj/LR6V0ubzNoEL+cVj8lgwyOtrishUMIQpHAu6EflEWY+w4PD6
25Px4C3zB6PfXuEo/dl26taPhyM3/BN1eOoUV+AJy6qFM4thCcpjA+IESDoJb+Hd
uAVEYfrwro/O9nLx49XR3aRe3DCF4Q0i+f7rOTPexv+EUN8Ij8x+ZEAcGRwQ8/CF
mHqEKtDxyvNs9aEqhvOfLLoAE+1LZMPX7vgY31Lk9oNFn5ZUTHj0Nubdl0VydxLy
yc4Do8gMzwy1n2ZZc6CzhFYvbz4pITzbiP1FDCafZrNgeP/BQ91cxPqu0f6BBXAv
YQrBqF3X+f3EMLgCuYOH2POHq8WEUMzR6aa9ndchOgv7511p2TaQITG8vYBzwAEj
xw5Qelc04C1LtK6GxrKT94+eeeO5hT1RiQltqneHBW/8cjQ9ddLYuyr1fiXOgw0N
atUuOih1SY0r9EEkCDAErTWDGo87PhJCUC7AZf9TxN1Drl7Ly0M0on+6G4L2t1hz
6F/jKrE+j28bwL2BLGVRlXhnz5DmvEP5zp5Ql1qMHaJSOdjbg1tcJXrOvX2IYLra
8lwrxYZc+zlsiOI6i9z+W272xADTKevuFIsmKi8t4zaIVseacLeuxAZ5MFYqjo0+
R0gIp5/Vd4C59+ajbYed8crI9QTeVYarPaPJQzsgEd7pB3ZvM6mkoWR4Uq5/+gFe
2mXOsWeT21itvCxwj0l2vvwBQ8Q/2/gWp18uuD+vstrDPsmOBcL2ZjLz70NdeAIr
bLp19DcuoLu5Yui5uvXAFY7AbY1/NaVA9GvFgb4KvveYTcPnzMbSKVdr6dzqd2Xq
WDzp1L2V+W4A1g57kofU72qwlP6ilh8pQvLH41OFzSsxr3AnfeWcx0NnN6Al+h5C
f+5F3XT4R3GFVQVPrLVkGYkgQ1H+aZfWrkZgqGJZOdHmWo8TcliGMrqet1Y2SJxd
lncfrTuN2XCJOOOFvfr9ZySLOBtdtiCEIlGizj9heHlKsBIi1Xh7U9g08UBQc9Ij
fJ3Vd5ALSKK8SQaCfMyvSwgXGoZSnQ6guFvvTFVuetO1zuNILtti3bQ6WVYLgfrO
jTrXPLTISvugTgLV7qZBfgf/XpeHs21ZWS4lw34sN6HZru6sMSTQR3opILNW8ZnU
4xkdne6k3fTPCLrJuOiVynB18Q3ZFELj3iO4Wu5+sex6oKVrBgV9xamCSP/Kvb0w
y+N3ofKJBYCh/GzrA+610l7/wc4Owvz/SkUr3mfSDZzni6QxPxhrDFr9fP0EXc7m
lSTGsTALfwqt14400QuhjBUu3wnIm9F4VtNRaWLe4uL1koDAYBUKXmFPyqdL+4Eh
trzHj6reNS9tzdBpWyEEs8haJ/RgInau+uPv3uqqwDo+aHWJhnG4lKHoiwVd6EUx
aJk2wA2xRvRMmvnQy1As+gdlMna4fWKOpuBhGzBnIB0rCCBlcSzK9S8ncQw4wLop
UI2hOGCGblwMZhl55SSPckd0lnngOq3yZTSriRGsx1UOy2mDCspkL2QkpGPMzrC1
yuzQfDQEI3XsQsDsgXZqL2waMoEef246pTU2HFjAcWJdaVo9u7EHp6zhpEtPYcxy
c1au4N997r/yOg8FlWHjKW5OSqgW5OgGlTABbeTZHiWlFbK/fLy0mz+KqQcASWDS
LbozAyAojsuMTTf04VvJ3YwBh2pV/FusmNai7j/7NFXA8H/Rk6YvvVnD57Qr3Vpo
fthCZRfkeF10hCkNs166RNRvC2vuw2I9zZNY6QRCe0M6NIiH21G8Ts6nsks3OF/m
Dh/xxQHdOhmKYkUpwcEEvNwVESoRv3ZHFZQthc7hcVaYx7LNxudEXvz5o5B5nyO2
bajF6YktXt4z36cCdrsVSu/ujgAto4TNNtcJ32rEyJ5wA3M7j66w+ff+7lu6UsPq
N2/RaiFk6+H6wQuouYDtbmhLu6dNBB0c5mNZC1p9r58PpXeOA7f5yzbwxS/Jhdo2
oqWjzAFz5RuNQRLekkAdsCVfTmOfoBKJPTa4N1AN3E9CHFp3ObJbHluIptmQMr5t
YA89+GeGKxYKnVcs0tLovUQupilNfcT8iYy1FPuyV3wYyQ9tdS8/QOTK1+fN/wSC
Lolvdhfea4tLFjWv7fbSBwHf/HA596yYO4oNLT6oRaeD10d/DCVi4DNf02S+M3jB
7hZhrFit6auK+DTjTA31uwh6GMjAuDDNEK5FLczWIuUO4TBtXgjy7ZCa5Ap1ZtW5
WzDJYg7I1AF/BJp7+Mb0H0c/WDTaapCEn0Cz3dw59EO6RrfNjwPx2d9Rr1SR9qC+
L/wq05yIdyxfwaUKgtQklEMJYJ0ErimCWhNdDYyOSCVDu0UxfxWXrAJJ5lABgDKi
oQdMrsJvE+q3IK+1T+ooYfrVmREAzAEyGaZ5wq9Ti0Ww/cNVeNjOBRQFDzW5aZAR
XYrCRCqwOylOzIG1BeQhYaNWRI74eb0kfvikiiCGabZjB9H3MXw73BabgoraSYyx
MkrrRB/TtCPpJXAH22LYxKa7FXzTYZKhgt/2iRMam4N9gAgrVnq3b9iqjiEaa4d0
by7Hfe0kRZEkBL038zLPlohpSy4uZrtgAQhW+W+cmVgbD2vUysilRTip9xuXHyy7
4MURslOxq7eWliKoeUN233w5uXhj66dM6gvbsNngD3eZBhRtYV0tHX58sqyYlAfH
c10RU4cnQoChlhjH8bc+utL51/sjzbJ+2oOkdRZaNXLKVSmw4GkLAEHCXcoWIABd
WqegzxQIOYai10m388Y3wvY9oxHnI2H88/aOYL7nHbo4h0pmvN9OpSBWn2eHGq6s
rlLp32EnwvQVsMpwryEDvP7oTJBRCMZAf/O7sWZlvDj4iVBPqcYk4rvCyIKDP44M
Ywt3+MF7EAOBp7r6qwN+kIehVcMbKQmDK1t5vv75r2NgLhHpz2HaBcr4yPQSDM8e
4a/50MJ3OOLOWQoBoahwfI2zSCyQAQZQxnr4FKiTGy0+OCEZP/JmZWxk90PP1Blz
ltRBdZ/i2/2q+8JXc5+oMNMD6yHFMjKYRHAxqfMxYzqTtcJeBCrlGSZLHdnRr9qm
hU+i6tn9UC39ceL+m0lTxLDzP5eiHE+VvvL66tQRMXQ9jrSHxnEcwkbGKXSTVBdT
mQMS+c0fcix6zGme+SXiXehfE57O648h8TnKS8WUuB4AR5xibWKFNTnXSYq9c6Ut
qYn9goi70W3r337HjJ7tP1ix/GocSetvMyUzjlBUu3KNSVZQukXryHSbS/Tf59Nk
MY0FrZtfjMTco+/Q9zsrEKki2Ub2mxCJKDOCI8DnoE34lZgl+6//Efms8d6vJhay
ZPHOZNVd5wT1CFNmKc4IvnsG6xUFwuTbG1w2VKnQjefLOIsOBwYx85DZ1WnPoHIM
/rbeTV82VLV5YsBXGfT0D43whFBhwE7owyWCpJC+Boe1zzbI0cBg9d/9WO0J0ePg
eQUV9j/3QAPKek7npRpOUolVe9TtLGhw1XkJTzXizB19m/OksHuk+emSBL32/bl0
PCSMJq74fD5ehVIfMYwx5Fv3RXUTksFAE64WINMiLurR5w5DPCR9F/rvMtfb1dIW
0Phm/7yHbtuKIuQqa0G0leC3EFzLClQcNZoWQRcDJd9lRLF0o/Mn+QnCarD/da3W
3+8AuYa7BUqtF67HhYCQQVUZ6f64zk9yLEveGyuWe6WTgcAfwgvE8dTwFM5kbSSz
iJuN4qGt36jVRMezKm2qNmw7vhbATqtgcji6fXDJwg7kX6Fb28uCS48K3neUP0DV
2sRMsRyuwnbonAVZzFTr3bUSSMruttYKOaVay2CRYecfov/6099ahaeXjDhNr8/u
Pczp668RQvDG92pdcfToZNfDhxTC7Ej1Mcp9bPj462jKgk13+vit/jpe3ZA+FGfi
zK3vAQM1E1KsGE2KGmKkAe3R8bVa7gb7/MJqoCIcTc1bgZr+voFjbpEom4l0yTwt
4pSzPpMr1iHiinFyzlKGZe7JcsgY+Il0GVZMfJno+sHstNVk6VIUq7C41kBX4rbf
lVemcwGSMelV3tX/q8G+nVmglgt8Os52psOAyI9LiIJiajH4nXKE2TxUq/NX9rly
WVZ0adDkBo9HrZmqtU1O1UZ+Sqd0ZZoUvquh4vsG4ocSrw3D8RQqPVaOqLCP2Ov7
Xx7go45DqpZFIKrQvovibgAf+yR/f7uESYDjYbtgdAMMERZS/Qujc4fEqKkx4YTZ
mvI+Au9O1PDs0xJlMFt7CsQISidAofj+qYmzj0NX7q0+4ypr3O+wV5XdCuBZj28m
5pQ3faoZ0L6X+VnKIYPdKx+GI1LB5z3WHwbfz2m7xBQv5zVgbuZL5FABlqaA7+cM
WpqyQH6d5s4MgvsmSSxJ1XlwC6epIesOCHRqLmYvDo3pj0kXA0YkFKCuzFTYqV99
VI7pfptxjZGNnqceppduuY4ucGWWBy2imFOlU3ol2ReQ8TLS+unrBBntR2R9EiNd
9MBYOuTsuR8FtgQIzrU+EF/3TkGApYNZVoxB6/1ulobf8snMvqUpwLpqH7KIt7xb
uxWZiyPeqyorBxnuwbDLHL6ubojLJPrqG7CsBct8aiDonLleSiLKys20JlrePkoa
rdpjZ2SiVhitEzre99EStY1qLMVTQHwXyCGXYm5GTRFWtmtzuBKE/5Cnf6UnoulM
ZuRLaFyYeBZnUUdpVSJpHvpJFw1m201vK3RZ29YkYiC3kU0hk1eTNsshAy1aXOal
1VIWd2W1Atq/PyUI0uK2UzdoMs9txz+8Xar61vdHUiXafkSv7349eCkCqEsdBM8O
jfQxMjT+EbD7TxP8JK1C00v5xm166r8wWM4bkCh8go22nFJVYx9/MIvmqhPUqxUE
W+stztQ6GxVIjvxh9/hCKbNlFMilYo05FxaKslir8RvBl3ijAg1CyLFlaQG7CjNT
vUhaX6GQo6g+pSB+HdhA5GBSX5Y1UlETzatqRCS08SSyr2JzCVRo/nVLL2EeZzH6
vOvc7kMV2Vo01OQWtpb/HI3TkkFVwxjb9Re7tWIGxTPG/E5y/6/L42ryVInsb2qu
RO/0sR//1OG7EC7AxGPN/a5x1G2YuDVn6aZoLx5ArYbwn3xRIMsmhX2rt9DmpELW
/B+iscHed2+k1NbGA5yEwbzYd9mBzgprroRuQHbh1bU6WTHxZ7sUKhKAWxDXYy8Z
b11q8b2NT7tnjbe3gNQlguwFPkE9Z3VH6IxrLXcMf1q2Dcy9f14auT+efSpOMsOI
OAR/wKxLFM37h9V8+Tcevy0VfQNVup5mGXIYss6i5IYIxYrbL+f8+Lyc3FQcD1zH
jgM1xFIxoNl8OwH7RiNY+SHGkMXIYFXY59O0nMNt+S4zZwrcVQokl7YtERMFcU6H
Z5s9vv5Ry4RneCo/vMFgeqLfp9KwIfJH9J82VO5TeeXfbXjRcFDP8L5vXyK0jJ8k
jNfVb/MHezdC0iazL3c7edCeer5+XQjjY5EKFBhh1afSWShE7KIWBFF0NloKesBm
dj+iOvy//nMNrYcOcrNrJDHWjs/lWcZUgM1Sh9Cu6kPGTbAXuRdw+S73vo12YFN2
Rp0Fl4rdEQQ/ZJpIRLmslRryCkWQw3KRpCJ+Fhi8X9x3NEetTbQsYDhmMPPVSivd
mX5sM82F0bJbC05jRl4ig/onO3ius6gg6J/g7iW87uTxpRSw5fNfin88nAXjn8L1
x3b20bb3dXGggWK9Vvrg1J+ZhLSyPj5rnF+A9iHApPMAX7JWFud5/G+pvzkLTFT8
/9w/qvsKth+FeBKgYXjj7MsRPsLI3BFUhgnXHcK1nzR/cIPWn3+ALT46gJeD2jry
u2M7Po712d0qf18K7t1W9s7hMEMb4VyyQBbHgWlGjCN+C2nRPC/khjFfe7lqteWI
gU2QOTj/EGFdXKETAqRmpWlt1TPxtW8NflkOyITOzmrVhvcC/PxYp+jnZRZagl0e
8rrqa7IpR0R7QK2LaSjFZKfe0zCuXhCrQrBDtDTl/Cbr5kgYYmXRNMnB0PaSDyZl
bvhnyfaKaKJ5lLe3/0hwlUKCPZweRgwZNKizQ+6MVFleJaezJOu0ap1vV2nSJN8s
u9malS5JvAcwY54R9ruB+KhA7KWRiBDZXxIvFi66V+eSBZvT0m34bHJWgLqcc2gm
Lf6TO4b+FR9Nl3oRXMdrlryIRvvuHRGGDVHGI1TxhVgXwnwThJvmX1+k91r8IsN7
LXiGEvzkTNRjftYDiQLpwyd7cr8T+DMg8G4ZVDiS74tR9Woi2OTGxvAW7/YmaRvb
5m7YE2FlRGDubIOKIifzs4/zeDVbiOVZzQAUgeV24DDK9G5VQvBVRgYbkHSC7y+f
PePzs9Fh6iU2CTxrOZ0bjSppRx9BeHdmVUcocURpB9ckG2NWatNK/og7wyam42cN
Zrv+VaVSbwEaEngmsSd8qR9SsoPtcjGwXOjg9Avi/PJO7TyIazQ260uuz1/fTFPd
ziTSjmAlblI+oSeG4tNDFAdW0h6BSTOVr4R/oXK1kt2Q+e2GuJfWUD+dKxj0yx1T
WqwzRugsqJt5tVjAL7YOy+ni2F5qssFDQ/yyIPa0qKZzwvMpmSDw7QFLCyWzB4ri
gv2z6e9Iu7QkS4/DFor+wVX4vj2runt0jstDhbsebpTizkHbC1rpNKt6mdErRuVF
P+vAN2QlV8RvoIO3Wr/IjFUkB11DEVLJFzn3RFiwa0lYK4STu4N0skQwb3c/FxaQ
I4+EbLitP/gWTFgzYZ5QvzfqCM9zZ4Iov6fXV1730E+jOL9sOzOTcHIIQA0qNI+f
3DgxkgTD5GSQMKHGqv93ZoHhBe1vWS3F8S3VseKOoTqA/CfZPPyufOUt9+/pA8NB
e8OFDwHVdPnHlbhXLbL3PKYAK0jcXXSgvYSqT6DjNrVT3GJwj271n5Ga5StzySJK
/I5c0ySoBXyOD8Y3FoEEFQzsiqdz/wxUDvAI1+LC+Z5bWgpNsTaKNqmfbCG7g2Xm
9/OfqYJkk6/G6HmUM1nwFHN3kIkKoqmhrP4t/fUoaBbpLO2SeVVlPcQRov07FgzH
9FHvJfYLOYua2r0R6lt0o6pcZoTK4LmQ4mxmjhoTTFXrE8qhQGeH/BIviq90FbFT
MTKuTLJwAfchLAIlv6i8dI56/N3e44KXXetDbx8kbeemuX+jRzIYOhVrrMoSFnW5
bqnGSfWL5wJMiHTw3hbSIOl5IVgaWsphbZ5Glne6zqtllD4mYjr1rx1NzW2KK6Cm
Lw6u3bMlb+Om1aEMgby4u1nhX+OvTR3Gihm/BeBms7rHVNZ9D5KDwmJiLomTM19v
F9I8NK5P2KE6Wn6DOh/blEGFOQR5z21Hp4dC0oFpkHC0jb13yBhelpMZAhhgZDnz
K2zXTGJxctbaElx7lhqEnjcYIliUEovUePWPAFHhljZZLV3VPzdbvgu0CxALfNhz
w5j47wamz9DVRxwCTSnoAWvnQ6Zsox+W8tdqMbojHDO0McmHcaLibGM5p10crFW5
u0bvZa4hhQ/4yl/mrt4CXJJmvC4GNEycIqaM0IOx9TmrWosaiGB/m9DtAzG9vxFU
l3G77kja7vk2Fx6XS9FFeUdosLTPp2U6K7ZyyQcmqUCWXjaMZBpwvZaoBkVOX8RR
xKBjmI8niCguwdXn3ppg8LBaOpKOjfUxseHP/XsKqa9GjzXMfCWHYzcqsFNJQgLQ
VuxnVkNi2k0PsRrawJa3d0bJY9e0q+frCEFwogTlQ2YaZaxHVuzKzEGpGGvqSB1r
IYZiMk9aAUQnoBIgj7qQAEFpx3kO9p41/evMaSEMzYburLj7e+JfhyIz/2eGH70M
PAxMKvTqmmHF8DntdSDb+eYgsaHiOKZADXbos3bDSHNMPUFM6Mq1kbqL/yQ627Hz
03c5+T5Q4MOOFKx4Xen9L1at4bwBjjQu/8QEgoa1K3oRdcKDvise4ujZNGwWnB0t
B66wEaELl/rWLhJ9KEwIIs88ETMC1jponJqgDCfcU4AXhzNuAmBdPimTEjKCL62L
8KrKqzdIKaa+t5fH2I4PKDeyua/SlUr3pdeDY7NyjZEcgJ6tcez37FxdpnFzb8d/
TZ/Y2TqpD7x9gLPbwDOWEaDVAiHZiatur4+R+vY90qCOXZd8JJnx1SxyZO6oOQx+
zmk4iJirFYHK6IGddVRRt50Hgaf+NfPaKNZQGybQWSFCd9b/1jqTDClDVQYyMD9E
6UDO3DxQtOE0gJ/gkoYonbc1/dJm+ERSYeKcs+/RRXRDFXJ6xu2evx6PlacA+y9f
bl57YEelUsddLESvtcKwMh3iyoYpTrPCVy4lt+vdVA11tpOexETt5woZrQqLeRpI
N9rKXD5lstLVF+IVDeW1Xb6naAd9m/Ssq7meAt0xXEyCdl5NfLhkdZ0vHpD8kFLd
hX0MCM3KjFPlIlMV4vk6U2ICdF2qENFBlG7c09ev13kQRDxchAhfeR2r1xAdnP3x
ZlMwIJGfB2qYylLQf7JawRNm4UKA0PO1is/RccIbre+kZrkqXOZWY6d7LhUkLRAN
ufbj4+N03S9S5burwQeiBZvsfUsZd9GQYjn6HUX1OnosSugLh6I4oPuA82wVtuG0
jtMqo4j+3W04api6dB54EM2L3zx8MVQ8lnfLwY3TAnP7pjvdAive4Q7RH4UtPC38
v9FVZFMQAG0WvEV1nuPnK+y4hLc0E0946Hbr35IeqIJenAO9vxfVJx0/utowXsHC
cslc2lUCb5xkJfNDHIUUxuLVfLEeWbd1vMeQrRO9YL4Fy1MlrkUFucDbpKKKmqBb
wYudCtro+9Sy0LMvL/1yoyQUjaxX2gxOc1bTv7+nIoFv781xz5K/in3QPtSwWkxS
tXe2aLf17CCRoE3X/gShexvjiOBt7U1Q6XaNzFbxsBj5U8/VCvfYcaMO6je51q+W
RRncph8DfgT6gSd8e0XxX5bNpS4TIgW/+sO8bRm5xs3euTiQfbhdw0ZHWSyRT4yZ
ZpgFTPoCHUFqrxiQtNQyCc9FQbtrv9C/q9jpKMxX6FxgT1NSM/IUGxzUqjgojeQE
N2Z26BXDO3kPwSiPC1kcgAmUUVBm/GqnSe8OcteTMYc3aqMLNZhOSW03koXjZ/ED
n+xGNGqc2WssJT7uEMUvMQjPbGsW1rV0PS72X3WNEFYQwVA3LO/zaANBoWestK7/
RnJ6yp6ko6/VtC5lAKkZzYtQK1S0hguUjN4I3iRZCirVmQ8zcndpJj+InoM26Sbg
0EfPMCegGhcPHIjcWl42bwFulN0RUciKri3EC9EQPU7ok0u9RODgVI+FxPOkLzAa
n15uxQ7xGBb2yet/vA+9lw+ju+Ieraa9FIV88dqgBRYruG4Xmbu4/+R0Zgj1jQoP
nWfnLc/lSTQMDroi679zOy5MgJ5a2MQpkW4J5dftIeC6mY++jZQY4ozSs8CSZuqn
wfDkMKNutn2HeuyRDYdQ3DAVpX0WqOhVdXjtOlY4DjmpyM6IE1bO4TQrijOyMizE
bNM7OR6U2jzugD9GjHHcQurD2BjGQ/t9ot8RU4KBq/GcwI31sz7eTlilNSBoExj/
7s5EjyELXthTdc5NUceeANsmS7PyRhF6zybMulMsIDQuQtPnf4GiUjCDmybDf8cC
soWBOAPOqy9EOko7qFVZxJ6n2WG7s3uYtTbMlK7CsisPy3odbzsUtmBQBDfI3mml
/L7r5jiLBt1zVd9ivqWLmmGi8GZunXq79tkmcPa9nU2dybuL8M3n37oVUtH+0W58
QA09XVyNs20Ml7u3TtLoGvPxjFUTjsIh+4ygH2o4EEIIe3lMfc/OaewtoZk4hxQU
GRS4k7lCvSN+dUGcvA7NfPc7On5tLMnSkws7TTkyXkEWTYM3OYsFnbReaop9PHSs
sD7IMq9x18f6bQQ2cdZ6Wbj7rbY5tPCTJbRS/TERwBqME+EekN5dXGuZ8j2vkKye
nrh2h2BgVSXscrk6wpwqXkra3q8TqqFgxE5EE/m8RShOm3XYEEO55wM7mT5Hko4K
HcqSIJhgzoqMq/Ww1afJ+sB37tWUpZaZr3tkrLVNO2W+dZVKOSD7aZ+Q+XiUSwK1
/kjNFZax6lJcUXE9a3XrgX/wiYouw0kp2FTz8eRUD9PwSQg/XB+27P2ROfyJe6hB
ZC7bVnEOASPfNDoVwO15aNUpnczcCPCGkIasKkBsDykZaXHYu1UKAms69aqm3a1i
G6Mb0WzMNzcvyk5FtrLKGZzUakrnZGXrYHh7OqhFu8tNgtotIt0e+3QaEr0kpyX8
Vxke2VpOhvG8efVTJUyp9VL0+XMAIivgT1Opcp7DkOyLfxcRwcN5N55F//Ak8P+R
WZI9aNmzfIkP3xyhxCn++jE5aSriEACFBuAR1f+o8k8cSKCWyASTLmBlCf/SMhBu
CRoaF7iZGTeySfZRrNOlmQTKcrow2NE7At4vEAVYtBaWFyTcJwtabT8lGEgVJmhF
kQMvdWHrB5vrmxqJBeZ+2elaC9Q+FRBoXJf2FS6Tdy6UYs2al/bprqp75PUOog5n
fWzczCJoLaFJhTTLlSx1WtqWTS7AjuoCd621ceycPLNC4nxRbUhgUNsC4p9TvmPd
RR1i51JdYpseatsZYBX22Y/XTNFOcK/YbI4AVK+io1rPdn2VJ9glVepvj/rAdiaL
r7LxiaEWSNzJdERrqYLFit+e4s0z3Y2WoihQ6hmvLUT3MsqmUvcmXN9R1Wb6Q4wR
hqS3iJHBJlzZwrDs+1Nk/eqi2nu/m3ZEc3jbZjvpcxwbzlRsKQAqWb9IsVVolCq3
GdKoBBCYGXaOqMswiU7gH+dJWw8BJFaPfg9HaywKNqxIKDYaRZAoS5LoSfqFXrXK
NlP7qJ5WNUJnnB0KhQxvLNUFWHh6VkmDTRfk/Pjxormo0AtKGaKOOKn2sHc2ADyW
sfRv5t2R/kce56SORAV/bR7lJNKuNUK4fuGEbMpYQxDZwU1Y+oXmkm/GU8vyWJjq
t6QDAEfPJ0xUJnQqKgBH4BYkLD1msjztVXegOi9ujmPgJx58gUFYfDVkhLH3w+x5
K1bRL7uGmDYxWa4rI1jTNJwz93QGHoTz40JiD91oOLHH6A/xxBeUOFZ2b5TUHG0Y
bqQQM1d00odgrUPdQduZhj2YrL2MC0xI2a0nsaah+5ogqlnDmUYcg5WMtFNReGoM
hrWK+SJ68DV7eS88+MIHN97Dm7TSz/XGYnYLOIOPCtgkcndG1ZQdXJf1FJqITlDM
VNl3CWufmg2dg4ztxnjY/ov4ODxO/wFl9QEy2w4AyLmFej7zzuKc74/jbWHn37Sa
ct+q9J0TH2ZZhAGmPNqAzPFynTA8d+vVHWzLeXAezG48Iy3WpIy2OKnDpES0iVtG
8gRtA+PjMb/vOGbu43ABxGWFv2QxxTaVSqeV2OlHdlu8FHfYYhHHHdLaCs+3WTPC
URtN3KqXZ4Sd+vzkO105nq2pJuWy/dLUR1ABvO5E+PsfUVMceoNLqrin8mpaM/UU
F2UO/nCawkXqwD1QUnmL2/9RITOGdTq0G4GY8eDzZhvhbbi23HDBsh3AxQMiS4Cv
Z9l5oR1ElzKPjjlCfnrgBmUa5Tvsc5kUla01jxCupaCFQZIkSi32y31qVxgTiWXU
BKjETUAx5i5BjSDENTOH9v2tEAJQxyBJzCvizhyLq3wW7juPfAMKDXk/RjnRkV46
cNfjL27Gemir6uqaYH9fvGTciVVvnQeNkxBKLhmZyFxYZp3HTRM+wVFAm4Wr6wBu
tZrURPrJG0mBna6LAgRUKteSMkzdm3sb1wywhpOMJtAdqfYb/UkHJ+HF/LeXOfDP
gDurUDWoCkbdQQNnK6J69pmIJVacwsQWzkYWj9b4QgfdFNfseIz6A25xDbxivMs9
dppAmaIeCOuezBXjoGTwGddTLtxUDLkj0xzci4m0Nl6pQr6ef2XkRYIQ5uSqRuo3
pSsi8T7pZxioLsoYXDqll04/dpiAeSGMQNge/GkqAJmng07vIyqFhRBppayIG1Fe
CTM4HrDOWofpI0CaeAK/JEYXsBXWmSnuxuJngeRaPFfIEp42MHaEplaYNnibURun
vxMzOKqviJPT6I0fKofz8bv5PWKRxbVQhXQXspwot5kyDt3U6ijZF47x4YlVqiDT
0wP2exPseYgtXSVuJy6orEeIYAWKE7l3YFymdeTSHkt0xGnvFLWztMuZo7IZqZXS
gTwGb3dfp52JJoJKFxNzV0QjSR/2cLAaVHi2AUzG1K4E6lu+BRsvnSgOcffS92A1
f0aTmgd11KaFnIipXc+U5NWHX6uLKrT4lrcBIO+ndJkMEkWLUdwLfPZiY5zK7JeN
Sj4JxfbfUMF190jatGjR59F3w35kepkBlVFSyEzHm/lCjP/4NXmsdzcCDLbp0W0p
RmNnL9Zb5CNoEdeuNcsfR8tHMqPvWKCWLNgHJWx4YbtTY/hksKZ2eREFYxxAWXE9
8GhLb+TqWvL71p0/LtgmuPIR4L4e9TZ9GrC3Z78nXPwdQ0tDpJlbxQ/ONN+7Xt7f
6c4QlpqSIGkkOa/Tw0AiBBEdedsdNEHaf424u3VTqyV+A8Vt2D9HN3pcAMKO5J4R
TfOPp8d/PokiqQBZNQtXQeBxfIWaeni79W5LqrZPJ/3XL10wh4mRR9A77EzbhwRl
BDxyPmwsACFERvvuq9DEUbg4a/lv9hgLyd15de+GLYYWDrjPlvMD1eeXA9f/w9S+
yr+upQjfdWUzAGs2UNlIkvzE0IrOXqERruubVmRYB9PtirnQR5axQDivb4I+coHu
QaZSVWrjespd+rT5w78Iy5y4kik6GKbK5nQFov/e5u1j3I4tXlkFLf2qwQsBNX2x
7M35cebcceWzDXBET+DWpIsJ0NE/0Su1vA7elvVa+Of9zrBPY2EIH+aBStJR7Hes
l3/hDa746tOk8e2N9fV/5vOitOTGbrsruSIaGl5zuNXlLSo6C+Wqi4ArrleEjBxE
cXr9UEHdWs3crqbD7sKtxV5sgR8/Pz1m2OQ9krg3n/9G9hFViKHJsq5klpmva7br
nhfjVh9tHZTGltwIbdRc0BOtw8J72tqLQ3ywUpEt3IiQt8190ppFfAd+JWeGfCnl
goMR6Ar8uzn0MapWNV4ReUgsvb2SwyhcveiSI/TIydvFyQbEL3x+jv7we/chyA6B
oKofp2xWodx2WyPm5keFNU8eC3h13pYiz1uJuZZdb7mF1QBMzveh9acK20ivnt8i
kF3E7kgNUuRpQI7lOQH0xJ8X9OkvzslW5d6WivVUqQA1ej9KFlxvtT6LdLbbWi4h
teJm5oXlrbY31udV9L1V6scGJvC9gq9xAiI5XE34+CfEReyvVXVMxXmxHCeiJI0p
n37YzQgqBm4Vh6TnUecOUirnp7+vkvBEa3lVfKOIxYYElK1h0MXsjwHmqWrK6f3+
rG1BJ2LF/T6ynww5M3tkOwn3EgOwuYrLe8ZECYFTMqzdLXne+Z2g2VrS9fjFOBSx
HAJgqurbBYi47jTrVM4bdq2NbWGGIgbfEAADhypM6uxblMJC2k3B+///AQ3oE0Oi
S0RgWZg1d/MGlfcVPjuS2q0BgSLIYob0TVkc0wJGCvpRi9CzOBsyFgcBgn1+VDUr
IypXkOrzo/V1guo5W/z9y24C41r6PjFxQWY/qe48MRGC/aTd415Y/DA1SvcgG5yC
vlW94F5DUsrNKLG6hqfoV46LBPmFrcmEERLlrNsZpSk0XnMXxDagHA4Px2rAPdHH
x0efexPY393GgDdCrqLXkBeeeots4xmwyjCMV5bq9YtZpvr0NHEOT8JybjGmt7KP
2PeKQELj6GFdVeqMeWQaXrTTLf8VOewNKL+Mguw2VzA339jgwZwkUp3A2omu2lF3
X/wNgBD9L+q59jJ0t/4BzyeBj2fzshGf/zsLoNByDvscDxxinf1IFTcFzugXyM+N
tmrkzuSs4kAgGrazH2tTHVnGYPHe35Q7MZgNZf7WT5VB9wSnI8r1e4tqv8ZIbFa3
vzrO+2nndPYVT9OEjK9Ip0KFdogvAihFijEsPU5qLoyZW5TYzT555LhiuD6aLMy0
xxU+iCmOJ9OMOieRzds5PZBn5K/EZZgNawL+DCom09KVqOZhndRzyKaTLmXsj/pj
y3FDjQz6UHctfnQkzwDnELNSHswqx2G6qA2oRrcT6H/gYfeA+C6dhxq9j5Kv2amu
LlpsfuJhe5Hfy5ssvTxT2q3g7/w8RtZOJT+9uI4XyavAaKnp9fS/v1cYl7M00jMv
EvMVB7QyXUTN1R4Jkp2+b/HRdg34DyAruE28ff4YCCcMKzLnYop9GY8+rWn4Y++G
gqAt5P5eFsBMvNjQ94xBjdw94h137caRYm3W1oDxQZSVf+QDOlPiG/qtd48GnA5/
x0FkIjSSMDjo5KCaa9vnoPzTfZjRjHvuToQSJCHaYkspIz7XrDAaQGVOgn/OU1tz
CIkePN+lTqyvRGC1HRmjzf5LvPfT6UEdV3TFy5P/oJN2d5s9KxmxnhDy1nkxd41q
6BA5EBW0PX4Nix/FMzSSqrncmsoJze4AAEIKICSIfDDIY9TAXgj4c+HaZCL4Nh4T
Kj/sKQb3SZzm9D+lHjbNnGL1V6lT72fInHPpIGhYaPBBsr/8mX+oZWEGAB2HoJOf
5vYoahCORntqaoKsMdb0o85KzQCrbaHati93mDKwBu1v2YEShZIVO9/sBOWoFQrX
uYI0ANkHFt5rWwLSiLiQiGTV//jX+c+09+Eua39QmTzDxmeT+PIjRWNgsRcBBoPv
bwCQULywFvxrl9bsqd5kTK7CQWAzAxjrEYE+swBVTT/xQhaGEy0ITwrH2ZwI6xg0
km3xUwKHK3K3q97j8Jf4EPrsLIn4iZwrAEUPimmGMu05xEildKD/Ie8ukymVPWNE
bKniA2cGcHUjecdd3zBLleThe0zBP6Z8IqUQ3gVH13vu4SlTgtOUTGeOdgNBzA25
gZI3zpIQkhQlvJlgO8KTKDRdFM3+FemZWVhzg6nzMEzHeV8Kh4LeqLD3m51HjqLe
QwECnRHFv0vv1/hQUQnLtI9FL21MNKaT0pl0st5sVeBtnwjpdNpMBAdweRHUbB1b
e+slNv5CAJLiUBxdiS88wrY37ege0Dw9BZoh2XdAfaL1mTRmPWYE7Ue0+5CkhFX0
nFkMu80q56qDTWyOlejHB2kzIU1bO0QPXU+j53UU6BaCP4+F67h7QL8p1CBBVlor
GMlq9heJEJS9ubQTiPdTO/81kDT85p7QQTx8VG+F/xF8ufoCzIdTeVE+PPMnxPs3
xvt7LMUk4Yy4if38lpJ9ku6r4nKcAVV+38+lLKJGDkck7Rsjr4u+BSyql5sLeYBC
8ChGBlvSqGvByn3DEVLqSC/iNwwuwh7Zunrc7SldoSmGRaaHRR52TaO50ZryFVya
6KZ3XnKK0MUqekUmISAok6q5iA0mNiYQusyijymBfdYe3ch4K2RPGphOurwRDl0c
OdcGGko6oirucKZynrtK4kdx1yJnEN1QAgogfysyApQ5leumgiBf5E8UvIABw5wU
RgKJlnkMG5ep2jh51CcAZJu4z4vcv+K3BlozjLoZXhBMR7Xo9VqYXyZuNpIRyn36
v0/OdwFSsqGi33wJJ28QRoEHUi3LC1S+uTbmfIKpVb8fnumd9uHZuSPZV+kZAghI
kmBz/1OL/6GzGhl/Th1EWzr4hMSCSjtPihyE/csjNPlBj4m+Kp2BHugtGmGlxd9W
UBYItTrTx6TzNXHo1EGNDZl0dWTCVkXSx6vWuH2UKPYezZSIJrzVp/HnfbjKW0fe
Cdatbn6Dxqu76qmfw5rGBqwO+U68aHxJD//eUTkkLJEYKtOFD0Uu5KWfZ3BiU/Uu
w+laAzK4MthbQLDu/p7yOXh9ULG8OeKWAp09l8ZJHbbi+i0H8JNvMFiHtyaQxASQ
1f0j1T0GIHY6yflbhp6B4KQ4x3vHr9MIbs425T25EDzQkokgOez36g72ycs5jAe+
dJ+6I84rtE/0xrUKcmSnHRC+hCaR2eknqz8KPPq+GqLJknth0HgRvpyCZJzUefli
/VKBdghdLwRBBcrHrwzPFra7t0fD7FXvqBgzeKomHaNgVWEgi4++r/o4HUQ5G67o
sulb1oP0GZ7rhe8awvUEwAsWzH8NKtGPzZ3EnMJ7jIEomkh1ET00rQ8T7GMznco4
B7GZ8lQH9b8iVxHc/qduA+XL/H0wNemiFwX+0Hx2Qgt/1vXKBhoXviSoSyDu9rul
GfvGhTNLlhBnWcJLAtrXdg1ycbDRm3GWv6HZk6Cp/53RJ8IwhahIzW8mITt3peg6
KHPbIf0fYAj2xyN3oDYzAcjuJTSLi28v3jBQasxljrCwjDiaJFq/ob3xy3cctsze
E6ymh0VYmCt882Q3vXqfw9FghyuHwY5DoLAx+ouY9oM5+qopKnpG61W0AAjm4Yzy
PSzqOisptNPWkcTaAfRfbkfydr99KkhrMSZffKJeIh6t/uwxt1l55bAWG3fV2lEk
d2tmUaSNeS2TJXhZzCl1VLp2L+e7NZWgbRMWgEqdHgfgcljgKvTdr+91zDUVd6Vz
BVb0cibGmiS4yIDAw9fBUxnpw70Rjm+xO7zeCLbHmhiwxwaoWBUG9Sk/RVnc2R7o
1VRSJG6znXcTNB6mIhcLfG9H/OamSoRP67J/+lp8OJCBm6s2ySWFlklHt0g2st4e
0n/zmlq7AmjX7x6FOvH5XA2B/3XXugXVCSQ15W9O9tuCjSJOFfPnjGzwdPfaXvXa
j8A4FuhHV6NdWbgLkrEUfA+bPrAv8z7k1IUGaDy4QOzph14QFa/eYFHoP17V5/mk
lmIvdSCS5w+4gsE5KjQY+8afW758DuXQmGKpj18SoQptRo4kWQpNzCEsK2EaP0u8
PszpbvPRiruajztj4cdsjHNlFsAFjDOm6HonMEQvIcBgvp1rdnbsDsZuWpR4tedY
SjOIprf6Ms6ebkq2zZPLALmxg0KsdVoLETYaOkO8osiANTugkiyQPzGf8naD0snm
dlmVIa+sHMeDzeDrWRGH/2mIVjOqeFJAO7k0+Xh8h0mXLw0K2C03MlBhXG3lhXEi
kN2cMRTkwg2+AFTriNZJT9SKWkFdskHK/QSTQ80grvMj4rp4OpRpz+UYCaIQ5ivT
YIN+TrKeiwGKz5PoVXv966IRlT6Sk+vZpYMb654DJ3wIZGVeKngNFXejhheVcflC
/CYnD4nSXIjSmYqQBcvZClAyrSw/NrKS5lgG+/QcyAej0qcBob7S//SxP7BMfTbQ
J8XbngZzN1wAmQMg7vq2PBbqheEDbaX+soQ6jQvUuuMQQjij7S5+QX5StQj7Qz8y
5zqrZcouBw60ddNGc/TAL4kcpJ7sbPVukJBP1z3FfAmm82FlSeUaZRC/JOmwWo9J
csl898bPpqBrPAnpBz+GpNqV66UM2p9+222q2oQeDF1Bx2AvF01hbT6O7Wo3tJ9e
04acDKs1TP+cngAmNo0WXVYs6RdHorbK/DA95uEj4nQ1oDcarY9LPSWGVXnSrZyl
h5XvF2XxWphlgNaah7s6OK2Z3I/UZKb+HtzLRo6JVPj6wv063zATNq5P56F7xUzh
EZimAKQ3AzEi9VqiroNxAlZhABKuHXJ88TCo6cjHj6z9HqJyGMIE1r7JIDqRtO7F
UQVlEJjsTPLSkQ5K769S7vjgoNCI8zNelL51tifmDuYRjFnPIdYsaYjHHOZ8P+mX
Ugr8KUNgGAvWTeKS1MfjmqljPgWiziR/x1miTKUWRv1k6/ChnQyA+5YWYK1o0YKA
FkvAg7xQXQ+84IxVJgnH0Rlwu50NIbunrs8hGwMTeu9a8Uqgyuu35Q4GDeJUFHj9
LryPa6gwxtkKO4yAtQGW/y9CXTqy++N+rOpJAu9WPxVGhH3uq9oKsN4rJ0eoHVq1
dxHXse+71gz65TgtKjDTPB7tAAvQTxqmFEtgVOMyyCC/uoNMLEbvoD8awVC/YHcW
aCCHyFIZcALx2P58Se+8F7OD95Ion0d8X4NfWTpTbgIKkULiY4BYKAjYi7eC2AgS
ZEn13NYJ7YXT5X/REXFfBCRLDb8QRBeg49mQ9PZqsHX8WdXAfDepLArYaalLkmRL
kjrX6i7L2II74h4SpStqxlvzHOcsyuTk+PdJtCFufVdRh0w76lE7/p0lLLiIQtYU
h3oRrf5KiYfs2rI/pNmlN8nM6yZQQqi8Xp7VPM7dZEO08WxjiImJkj165LGSX1Xm
ufosNP0+o8N1u7DwM5fDaqOh4QCiI8ib+b8aHfofWfPV05dwhxyGUaahhERjvo61
60r0oqc3CX8wCTRE5w9m3W7JR7iU5pougHRjTQj2BR7WHAGXTfaIEc6Rh9oQhz6K
/507HR4NS4JDRVWajYnKf8AP2jE4uJPPS3Mg8sTlNopQ5zXAlRNSOmpksLwIBWIv
DnktA9Tw/ES4B6HD0bJr11IIIQbxfpISTJci2f5cxRSiR/kX1s5E7dD2JLJhkw53
A1sPOqxubZhXqEe2a2vxSUQaX0RnuYuEU2FlvbanpQ4rhb/tJtnW3fT89q1foeBp
J85AKXIzSCj1rSH9Xyl7Wf3zYkBZ7PJM7LDfqWKDPivjnSieEQ2PK8lf1pUF/rqe
OE2yQ52nwwBIf5C/9yfrYTrphHKa45SMXMcRRvQq47vKdNBY8MCQF8HoOqDVXuEA
7ks/4dJ0VAGOI6T/a8NCQazv6J0UTm9snalxWI1LtjoJZ+kHa20CM+JT49JqFObD
rTIHjiZOCIDZxdvcxjlPf6mmuJEK48eaao/123xyHvHwvC/d2FFaZoaBoLI8v3L2
ItHJFCbGmhgAGvDIdUutspgZWPXEupX3+6yoy1BoXIgVF0tx0flYPSkaQ4Cejs+i
9Xm+L2WPA3DaKvcPulqPSLil5nZDX7MnK3RtL/tciBT1ijT0z/L3CoDYNrZF7S6m
zbZh8yYJMjb3gmlmTW3pY/mCLC0UjqHNLB94c3hFhmHWx9H0AGqAolx9bDu2+mo3
tAino9OR0pqammtKNfx/iuiIgELuTCLaWZipF7LAFPZyijbQcUtXhpCAkIhttabC
DBAwQ/ZqQ/cKvRClnHD5wOoEIj6dxUyqS3/fDVlD5JsmHIRI8mB+jIcYG7NucM/w
dKJXQz7twXgNO9pbvxMeSij1uZS69nN04xx9uKkfJ35cQ5ZfbWE5Eqw0IFodr557
JYovIGY4qR2dwWaY8+sqwQFFKzCeTR7HCly5GkT2Kvr62A7Bw6dT3ISpapnB3yiH
CVYT72XBozsx+e/m0eN6oszoDNJag1WecILqC9YgF++wK/CEliGjzaJChxM6Vm3p
ZPlp/jAJg3wDAjWce3ydYvqEbT0usJLyFBSmCsbRdqUiHnIFG4v8e05DEnTui4Gf
cYFHXcl7A/CLqESBiJvhLOqxr9gcDwQ6gZOPxZXM/MfaW00IA7hPEgkkEBPgcRIA
vOYl2jw20NI4FA58wIExG49IG3yAo/VRuF1UKdEobxH54ef8MBkLdfk+/wOeSxLa
IocKT+caEKRnbRtb0DMQ6Y/XF3UAONMwm2mpw0bQHTri4HlMwF1UuAYfL2M3nDyb
Uf0UUATSlwDvkkbQs4SDFyUlhF6o1LoF5K5rxLaH7pDU5eaitmMMZHOizXHV8MCF
EOXa2GK32N+baFyOa0XxcS7ExiA0D2E7VFvI4alXZXNaL1/QXZeX6M5oAgt7d2KZ
Mb3VoxviPti+ZszDnrCR49lt9Mk7hiVkGZqOyEH6H/iyRXHaW7L5oG7bmQCZd0FA
ZBfmkKniHGYytCfuQkHAHQ3z2LCy+7lW0SOMMWJqTJCabkYl0K+ktL6oO7hUYQSj
NvuX0IKm33961th7H+LnePHzq8OXragdGYWkHsoL147JSu9I56Nzjule+tsmPRdP
wJgF15089lZrqZBP0K1v6iZHJBbdzmBOeVRTnNcQHSRLRdAC2HiQEPc5hL454p6/
HQYx4Q7HnSMhAZ+3nAmpqjcU3LA5ntzOpZw1geOlAN9OScasr44+ARh4oumYuRMT
X2Cclz00NObS2MVytl1+Qs61tBThO+/FkaAsWlPKYtoDITKS9L7LBDASPAlikeq6
Nifm5qCr/yQWbYZgcCdVTZks2b8YBORACOLBpOYzMWcjcCfyCOWgUsc/gcNOxWRg
dBfW3AF02FULYM1Ogw7dFkUdHqtVWmjHcG9o0fnGpeqLUxkhnsdNQ7fhnJHtjGdC
en/vdtAoO3ljP0AbVcL4w++t7BZUfPppRSYTyzuxGfLtv+MwQUL6AJ4FmVVV6iPt
RjDp+7HL599C0nn29X2kiON7dt7m5wfLhNLfoXuaxWRWElX8bAe6HeuPTH1r2yzE
8fV98GvSN3VJWpvxGBLn81r9o9FFvcaXSudjuHB3IypbWLLnK+vCLuAysPP2/Tie
HmVt+EfzESzVD1XeH9LPsXtEWF6fCZZHecSTTfuMiU2H+ZrT7Jgr+KWEewkRkG6C
vRKXx67nUzLW2DpO9hugNjhm7l8C3UCwG07NVz2YMAHFc6k+TUMu6aaDls/VpbbS
l+9xfGb+9gu/RLf6fAcrE/EfvRT5oPcMzdrxdlFzAqfSSaOnxIPnjWoN4rsSUBiM
3HLHhJjl9YUXosCR/7DI/NbnnKv/j6HtYmwbbC/INtBjs2owxLfnEtPKovB1SXEg
E7j0cCObcGmyuGST5r5wcGtzN1rweTv+3MQfQ258aLbd4/afDOwdHYQCOizcgXJH
FrQNH5W7CUcz/50YUDuW3sYZ+xm6ICpMcwjuEDDA4qIf0SkuAOcREj32zLnlRpM1
Hbe9Ty/D/wbl5T6IihF/s9+lKgi9fNq6dS0wIdfIL3x/Sl1t4MVI4RIehpgLfpIe
SEeBUDMDweeeezXdADA102oU9ilzuznWVdmjsxOLDgOYri01xJRG74wZB6H19HFf
FoJwma4nLBihbcQzueI+xS1bWVhp4L+xvG7pCVmmzAftUHGFikoyf3RIVCxJztm+
ZdmoeHw2hJffDM6u4+Tf+sUjkduFlRh+1ubYEKb5ZmMNRRPheFfWCmnEgm4U7D7S
6SGfBenGi4lwH2PmTHpwsu2lzGyGWPX3+kkIXwMtP8C2PUMX0jI85Bxsm+VjtT2I
bp4Y95H4lRV5yxUyN9SJbE7R0pcPxAPaPxtAgC4Sj4PXYOKpfga3nP3eoyLIrICd
JUaYYMrJYF3GpND2ex9TnYaYTid8b6hKciIF9pnS+96ijuUUPj+hrygXjTmXvcL1
KFhZL8i3aZ8wjvmpJlDblLRR4H8SHimpztnNYL8Y7eFYJXjTiI+bu0l2yRduaGUT
mz8FiZQpeUaPRM8dpL3xW0BptO5RP1Cr0RZBFDqJ5UYaE76uutlwBYgqZHOWojYA
KAnIv40iMVx20xU07oy09t75Nll6BHHxJqQ/UXt1wJBISZgdc6TaduPdQieI/xCM
WB+EN1bOorYeXt57XUCGby4WYHBuiijulbWHYUEnskvqQh6IoGzse6vaddYcHJ13
dm+i9Lz/S8HsqGxtOXLDi02mkcD3mS5kW9AwEyVDimgqcYGVc0Qm8kHpQjcWvrTT
EAU6m6ZLIeIozOEdibPoJk1KN9bUhnHIzr5b1ipjrnK/TiL6FrjS/uPtCxvT20+F
IYOmnO8OgDjJeiqsxAS9VHPVhuoi/f4HxMRiuQDP1UrXWmk3C9GHWPNNoPaHOVgP
voWrT3Wm+nuJLc4RjKvnq6xZ6HRTFLqdyJd31fzKqj5AJbN8ZxhlMXxSfla6HxAX
674h7w/6YhfCo2JaHDqUxuG4l2X4Abuxwrq+BFxuupDrNqthuEqlukm/D5edgbf3
+AHDPNQfSUDd5pUeUuELetnmIcmzRiThKiygvBw8Qlgll+DsahMHs+E9LzxTZ4XF
igLk6nThXAqF2fv6m0A4lIrqRJmq8T2sr/GbLMeJ+2rGXVxGZarXeq0YzXQlXfb6
nQfUKkiO2PaHJvrQwBYau/HTKJZzkzwCGaLpsEkQoL4QZ/8BJUp4ozAvPCMkNZ/W
fqziUl7FXd0bo4z7UlEC7ADpS7Z7IGnIXcGZgPwqn+b9mP7Ylrih1EkzyKJA0y3b
N3klpXC3bY0fEGWKzh+xpWdOLbdf0lpc56/REJnqC8vTl8mnRXJQo3+iRZ6TCuxr
WoJbDB8FL6bSEYvVSRIc6u8cZLNNpIRV/dAz55r4nmYmjQu4gA7wAWozoS1RA+Ix
KQRLHIXvuVsfL5Ri+idckxBXDxF0va6r1S5zlQlV4s3LuYgqaf4Y77ARFFwhGKQI
9kf+KjGTeVDIloufHWOEc8jOn/PkS+toezVhZq6Hm3fye54HpR2sM6YYGu9JHsH5
j7gbZ7aM5hy5fM09DHGAuLhMJhde+LLjqKVXbMc3r5/rT25ShRT9RFldh8InkFDQ
WQwFneXLctvhVmd3NHFeOBYHYircLxWKuH9dMJ1sPkP6IQrSbz+fcWG/9dsA2qEd
FPo+R3ojJreDgFIHZjMPG6NymBrSbK+eeBYhB/V69O2LVBFGQOkhWTf47GeZlBmk
UW1XzBuQ54KWXUwuYh+Yzsib7Y00T7UfsQVP/p6JkhAvRp+Z5m672JXTfPmiwztI
Qci3Y/Q4zVLvmQeFl7D/Tnj1aWdLMxqbA3ZCyAgFbjKBuemhDh7/2xVwdgGV4Kbr
p1LFovzVcr3rrXMDgXlvOdoi1DXm+t3W5XPWG/hZ3TyjDJ3l+FiEfCTU1OTRsjsD
Rip3Nc01hj8NYMCwNBa55pCcm6d6JQXcj2L3ZX/FTMM0bXYK0lGOaQvxHTO6GQV9
xy9P1A0AO9s4XWY3K7GSuJ0icyPiu3pY0c7ERtzZZYIrzeOReWo79kNVFtg9WJRx
3z5DeP2D28TQ6fQIBnmvic7IvfetNeXPzipYv9bxOtUF/pmyuTpO4re37OS7FDia
0t++kh+CuMkQraCbrddWdx4/MXblD4zNXvydBhTC2MP51LFIFsQQaBWFSeUkSaGO
888CMl15PwJSgA8pPDTuxSueMc6T6b7x4vQ3WP5v/Q1fVDW3TOLnNEgrh9HyR3Bm
e3Q03mOrQaKde4CQyYkL7Lxh85VuKXn/Shayx/eoFARrs+xIMHjR2ItCZ7+bJZnC
C8r/GhAHGR2MqZ/RmQ/neDnPhQJ3baugL5uqPH8MBsMV0MYPPbYCbJGNE/12SOZc
jEpjTgCrGqdz/OC7dIDy3kib1fFecvpyEz3mkOd9dwLYF6u8ZYSOP0qxhrLDkZ9X
95/DRVEzg4BEN6+8Y6N214A2VA6sLKX3TYcky5Cx5mI9LC6hyBv5Axwh2qadbEHT
eS0iyEUOhhx60x7Ehpkm074ja29rv3uym3XU62F2APCc3A8VE6rYAQNMyU2zAkM+
bSRsvLJVuraC0mvTgyqwh0z07OnVuxsmjYW4htjSvDjVbL6Fk1/ELQ8NMldgg8pk
nRqIeThF3kWild59zUAJ6N6/pRqPRQiQ9ZnfAlg8DEI1lZDucI20bgHzBX3Ohq8f
m9gmZMD/wYqYR6HPGlGo3tVtt9SD9sBrcnKLGmAoCJgN9PmTdaEi83ngcAGA0rpa
C88qyJzdPayDtqHWgRKY5vu3JGx/QY4dMDUihE4bR3CYVIGAleV7vfhJ2W9F7jvj
3ASI/cGZN8+Rg4HXeFMMWIgHcIezzxnoSXnd/Hr/s+PtrIHiDUcLE+V4bqhIIUAo
lm3TKq3lLUPlAUoHbgOR43tsX3IAp4bnADcQZU5RO77VDVxuHpGfA/Rk3nMPz1bw
RG1+I3gWbmSZ3MQKVhAdoHorChnpOoFd764XA2heOI9470PnX3K9mVIMc7SgrUDU
0q9doksPOoMmrEQV6h40i8NKvI/JZTb8gGEB83pSt/e8gi4+WCXLpPwJgooS1HOO
2XvU4byZWA7Pk0Vg4hpoP+ACbpRdUbiU8ORZIEbC1Yj+2fCLmL5A2m4idGJhZTjT
r18hQO9afzDQMj5GxCECDcop2NgqhQ6OsWx5zjN7bfUuchLIhfHAgr0lQcrRNUve
nwn3H+HWyg8mtxj7nM4duRZWd9ZKx9qyzVDWCorLPKMC0G6/NFm5VJ79huATYIX0
cbaY7CgW5F07MeVFxknqrGLkVeKIV7R1HOUL7RqNKJMSNtVZLL+ERV8yogkGJX1D
zi6W9eYWqtS8wfHWEIeKfPPDjxbe8inzD6+xSB7IyJxI3w6gEF3g/0N2iZsqaSnE
jPcshUKxyABR+LujBUq2Glie+/okJrFdvR8/41yo1BPuRA5R4miDRvQDQoQ3iHEz
ASAQ6A1suXnLbEmr5UemPnRVwsytVHfVYTEzz+Q+5OWjO12xU1T0mYlNQZUAiqhX
1mm+oCWpmceCSx0c5kCt1j4euSNmPKGrOM0bAb8rvCUXaI2M7Sg5Qud8iBT67/DW
QYrH95EDEBHex9sAhoLEip6Sqrn0HS9kYeNaUthO6qThiANqlqGEBpiH61ClOlJp
nHHIRtDVZsmPw40mNt7yALDk5jyE1ppF0xpvHLCGoNFm6NQ52fidniDqk1Dt8fur
ZP1QNcgvdJmeu1TWGwH5aJBwmVkAK8Wi+3vznXMwwnmV0VuP7u8Abe0EnsBM/W7E
BWpqZLCx5C5OV1Jqqpa4kRldEOcQtjjbDYjS2gEJE1jAO7MvRYyzZNKYnVwTY8kw
MOaD0hYHn9SK5FECp/MqDNxKW8c8DziUmnltreOqK14F2x36qzj1Lqg4xqbRJBz3
bK1Z89/Bhp0nVdAWL9Ngv2/xb9v+2zMcu8L/lMxUxj+hlnkp3C5RG625CNrNt6DO
kSlsaplJ/SqMvYEXFazYz7c3FfoOzaggKYxeL062JCuLzHD0S0+1tNbneTnm+9oc
yU89IvmCQk1t9Gs94Aw9CLuwQuZfv9GpWGkVY5OFIj7gQgiFuj94INxf1fiVF08t
ips09u60rAHsjwFiSTNen/IVtRv8oVbzKkGUutJjB7kPdjvoy/faX9bWQeikip/+
3bAkJdaC/LvZonZaLGA8QsQTA1YcCAch7wlgH0em+iT8gJNRByVr0OfBNdBbky35
sViP7OU1mYRXI6QjaSGLZISuXR3wARRS3s+xiLvPJ+OL6JEQbiF234l+BwACuQ6V
boH6V/wsPDq/yeNnXAR22EViNBBY/5Q1x400i569ZRMC15LlMmnRgZYcKa0RDDs7
8jCR+MDPs1+2Glit+j9f/Tzy2peIWU5qQLGSv2FLWiqC+dvCzoV/1A2krXiexg2y
N1PWPHx7ctoICobSZed93LSUBXmUTPwMedwJQG3Gin670RsFI3GZjwNdTmdWBJx3
BYu6X0L0xM7eAHS9pxIAsYKLkWnviQXIrKU7Z89E9ogXh/XkLc378ONGBZ3SmG4E
d69F3447Db7wRzP+aH076dXME/nbUFNzMHv9UlYuKqPmyEzoZ8gJiJnrBx6Twm1F
wlgGZblTZFqHasIhij097u5kCw+WgAiN1g74wxT6Yx6BxS+ePeKHVQbTise//cCh
sFX14Q7e5Qm2EkWFmwGX98vbPqNAw+Ss7UKAq8T9TtvOURK4h7Y9MHehKzVgDT3L
QIZtDOvFEJoecOYQ8pTTOiYDfvvjkpcEU5fKuXAJlgzUV16DQyOM9QfO2F69Urgm
iITw1ugigwN27B9/5r//HAAAFzmNCTd53Z/1LPPiHttJunlvFcxelRmCw3kpOcMk
ETH2xcbWa5PD/gTIpkbj2582CpTj6H6rfjz7MFvjRhGNTzzVA4LPWNs8OExGzF5x
bqM4R0vr7VXuXmOkPX9g5A3xigU68m+etIjaT93taHh1jOWnWd0bCMSe5161cpFp
BaEx0of5Eo9fAjRGjSw+wogi92nz7XZgEBYSzO4q6RMTD7vu/X+bLPC4Sivg9AcH
MXacAxM/iPimO62YuVhB3pDfwoRQ5QTDR6Vagm0PeNf/64jovNgP+9i1iulDnV4Y
Oa891zmtnmMiURNOuvCOVlrNiKP3ogOC4c/MiAZitBeV+kAIacPIRm+KFn2hz4iY
jbVCI4W/7/N4g2wv540/YzgjDs8K9uwZfntbhGwlzbZVVjoWJ6brZpEz1Ba2VdbN
gbc9wnYhOV/jnu3nxJq5gugL909b0ruN+H0BOa7s6eCCv7tIhrjGRhKr5Rw4OPBg
oPBNE+KhJP6mgJKWH2VI5BqGdCqA0gy/Gt3cjtBj+YD21/uPyOV6Nm3NTUFm65MG
49c614ZKElWlo/kk2usq4xNVCHd4DPYbohOxpzUvF7OU/HwvGrKD7hJ5OtpZ1k75
YpzXFK0lEMMe8PC0fVaj9wCg5B3u+hKyetpgiktKA43Al28DiTP4fsMmBAnYDvJd
GDUJjHywE9JU4Lq9IN2ZV+ZJZunAZ+N4kn1DVwzbAiv+2Mc+ixhsWLYxYbaffVTQ
hN3DiMNYigqVzQjT8EJdfL+gi2gP1l6meWIV+YYieoMmqCnzvm4zf3gnS+78Qe0r
Ma0kSRMyEBiTk9KY4BE+HIMyktsGHBp8uKOAeTlo4/hxKRogV+pPyxEnmKiLYsh5
2rt6gB3XF3db/WQfdtR47uawgF+1QoaanNy68MYa3Ou/LBGC/UJkJQJSD+V+swG9
Mj12SPh5cXvaXaVoncKAI0/qPIOBJmXHxdPpwqOSiLi09ZIw1myF1jCYvyCUkorf
JmE3TNChiFE4EUdUw2344PA9TlX1F4g7nPde/5XG4CCILqtdRoT82UE5XfsS14i5
jI8b9DrdTF57GTUAth9myO3x7TqZsYs5gpv+Pfcp3qIefGuZM3ZSVn2HlYeH3iQk
q7TYAQGEK3eBq7/l32rMCsQS9Yx1CU42C8x6jjCoF9zK7eQhdvt+hALvWwf0iwRY
9/llSSSkT6l0e1ldU7e29k+ebmQYhVPwXPpSmfMqyriw0ZwHrTK9anERUZz9sXiu
YDWEnLOs5fPfUeqx0mNRGDuNRDFMYGcZ4zmjqpkOrddXzKFNnBPAnK2TbjWu0J1g
w/3Xc6R+r35Iv2hrd5dfbzJArH97t1LUOfKhi4zibV4QSoxN0s9C+GanpgK0VKwE
9qmqwSAQeoHNm1or6riZw2IKcRzw1um1vSB+KcV/L1VSs7dxfJLzNJ6Qh7bGs4DF
UvNysQTerrlKdTEHWqtTek4Vb8uobDpXeZVtk09RWxJcACEouohF9vqGqBXPOPIA
I4j4CV9ejQ2u1Qyi+3/s/U6IvmNf4tboDdQeZIVz+VdY+UzoOu47hKL0eTQ4RXYC
dvONuGre8EUbw1j+wC+Qch7Oi0h1MBLNzxXERk2/Ye7LUnbEJG7E7aNxgHLLvyia
NhOzvZNk2E6xhf8t66Dd2rWDaKQoX1ntclwlRxVQtWwIE/WOVThD9nzfV/rKqmOQ
gcuA58UjQ5H3nqOMZK3flh3jMRlmvD7w4neiPRIfrqxBuSHyzRwNQE/J+aFoehJL
Cm9stKDW+rTKAwnh9wW/GU/yRmml9oyOBKO916pYQEq2yWyqe2DS4JgrHAbNBqQY
gVssZ96FPyBPiV3MNEjL709aY+Kt34HL2pXxlNaXtY+/M68tfOuLGbKj6zvO26jm
hvLrbQwvgV2HOOisJv/3qjfPH0JUll6BgnoR8kIAPi7DyIwZROkTIYnr/GPEKvdH
Ugqkf9mwuJpONwQbMGdhTaAtb+4GT3Z73vi2R2d3VH3gXWNm1Dh+JzLSf/esZVms
FpmyoQ70IJws1bybC6LdWRcPqXQwZJz738akkBIIWGLWI3rMS96ly++TentzdnUM
HttW6+oXBcroxQqYyPIs7OKrOLGYCgaESWV4aRIBVHBxeRWUQAO90q6ej21s0SEZ
Y6pHnwfmuWvYSBM0MXIptVkIkrDH9Ps+CAELdcIsIuScNpmomXaLXjs98s1Ie6aW
hqCYMtMZ6+ou053HExoPa71y9aAofdfgkvtYv0a1G3osmbyNG4U8Bmy+v4M/QUx4
HcS5nTSBl3d50CirpDiDdh8h9RqPRmjiLCBNbk98T2Ptty9S2Fol5VhMsnFTgm9z
h9Ti1Yl7xEgTROqfu7Ny5hvcncGp7KUo8rh+D/3ucN7J9lemYDX5vQoxXyGMF97/
PtCiiwO99XdLExtLpgRzqkz8NF13aOFZSWdHuBMjNC86La15Uwu+8MA2CSP+Qng/
Kbw+v2H1xCpOS7OnLWo2Rn+iLn/2ljlWvhvEEt+ZBmpJgNjwRuBuMfkqYJ54Wj3+
9xuo63yFa4d1kNUHkX3vw/3h6AFDCf56B6AmCq79vKDvRdfZatBlVmb4lG1iWMNL
R2yOyd1sARMhMMBEeEVjEDrAwOQS1wpAwprdsv1DKJeDOV2AifPWXac9r2VFOc/X
R/Tzvjbi/fqTGHBcWQcBw0WvVNs5BFbVKlZUBElFTOcPfvZffB0m7j2q847toex6
huM0OKkSTAxu8yf1n2/XQQCa7nK0Rnpy6f3gdJYfIfwM8qe6d+NJp86wuJ5R56by
9pmvMFj6M42/j5tvefMOSR/3sSfuzg8tUnQJVccnXUc4aFwaPKXS6RWQ4e5l3MBL
Y83B/C0P7dZudMgPCXUfgkfGJhvLesP7+KKdVu+CQVzQjnntbi0pfEmAP7z4L48a
OSe8yLV3SYijaaXdx/VwfGF9c0K9LFBsAnEVvI3chqENoNk27Ams6UZEfgupb8zm
UCLTD0k5ts8ufTX8alP84BcJgIb7RXVtj21MoImxFzTW9e2lh19fdypqWbhn4rWg
P2uYSiQ7eCeBChg00z/sKYjBh7+c/ReN9RH0AeTH6938pU41THhNJrC5v5njmcPB
u269FcKiWUL5q01ngGPGJS29GBSn6zTsEHtB/cyuh+cbLicN2XaKjGDEcZfa3XnU
Ve6d9m3+mq4xjsxNRnTtcKMKTDsDiBTe+el7tj1uhzg0gF2nWzAxlGaDsxhE+xMb
5u6W+TftYOz3swH6xl6y28aygej530r2nwpOxi0mVGz5Qh8Rzihe2f3aswtUSsQ5
R4f3h8dPmit2RFNStHqBCK92yupRGuouK0E6reSenS2/JjLm2Hlrvmy1KADhtzzV
YhMi7lRSy+ZYFkFXLiwIrqY6+BgorYetiqyANM/+apjH/6O1s9KYIGs4jI00KlMl
dFMo0XU3luHdMH979+eo55ksDYc0lFrzkUYdtcXZ6okjH0MNbVpj8AeRWF8bOSP6
zK92/wW3OgQ+HwtbGG/q1DRtNYL2TZchyFD93caN3/zwWnR/I2kYf1VKAw6HLR39
MdQAnk4eqwliY9yghLzTj5cgSnn3C8QPA6I5yvgI+JSewNdXXp7u+Wf9DKmSGnF6
MUefRfCdkLN2+Ru3BWgNmNM63wWUW856V6A2D6cduGgP2A0lJWv60f18BZ3+3U48
vaWomxcyItBdB3EfbJvPxmo1H5lcq5f0e0CATYYwiHIlS/D01YDAYZS5gMmq6/sQ
NhfZRB3wN7+gyM9Ui8sdmjS1A1hLCrgELxkvK21SZRBx2nivQoVRRFKpMbbw1ZAf
KJMzbDyqfC9lZiQ8lHRGE/5jHXi8C8Z6/ODJbLI7SeylxvQxJosjCf6X6Z6W7QQb
hD/lT3pvwZf28+4/RjLQEU/AJq8RZ08YtnBT1e3c/znyTu1C7Ce6zllUa4AUyhHV
LwUod4sdemxCrCf33ItdKTBLDiNDryFoAyiYcLV0YTe3upUPFkdnc+blK3GtUWkG
GwU29Ab3wHyfiiT20QgfTQSSmw6FaBdqdRDQVKi6wmtQiayxI7e/fYDGfFw3WctQ
FvsNIjj0Bj2pz/P7vk5g9H63UW7mXdl2A9gEu5H2XJ5QXKN/S3Uv0cjutnpJlCvu
/P0M3cpoF0Q46fDSvWOQoTa0xg22uiegAgtDcUlmybwG2O3aat/3VtF14CpndKA3
lihQ8mHidopuoSk3GSkrnjJlzw4z5TrJdh8bivixmgJoS7iWFTanrMDzZLwu//jh
nDcjcqHlMqYb2TYCCssEg1XtTE/MApPS9Ri2W5BP/tuMgrIe7Dzbsk9OMX8/i8mN
bpLStVEco53oeTW4qybXwJX/DSGxwVWe6yd1H6vPifjhe2jeBs8GIAOXXX2BWP+t
fXpPOfd7Ty6Wa9eMLxk+/TN0M3otl6RXRfqvg6mP6HIFVRATHnW+dfkabJiIiSRB
nAi9yC0XdzPC9TwQ5kiR6shylePURhkKedxSuGMU0Ysg7lJ0vmnyxETHA0PirISJ
TnW23bHgtFQeBs5iA05GO3quHN1mmXUJw5V5c/d22gJrKDbNJxAfK8zBnBCAPgxX
hWqIky8WvayygZNXD38qsC2Tpb2dGmwgEpiL2Xo7yL0xu4i4gpU451nyOAyOK2q/
R/E+8nBa7PiY5jbUhSLwpBN+Q35gT0H5kTufW88APLiidPtF0ePrfuuM+sTdvEiT
4lYnDOpM7gasMGEBGwr4NvbMjx2Gw+LMkO4zb3UfHS7Bv6sHbMShjzEOykRp95Ak
9FWGc0RpWuIEvSkH6uPXx2IPLR+iOHO46A6KUp+D99eCClfVCOFo/bNSPDTuzJwr
PpnYmRHFe9FcVWEgHbk2nKDO3nRFZ1hUqnuqDtFA1IEM/wc5FxMdJhD+ypUVfQmB
v2bWufD3AgSUM9+n9hTteLYn7PA4LVgSEr40asMYIBtvHaCHGzDm0nb8LiWh2sPe
4tAJe3Oppk3oMoieHREeHe0hWtQXs5e9BSx30J/0+l8FQ0XN8XH238ocNKlv5Bnm
Y7KGYXjKzopKfQWdj04k2jKdwjqbcuhSRyqsDiXGgNeyVM90MvMvY0ee58ttpW+L
Qg4d918Khest3IjCtICGnqPXnREKBwCcbZSEfgJl/rQy9sFvwCr9K6dCsrfvWZvb
OMJwG+BDfe2QD9yIVYZCzNALXCk/YUgWv3srJA/+cR4sRymRVgeVCVmVJQvDDiSo
J/se9vtx7yVpS4y+FUGsS0CR/i8qcHxyluvx+T/3U08JAMdvGNPxfMLjshVZzIdE
B+Pjap7wz+qabfB8gVL7OGKuf829gg8UmziNO0mryx+D35lFQNLvguPx30cZWL68
DwjiMnsHDhPuJuSKWPsyBdCJPwIfl+O/lDP3Kh5xf2i90NTisWNuDm4mqNjnX193
mJ4zW3c1fZXaiJ5KCgRjjEWonwShWjumCllNbj61F40alcTDMcYTzYlDpLfc2hh9
TKjdYpMDR4FwNY1W/nTnlSnwlIABesrt0oN23GuQWFo+ta/HvPzFodDWwsfjJfFo
lRPxaKpOpeOxnyMRDH4ituyJPhdnW29yLTSBbx3N7GUcremuAYelht+yR93O5E8R
0pUdijdAGW9c7p6ZBY/mGtrrDcyYXnoJnY6G6rV0z6Jb7hh4OIAuamISu45sbT1a
p0zWs0n+RlrrHMe9ZDYuJkKjzkf7HbZPtSh/aa0cNIwmnFALX9fkEp8Bg2ju+uCT
RVVhWesmOXrcw/RqyMa2oVgeKynivolOkOXSdMJD8kw/D3TuNCev6HUjpG2ZOgTv
5ZFGTXprnWPwmDzQ0Gxhs1BDaw3jr4FeutaZ9/CEeajxxTFjUoSnEkQOMwYMI7nI
/V6p/ODMh+QdK9W1Rp9zPjc9SPz5SxmAJtzKJ+S560AYzJP6R8cO5wrsXGo/LiUI
P4bJjirkI/JEMknEZZfEAvYcnIeDPWbIM7QboAr6afTgISjsV7YVwpJPzcWMZipr
nAZKID4gqbhfS3xRqNJw8at5N9FToWy+9qk6ELr+TbHeq13qd79uv+5epK0nbcQm
37cWv8nTJUpB+mUMvDLEoe2hWPPafJLziJ++wfSXj0i81cOgQrYfhBzvQhHlLPpy
uv926IEAzmGDGEI/6NUu9BVptmX5W2YjjSSfl9JOFW/2/fBPE0oxeuslZn5zqDSR
PL03zhzZGAs3wXpi0KKP1IslZooYPwSZ8q+KXz5sOj7Xqjt91ETsEQgt/d0p5O6u
yS0CngMYTgmAjzYyjRcXbYGUAiZTObmYHnshwtWoIvhspJtcB+ipXvg7cKT7B3Kx
SRdNEIsvh1xl/YeTQbie8QMeUI6gaLpBvxshM4rjTz6oWDI5OyHfLmE9sHAYL9IN
VFB9F9aWZxO8vkSFps6LKfQVncq14OfSXoI2BB8OpHQPcCnhi8M3NGHjcLT3fjaG
kvNkfv0rvjQJMkKJ+b02rTq0nhhaQzG3n5w5NXUYKzQ7NdjqlAeIKVxCc/4eioMq
zvZJu7IaaADcyaQkzQkA4Dh51XFgpWCetvifI3wbdcSZ5b2VcLb0u9uGWzu5JwPB
Tij6emkGfneax9tmttmPI7WkpSJ63KPQMni3e450B1sj2GCYzJSk+b+t5u8Bwp5G
iljrC9Tirgs1TdiWYNpYe3UYpHKCA2VdS0gqYk7ydvhoNB6eZFVakjxnACS5RSNy
kjC8kJO+1hAnvlWQn5vm8kJnJdEMUlRZEoDSayc4fQwRMKQAg7GXSeL50a+NNntD
Nkjbj1uviBnTWiAbDMPBEmvkHb7TqJUzUT+snhfKtDXyvrpa7s+lNsJ8hWcNAwm9
sAyo16AJgoZW5Mevx4/z63v5uj9iG6VNilgY//WwSpUp/baOKN1J90vLZiMMAiaT
gaDDD4dkbBHpGzHPW3dT4/FtF+7HWFnnqBT3gWI/HxIibsOWy2robFPJZY04H40Q
KGwKTE24XGeNeEXNqRRfwIPdrqKTjaQ+3RI4BNLcWb1+k60g9jdhV+tU5YjkDwyx
sfRe4x63+Ovzqsl0ZC6PKKOUHniUyOOi94HbGtQDLcm9PEvfzTR0lMHr3eGjEdVV
A/Gjs9jVxJqFmZS5wGdBDGKP4WLIM5mJLFbGsP88QZ/6yZmHYKu3RJpnF7e/NjTF
CQhN9/OhvKC/vacbi0MdfvQ/lbjuKUfeIGACDqY9uw1koP0i5V6IjprGEn8jreN/
Z4HOFouZxrXxL+ibe8SIHOofafw3WTZd1AWkqRuWIhsu1JC6aFfEjT669R7i19jM
Ajj/M6XY5uoWXHR5kax02TjQ5J2+KOiKD0ceNco1KcKIUadHO5eg5+WvkXU8zV9O
WKoEIuRp6Eln/drnrUgFMngv913+7qaa9EYZypynl2i23wj2U4ts2vQ4a7K2UNki
r8So77YIcbns9sBa4nnWZgZN1l1A5I2P/uUP6K30Ntr2oB2vHsmc/gSl2lnfaa8/
/sTC+QpYIpu9LGSzCEoqQYf49veEr1g7zugrUbmcgVlHhfesIkUvFSiMwvAs4RDd
WSMDhZy4pqiCKmS/zwGGa9ArargPQ9xCZvwhiG0kssGkzGRTcvjd81F2WZMg5OCS
8gbSrjQU1KcnmFP8oqINPQVelVhjPQIovRDL44m73OG6Kc7pnqZQ8vvzhRa2IjUK
xQwFXGzQ9fP+kSKDVHEnAV/jKXWtlaN1tJa/eS5Y6IrlJnMsY2SuFnFIy0N4/mw4
ArEEtu4JeBbVrSLScSNDNSHPE/ACMR4aG2B6T5NSf6Y9FGMCdHTJYqD8kVO74F/q
A4vaNDoAvT2BDRc2BpAXANzZiave5s2zt+N6+ElRd2S/Ouc9s8U827xrHj3wWmoF
X5+Unpo/hgpW5gKdbp9wxKeWIT1Jabo+UX9KFEhWC9AFgcSaHFfGe7dfBnhTUTm1
C1AJ3vi8ZvXsusXxKAqUmS1SHyipp7/CxaRj9YhtbvCqwUUs/ZgM39UBA4rU2bCg
uKR9Vfs41B9Uhqh+JRtqCKxnjwVGhAgI0/qsSkOOqwf01tQyw/VU/K0kBO0Kxrto
TPDunGlai23g4kISujWGC9VdQfIwpoduGVr5mWNiJ+fROAuitVsKXROo1uplnSOM
+q3AMNqcE1IEsbYOP/yteDMWQlJ/vL+AIiilzp4iDkNZPGzf/SUPuec7KTOMOkmq
EqX5Jca5Lo7Tt6IARsm4gMMEX6mGkgLE5TgT9sDu9cZuGWi+kIjdyppsNIP02fKv
v5JIi/dmw4Lcvq4lsficaEwrHCdyBqndDLKiXwaxkuquVKZXYjtXAcTxKmDg0fEA
kZIj0/gXEtbT9V4+RrhbUG8yMZyIbzc+EE7YRgnjttyF8w7+UMitS+2UCSRRx1zL
W/vRuull9yFGVYpOGK3eHuGwOvVZvrshc9AF/JWGIrUtsXjmszQ4m4ZA7lIAEyw/
3JVUUQnSSgar0H8+Kj0cVeKUXzo+w+j+G0RnOqYMVY7NW8qL95SveR0q35xFmcYu
hCwy/oBD9p/81NkEti7s13Ib4bzoxLy1jQsNdrun6aZpOCvTYlaq/gthtJDd+0U0
qmr/OKf92XD0uuRkgSeOjg341JMoPt+BF3Qm3/Kpw1tJgJNqkKIYtu1nh/V/RFT5
IvfnHbtRh07mAdQjPUjkEE+g5otiXvc+piS1chbBNeK6OXJjnO8cnlx5YrFGwhb8
Ge/8/qp4JJorAUXzyGjVfnvbfm7Kluyf/I+T9AvAMMx41/AwkVbfsQ4u+7gJ2MpP
9luSBf3ettva63CAAQzNeINoxyRxjlijv7Do+02lc32pIKnwk/KOutlixRlOSi8B
2GzBbvguNtEvcRxQnA6pmv3c8vTFklwMGww18B/cMrMbcDsZ8wyeBDGtY5/HLbW1
hHTGkiIyx45VhThEa8GzaqAVKNHmWNyJogZsLTXBlzDtcLYh4zu39HtZUYYocdmk
hVNBHBwBooDINu12Gmahw6zeH7MzIV5s9ylqkE79lkih7pre/675PKqH7ZhHeyyb
55FXEqUOQhvyKSIfpyL3dYgKGtqBAl7iLzNPVf8sluWlh80YvckDGU9HHhWyAim5
OGsaR4Ecgcu8Cv2xHuBsDCxa9uDgwTWP8skCtSGZ/20nk18/X1yGHAId5rv8W3sP
syEPZmsjnhfcQx4PFCY3/KDNy/pNXbmVeaxJf99JpEuPu9CQVOiR38Yex035bRCK
OI8xTGLwUk3PAzA2K+L8DB714cgJglaEQuBRJVknfIYd2Lu/KbwTttyRcJjMb9/k
dOitfo1YwY0d8VmGnhOo6oAnqAWM0aPNETPbXuWTr7YDrpLBYFfxZUAVSEtc7+7Y
5li9JU/qj9ITEiwqZpWvmpDWfl7UFY8jPzqNuPHJP59luenDgNzeaZnVgj4wj8qf
Ox55OiMEUQSvG3R+7lIitow6cP48mwxWJ7mOAvyCybafXA5sqpjtH0S5rdFDX5rS
zR4G2s3vkGnPIJzrT2116u5Eaa0x5ErOmIKjI5e4IEu7BwWuUXPS1VHx/KZJS7Id
WlM3Jj31cCeVb0LK8J7fu2qz7I8S7Qzk7VRQALF+RDA7eQypxu8oNUs/JVMcGvhE
JFLil9dVSaRlQPw0kKAWCHea2PPJThtJIeuHlVQq9HxkIsDWyn7lO9Wb+HAOJVFn
u8rYmhypcdUmaVzgr2SrqK9Hp4geXZrjyGUay3wrVGKS3JDgW1LFDEqjxFXJ+mFr
AavvcrCKVLbmD+PLUR2EoovEDeC9AI9ujWzt8IAmrZmps+YPkkm23C/hN4Q+/Qdb
wQ/rXbZv/alHRumkWp+Fz8X8UWhMco2xKkGvFIU0JJgCWHckCPQAAkbydAJI7W35
3VaZWUdEMcxPAqSfK3Cu8uqzxX9QuiBskN3hgS/CVlOTy4oatOwBhQYvv1W3rz8B
JepiwSgeHfg5dtKPJvEMY6z6Frh5k2W88EU5flknUjHOSL8BgeIjBlpX+t4YEC9r
pGtivbxAwGMvLm0B55gzp4Ba9hFc0H+t6x+zylDHqffm8kjvr4jRVIytVKfKlAPf
lo7GjxIs/Mp3mFK8QC/77n3g902SkYCdrp+KKUEK8GrcEb6NgDJbjW9C9PSik0T7
uDd65ESPOyXvKdPWFjoWkcQ1o13sM/gqnKM84HVimCXTJmIm1LuBJY4H16bSQyQv
uiX52B0mAiJYwajxHhOsk2QEuw3wYogNr2cj47q9UEWFY45A1C2uvGfKzv2ongDX
GWRJKORnmvRKxaWkzXpJGz1Sc7prFIZ4Tc/PDLa1u1tmgR//8ujwuLZfnbUJp5Xq
ri/Wfb4fMX3Fv+86dIhWonzjYkfw90POmQzUN+TBFLfiVqz2nWmk071b/X+MRQju
IOsr5mgSS2tY2VHGT0Qy1RH6dIuvaAKFil4xHzz3b1Wxwe7wLCB9AJKHWvVuqq45
F9btoT6/70ZyAm7tw4cewU6MzRBMeR9iRZD5UZT/1WWuYuNCmIMPUzrb5OcYq/qi
K4/hQfqHV0z1/k25m8AbQxLN/TwzqHPjvqpf6Slb+tG7c+hZ0Il/iTVRih4q5CIT
dW7LbUokS9IuJ4+XR6eLNM2q5xAbXyqO9d7WDswMm535OkYEgj1qcQJVHiLJLsL1
Tgt//VBUdY4BPB3XYhXWYCXBcu5DhXNDAcJBzPqrkNrwziI2nV8vNgeT7/jgo4QZ
kERpyyasMw3ofiJI8iHI0TH0FJ0NP6bT5i6fdOuHYUph/NEp1Pm9c7NOVP1s5TUL
c/xBR5JPH56IEvMcrlYtlFZiAuVcOrX59qvE8lFIFikCbiPXxsTfATS8m1kUG2jg
LvBchvtH6D3YNmcknnj5j8F+tSJTo5+177BoZY/mRHRaKEzbDTntl9j1U8TksLLU
2rWpDD/PuRAr/ohmGayZTWae5SI8ZEqIerD/j3iTW2F6iM8I/aEMF9EK2GmOPhBI
wwxnBuI9ggbHSjN5YsX8IDZHuqfiFg/UshKD51iIAYNonJYiDvTOZ67/s7U0eNY+
vHEB2b1Y6gLaykrILfQ4sF8rXrePPrnjLpK+LOz44ISfbgPVK3tEZIDo5KVHM2+j
tMHsVwPsHrOVQkXNQ/7dRuYRWaDl1xImrMTmIgWqsIdqro8mR7q7yaVmn0HWimED
hre/oNKMM5+F3XT88m5wJ2SZQTOxIG3iWctlySEmg3npvBs3Z81W9+pR+LuwGPYj
88PHh9MY+8o7RSzcuatStjWczEHfzdWmjqTiKzkPn3IakNSR39P2U36TRy5vzrTq
4FmYui5ueoe93BXhOFpJCcp5RXRf4ju8Nbk6iRJ33p0df3zOMPO21L85KB00SM6B
5hhScjIb+pW7YOKmno3BKYk6TuLoFaRJVKia48E3GrSzPOPaU8vRuGu2eqHX05W5
HgWE79P+BPEHUFIVu+3JcZWH9idMl2yKNJDSBNHvk03RV26Eu0U4QSDRuAJMrUBi
X+6yGr5+31EkjXSfO27pFspDQTVjlhYReFOq8Pb1xvGwN9wcHsTfbbziFLqx5vOH
mBtYbBobQz38VBUQVMgk8W/wtq/Pud0w5VZXJl83uUJFjWGwQ0mSgGAtean984gT
5jUauKkEfPXtFnPjm0VJMJJP9GNMbKJJ1Dzl9m0uk7c49BrCFzJeGMuBwucdWMuf
4NUNSbHBpcjy7Kt49h9AqczYewYTiLNsu8PpclQsJs1Vq36leHrv/hFajGDsKfbw
OJsQTbzWFOAkbJR4Tz9dRfgGUuovis6N5opdZZyxh26fNmn/9Jk/zSSAHlqDk/hG
JQkwwyNA5fLX3QMmZU/HKdEt9un3gtapVsen1n2alKhL8z4Te9/peLOCHhNz+erd
6ij+kd3YVv9RtcRUUbV5/OQ028WwN8rTT3XoaXkqcK5STWw25k/pyWUvL/RaJpZW
E1OzKhkjK+Q5XNL09jVQpt8CPM046DTO7aT2ULYKmHgm/Pxtt+fjRhnDTVfz4ZSg
MF9ra/0iYE7G46JdP5IWnkHj+5dzRYBfDythjfuFASlDZYtyHawzrCe+8yzXYaPA
4aed54n7qDin0nU5mJMWEAlfKhOD1IKgvHNP9G5w6mevscTjxD/nUZES3mN7JgMc
DAAc/eP+751bgEb11U2/er3JSQ+aH5dK06ymPHQXIF+wWDBiQuqxCelKjsIbzgD7
v05y7UoD/VE3x0Wm7uBIh0HukGKh3F/jm0P1MSluX3NzUOgtMeG3malm5QBdoVLr
KmsIMUnLCrdyeRQPEheFvn7OoquLDzPge+QmZjnclQPsrhgsXK/5VtBS7v9iRp4Q
SYenUv3uPj8osybIGNRzFdJoKykGUODdxpSEHWx1E8H1BCWl970mxfdN/qG1Y8Ij
RS1+/vKcDKl4PV3FLvLdXBpVXPgpRISm3TfhJ/mEaPq/AgwmmoSCa0ZBIz3xtErj
ORKWzejARqnTPOMWLJ5LEUpj6V10D49moRwrubUD+NSlSHyj6N+tJQxOzuTJA0aP
1xQ/FD/e7aeigpiCxb+ZrVn6D4JZ1Pbi/dYuNyrBwpOr0B+2WHc8oa4J59N59cky
5/YTX4qmScyNQXlg5oSKKNB9a7/wpLM6btfxM764TERuSHhwj31MXxQy47wvNoJQ
MzTwYp2MYowdjHORsVBg4xCGeS1RV7L86WMouQvHxhEgjUAQ7xwTl1FuKS2TT4UB
TLkB/vDthBa/ke5p3jVkvwieYVnNZkJ2qH7hzaWT4SKV0chrBymsPLd7W6Qil/20
Ja4cDrsumaf/Lh2btsQZKB6z4Lzx+aDr90tm/kepdaGlzBdGtrzFNk6M+9pQ9L2C
rXWk6gudtdQv6sAA1yiWEae8Y8Pydp7gItiA6hEFn/XCFROxjq23Vto0tIUqoJNf
JLrlMmwhSV9frxgPYTXJKN6Ajl5XYz1V/ZeJkzvbt8QJBJg5WNXS/7jBehE3BnqM
I1mt0YRTVxxZpOq6d1aq+TWlQS4fiRTeAVufHsO6AHX1P9djrX//wJca5eyYUS/u
OIpNEdYxzq3h8+QAsThbsmJomC/GUPt5yft4GQp6FnMLTbN6MyCPExbwTlF5Z0Tj
tWGgfvmBmOmxPxJwSFaJk0drP+uVDRBbKyPieeH+YS7i3H8PZVwrI9H75Nhwy6UV
Hdha+0kStWhenl8W1tuDdlfLfA7RYhHzfhFN8hwjcnh77/aqM4BGhfsknLncJFQZ
hHPFfhOqepouDrNpXB0ykvXSrlacAj5qIEtWGXkh58QRfAdXKK4h++VfODXfe1aJ
EYWoVBMlX6OUfJw0b15bpEsUbrqQvpNLdaRg6kaN815wXBii7gMky8kODX8oCQo7
C0113IVI3EuRDoQ6yFrvc/iLgUFgflwdpdUAvE18HVoGnBGDXv04ZqCHiz7CQxC1
LSqvSoMKwXQy8Ar6Gldt+PF5RdHUAT/kwmiTjp4Wtm6EuGriL0gXTOxqkgeXuvhM
fjYsTHwnPQP2cr90lx0ym1QxgZgLBT9AgAaz//vo9CfYmCUtcfQZFediTEUFx61i
EmYUutvMAe6NmjdLa6yHZPi+2HB5hE/OCSRxjegN+6xTYWIBaj9iIAiZcwu/IRRY
GcBdVMEEFtJjZODJlzdQgN+8bnSzRVITT/E2FlOf9dvQoNRQrwSYr7VU73bA5cEb
xvoqtUviORfonJrBxD2akpMTugBrF7kah5qJARayFSPOGB9ZaowM1UtmWJuQMLt6
3VgCDmiNfq7PsRbGzpAgAnwTLrfz4mSZ0iEM7impmALl6QwV85ARslsri71ORyqH
0mz6LlY1lxs7HAwnCnVGr3ivNC90XYRq7HKl92vd+Vtp9It+shYqsgFT+zLcGyTV
30dQmD4d//jLp2aXixGc+CEKWC1uipueXwSvjGvdKgtL1bxdlI19QgNTf5VTE1cT
3xcW+pHF5pRkaKlrm7XDNNbpfSTIWQmNNmxiGo8xltia2FU6Ciw6LccxTt8YDaPv
oQy5+9JYKGAw+8aAwFt3hC1FRC6bN6YqrgmA9+TheAo+Vu1IUQ5vT7QKX2MdwgU6
Cf/3JiU4hx6hgsYRTW2cfmqEzxrDl+tY7c01i+RkY9qbsvhqm01E8IMMy8A0VuKH
oolT3jx1jXe28GyeinmY4WGE8S3i5idAF1Ac3mdNnLscm/hU/VoAwrh+fLzcGXFW
Ne07oLtMlHHvttMDZaVukO+pm8f/pcuZrkff45IFJyf4ghjf7Ao9m1NWsqxRDrEo
pcs5KHLemRUmabbYtrk5yz6rD7fz/GjVY56x6FB06fk366Dt3MsHByhlp4BwHCAm
VyyT9j8o13/V0O92o6DljWEHP6y40qU9R/ZK9RnmISgfo5O2sGu+d3zhrSw5jAg8
nBkl3eQYc4QV0thQ3mQUSImur/lf8HWKT61QY6PGG6UnBcq223Sz5BNDUdbiopJ9
i5S5p0a0N4Rym+yIcVAtbCE4YHJi8yTEj58Ln+XtMSAVozeWMrT3UlGWfL1ra1ur
k15TB8SeUxBxwVU1/JUqQ+AuHAXHG0Y1kDc4sNVt6eJg6NhpfDWrZN+1MYmwRvhJ
qKbeIod981DsmICLEsrkLHh6Qi9bCuuWJJW+1uidHh7fzWW2EOrNi3J9Qlqp7gKa
jQBiKcWg9PZpP3OKL5dCVvDL+dfUOEfC+fYPms/qEkN9Ouckp3IEVX8MopcPcmpz
u4Wanx+6JUW13hTTWAlU4FJiEqeEYuGLZc4YcTE6MBziTBPEc/uSEKWcq73FQu8u
22zs8Xk4jCRcHeUjVSEoPvo1fgSDXJD9kuSA5SWYFocmVA1ZT+QdhQO2LUTHyQGc
LwqdkzqnTlCuhPxmj5ufT/HjVAPOL/1sCBqMMt0Cr3Zbi6cCECseHvlGx+Y2df4j
sDzsIDhuufMuQBZ60YyozMLFE092Ng0VkAH2w9jPhAI9j5lrUBgRwy6bVW9igyMu
Uetx6GgZytVPxrNAKjUCvuDRmHtpzAmhfOskp7TAbQirxCDRPGXGwKo72/HHgQps
BALTZldQckwBM1WBwR+IyCxC9AWMNWeG/PSnA6hs9IuIfFwaiZ76tPv8yTLvBiFb
D4zUP1djYmmP3xJGB/yV4JCIwWsDRr72zTIMQWHvC1KCkF5grsJFA219Mxttl9rG
7aRDtqMlvowEBAvpL6hdQI8QyC6qeVE68vHscehLMCIrZLP/u/Jth5XRsDc/Uf6q
T+I7ErAOYBfsjXzAA1b/6H+v8W510na27vQOm27F8Eavr4tV6P52M+VjyX7XEa/s
cA6T4XiFD4a7KE1cxZV9rRzgFnzqyZ6x1kYIauUH3HSpExoAUui8Yimjpk6pZYK3
3VMdhXs4cqUifTTG9Dv0ogzw34gYtyadUtfPkqA1A/DC7v4aqAs6BDK/dhKteLTn
zZY6AucYBNlirl7/493pAm0fkrFF46lXaNZ/EoG3fMx9sCWATC1C8erjugJRBJeK
VxDFGZ8YbAVuLvYRSSAUg2NT9yPIDdQqa0evVIB9oeekC0SUI7R8jcF/FPYPFTcG
u7tMlWTl31iX+KuXekgRvtPU68vxVVUtx5uJ8d5/5D2JSM+041lBgBDwUkI+OUgA
Z7dPWxDZRY51Eb4gdqI7fOI0Svr+vHMD0UmmzryRSbrlsIKHBMkUQ2/N5NkxjBZD
xgqlrPG6erTASmbQxBo/mwc4wqdNMx6OcvEL+Up8A06yRjrQCA2qjLTxE7zE3de9
//kM1n33QgcVblH0mutcB0h7BIeRr/V+rk4xZmRsSOVyjmw0NjU2Ajb6vkldeLAn
0xCeyAvwMjzkNXhsS/UkjxslouSXZ0AmJi4nSRBj5QB3o0RPFfgQuMRDXTEge5Qt
me+WMPdhmsHI4jc84xM+dOXkLblzXC9nPvDEXeZWr24CtEPxQoRJvR4HJ6/Q7Oso
iwPbMv/2+2D5ml23c133/0xx4cijxIm4nLPa4XH39pRUTnAaSQ3MKSSXxUAb0TOe
UWBUtFH2nZvimzA5+3nJn+S5WWxtunk01B/yEDDHzEv6BUHarl7KgF0+WVuUgZHd
M+ygV2/4CUoGtUPJQayGgIzCfNv46KpH6fUn/uTpX1wq2e5P54vyXsKn4qGrNhdJ
TSKOVBIJiNJ5AdXsSI4iVsyKJdJGGhVPS/QhmWoLzCjUExq18v7qKEUB25ZD1STf
AcbrKd0Gzv/vvS3Bri0rRKCRuuePuPBgD3fjEvks7ol7MI5RblpQUH6reIrjyTgC
e0WrXBAHh6JHCVPm1z/L7ykOsFejDE1rgpXrUCTE3N2DEr9Y1EiW8ifUQWp2j7sg
cCGIAVp3RMrlscyAycgpuAnvOUjdUMotLFwrBqG3FCHvWtmE9STsYzWbQ5VsQE8z
w8264478GF9zE96LhJ0Gjl02aGJm5fNRDjRY455avQiYbBTlsZgW0+8zENyF23fD
Vn4/3JJpYGM4VXVlorZLINw8iwQm4OJ1LtX89PQDj6xFaZj04kX936Z91aEVXwzQ
XkTEND0SC1DKXy/dKc8Y+pVch7ubFK7ptUb6pkroDSSJFSrMyTN+RGwHDVCV3EeF
BFSKn/YtDjb+bhp5k/3uJe/Taxeg5T2V1fIdaoKL8MlgZ6Yt0Ky0QgNqhVZmGCv5
2xDtYGPJAQk8eNXaqQxYx1h4obBY9UNn0moBDrUBuyRJdKRyACTNHnb78wAml7u2
l15gO0SRkplFwt/y39M8CDhf7eGcshgkZ2C770lHDBHFvYHAbhBTWdzKc/YOBv25
MTUc290FNECKTPyNNWbRwHFBuB4peNgHGND6KHVJHC1FnvEU3n3A1sczDD0DK2dP
637c4bte61kkfCCs/LcN//ZBd3OxH73DUs3Q9aZnuD9aZXpHixxyfD7SXa10xz7G
FpOmT9ClnZdWg+G460C7WvVQGdh7DJjVlYpycJdz4hfNs+iSkYPZZpTsOMQcca1N
a73KV820zmVGAi5PipNXpcrbV7piSY9GITiTBBwX0bcKH5xeA5NhzFuD8cJn1+iM
SnK41wMz+kuHULm6EQZa3fBx0v58YSOMcttJ/PizD38WjP6jshxB2sJPqxH+DPlH
3UL9UUM4Y/CSXgcwBgUsD522qeQ1WYj/ZIEMv8fPE+FKDJZ/mmeZ+h5DJCBQqb7j
8XywKI5R2uPA/ARXIKBBmvxePsQylmN8vzHUaZtKqsJpQP8x1yiuKmuDCwMt/EzQ
3HOeC8xqlXL1H1NANi3bXyor3rxFIeaftT7Sim8xrvpGwtSksMkdp3bXwqpbFEP+
T72h3Dgtpw6lzRJDnNbRhE6O5FItovNFzh8VA4dtCdVrYQBPJfssY4tfiGpsqi0c
Q24k8cdy+coRJpSeFY3BYOAHhk75RGmltNyAyBHfR2/mGS+xmRr5Pt9VhVXJJb3T
Zhr5aaFzUxTpcwBswn9ZA0cao2iwgYIu8Psy+GsdhxsSB9Av4nVfE354XOaWg+tx
BA1E2e6tulSsUrd/QXDJlEQ7R5RmdZ+VF9y24KzdYBqz3mpHOC+cEkuT2nZ42ZH4
cqxDL+akIll0ia318AZf1waYKS18AzmujJ+zNeaElRHaiech6UQZUJYbn2houf/c
SzPNulv29FMt9rsAarYp/fGgf5apMaZlq3DmvhAS2pZR7MXmN3hb2VlzKuJTN119
3vMF1ajHpIBgzVCKb8FRDdeM3mcBG6LjmlfaDB8hbVRkZYN19eiDdG/vAx3gpRzB
iyQyNr0KdVb2q/XLhHsbFCXqNt3VXxc9gOp3qrnoWpSGyoZ+ju5WGKPHMCJP1EJ3
pH07Opqg2x2kDSYVu9E5S7nUXh33dChyqu4TGDhOXUVROzJXj/CJGanh2gyukrK2
dPwxIWoEIdSKGDqUF0oiu7saTwnHjhfKfPCOR3HpaiSedmhUJyupvJed+lCE58Nt
13ku4KxMHhITomub5tfpykJiWHZ+wgTyxAr3lQuG7CEWaJ2a+5wsN7/Z5jEZqm2K
+Kl16hEP6ccOgcr0a63Fd57qvNC1DRywekxSGKLOG2eQdEE7C9IdVEDEsFXc4lmD
PFLLWyqyoUeYkP6+cJcEkd2im8cHp2p/f53j15toYXBKzkG1vzba3d1DNywSwC4a
+TDaimhBt/cQEQ+eVSA1rTZnxTM9dgZRhRllgVj92V+xV5rAaHj6Y5YKhsyB3pSz
48X+96RGL9VMA8RVStn/9NBduNT6dWdWnpUiVdWaFIWSLHHv79IAV/p7xjVeMWp5
kvd/C3mvHbHWKs032u0Rd12AJu3r2GffXSOwTOMnABWdOWcJww84dKsXr5q1Nifm
+PdrA4Z8umUw/wGtLYmFmGSRmyNv8h3fR4LEnXGUGHzS0onTPlAi9UpExuZ8JWae
bGvbUAvyCteinfXPPhDapKadCp7OyZ2qnmOVj/makZm4LC9w3Z45LYaDkex/MD7k
E/8QPBewnw2xgtJMRGdprZLbqWqG4nYEW29rFN0GYWTFbDXQelvxl8LXcr0R7ryA
UOSKUQnwhgF2ztA8aMw3YozQyXItl+0JyvDBry8w7KUyH6otYkUTEIrOn9fzcBWf
+9EwCmD9R6zvvopxKnukVxTBF0NAEbZsOoaf9JE56f2o87e9c9yD0Nox+7y1fDgF
/A7Pe+AXdg781MZryAa1BH37rBgTPYiKeuVqhEP9QJeUWpFE4DSSbnIO7ipDnpZm
fnvsLC3RdaRokZNqSoDSF1LQ35Gmc3u4uANJIcdaFVAw1/fCY3aiv3bPLRQ8fAkG
d7yJwImX9IYc8h7H9zg6StQwWG0KqfgyHSA02skx0/qgFAN39QCO18ST/4WMVvgY
zqaATf+Uj8lZj3yH5eM7ECialep5Qcgryq4Jg0OqAx1CvJndduPuVZm9FKHHmzLA
d0cdRBaOnUN0WKNMS+A0N5YzWnsvMqEUD4A0hmTWtrL0dZWDjux1uAD5c4Tbvirj
VBMhvmlC6EC7/UKohkReAWvWYR6+z0Jba9E/BU1E/KfY4evNQ91NLnXQghXsGwIp
aUx90YTfocb6QP2ZA4L2ET/8S1EVixOJ2/tRiJH+15OW5IRATANSkRSnoa5E4l6V
pQsTmyQpn3TKWLi00cBuqFx9vNFg2X6Uc9nbW885ltuIRI9kxcavoHlZkuvlq4ZW
rds42slXyBbkcNIoAn7aayELOTNT5xYFqhNFeL41Entb1hTkVIUNAaOFTmMw0w/s
Lmkamt5O8sXVnIRnejmBWbyBvx4C0igvkaNVuaPLr8lJYmpG9Zk1JQ4u7O4d6kbL
Iga+kpprS1HPoXrR33R7MRqffwcxJnDATi7MLMJrQ5GAEj4kCbv9XmSaIQfjAtEp
CWokhMXz1jtnDA3U2aMt+XVvgQFXEYH6aVysVzF2XPQ9SwyfVNTBKfOKFR0Qsxss
vNodOBpAo9Qt6tBqVGFBsg1V+uRzZrzkAJGcDFyiP3CHsfkrSzMlIxKVEuizATFV
H3mOD40ku4FNKxZsGYpXyxFiPx0zpA3U66jNj3QR7we3fSmbNNGIriDWAbl+k127
NsSn8b5ZgtZKLDxmrNgmUcLWxh5inRAp+ZBLECbWLd/HFGVV41PHdZFpRXe4iuRg
IXdzWP0cS+S61T0CpoMw3NIeY/P9UyM380M6CcQu6Mjg5OtvFUzcyaL/LmjIJr+4
aXtWbDInZ6zOCYwN8MMQvhDHDPOnJJKowPUiRyv32bK+4QvN3l0i7SJ5KaeedjGi
4wCw1zjJ2i9PdGASrHYmsf9UGz8YPfJkWsUbfrTpkagfSWx26w+l83/YX+8rkBdc
O8hPzLv90J2qJfkfXoMFt16/CtB+hrMgNUXio7Tcus4WRQBlyrW9F+8dcXoz9e/a
sZFr7z1xR28We5KpuK9q482quZloIRnItF4kWjfzFopfFpwE/zzOaMQquBxLMwEe
oMw4HRfGMMQt6CPt24sOyCFNUMIcS4wNOjrEG3XNxMuzL3MQElkLpyeRpEoh9WGb
TPXhFCNL+6/EnniuYqaxeSyVTU7q0nyCmsfpmufaVs8NHDTeAUTgE4ULu2XyxSp6
+c2tRHjXZIm1W00UVQAj+Q1gj8uoJH3SKe5FsndYF/cy5eaA5lpDDzCKjxQoiqPT
ZmSm9bXyb75R/LET7Uuoue1HPETbkopMclt96cBVELCUoa0Re1njIv0S7KbbDFt0
zAqOnf8bBen7o4rIJOv5DCJYg4757IKNh3lo7OvKDu9h5EV+E7UThu+RBx4rFbT1
na/ENZ7n1a9UeTuYV4m66PRdoCOdLI2LWeCAcWrjd+829T0A9C37VNO2Dy+JWea3
M+sY3NipoYD5UXyNGyneRlPNoDwkNE6cF2loqPQF+voJTTcXlPk71TUD4H4DfQXd
sCmg3FaN9+9VThIS1Olq25U7bt/vJgFj/fz1x7i+B6Wq3wZCn1QSTzfKn/o6YKfE
zvZGZPiu3ifPAk3YIAg6ARpmisiMlfn6dTz68F1FhvLojnOi/B6zeD4WBIeeJxsL
PMwuHwXAaxY9KtoU39+z3aVTiH1T9L63h+TS3yNq5JW9+a2KKQMAdQq27T6SZ3Hw
cpNBxd6+AWafE9om0TV/C4ZFw2yTzciTrIL27FE2wNDrd8Bg04gVA2v7AWjiU1mM
MgiCVVG6InmHqK+j1gt2z5X8CzMN6XPAvLScnt0PGkZ8WJR/WobrEWlHikZ1mXG4
8sIum1R20IaP1rgXLRRVD920bC0TnjByrO5/PJsbga4XFzD0oiVQeMitZwd/7eNs
AA2T929GYRzTyBepX6SQP6A5J0EYfEsGzqGKUxC451y2BeJyBNF7zIy68IbG/rbh
XsraiE+fW09f71bp0+ComkIVZbdP+OVyFbX7w/YnaFS6HjFNeyGONSqEHCWPEgoC
mhV2CcpgXXcinFcNu72xhFhJrEJb6nXy9qVEBiGji/KibqQoR905bssDw+IftZig
fRfju/Y+ItfZVkgiKlphGFa8xcJqPzAIiq61eE9KgojPhxBpnThr7tFyXTsJ/9PT
E5vs/TK4iisvVQbkRM8e9t+HhYiPsx8AmfwjTgk20gLKxEzxcAFWzv3SC74Zgrku
2HGpHxKP1w90e9Z9z82XEdvSRwhURmrmZSI+me8wIR85nlmwOyDcjd0wwrRpFcpW
6LtcgjRdusq68D97ruYZ3AyzSu7ypFRpk+T//nFIw7j44XC1DSbhbXWiseCX/dNf
6B2H3ZPk3UzHouvI9xA0RrlbdgGe/LMOQpN+UXtJW8tKLgKyCmtRXtAuWFlTSgOG
kPUXOHR65JNWmAsI+Hxcg9o/VfTBUsMTPbgc0r10MmdivCYT3XkWSMrhPb3eFipe
KPBV8U1jV75PRwx4hjSUBOYvLtGDBBmUBgDZy4M0L5c08sdZTnxcIXKNhvqVHUlq
DQKJMM/ISgIsMcufLJ8I2TlrQWsVt7VGoSj72c6h9D/kyRUS55+EcX7wZdUjGTkS
Krllup4FCKh7zFu/MadPnaKOly6Vlt57Xc03ZTM190M8rcFfzXzBnryjv4aFH8Y+
sSOASXC+d1QoN7u4FZWBwxE+OQ4czkZm2K6XalO2REeM/6mUyTFFsC6Z0GvuOqwK
xIYhyYAsIRdgluGPr1RBP7rlBaR+aqUt8ImGrhVzHSvmdKFjzPh3tqQDVuw3DLfs
T/GLdAyEkSi6KUFf2A7RDdY3b9DqlajiY8flbxpGPQjLpumvMqztofOwVJWqQrM6
NBoq1NPkS6ctt3yjwP0AYxG7iipZ+EKcFHMJr0nLQqzZwfQKXOisAhkl+i+9D0SY
psoKWvOk9r4H+XfPNxdPUQzE8Jf57g0vT2QGh2hyNdxPtxBovxXs2IxkhlTKhWMR
qU9cWATxJj+yukZNsTSAlqd161QEDzuYSjCEqX95izmpRlZ5yzOVO6QtSDxyTwCY
IjsV18f72YqGzcABwkd+PHtpGRBF2tkbpMRNESgeANTDT5TFe582Um3oOOUplF2I
8fQRlF/g3I1SeGzt9UPMR+UYdiqXgmZdbqy9Ti5u7L75g7bJLofZ/SdgkvuIJX/p
QlNtGJEQGNhrQ2/ocZuojmWNzvgp2af0PBSMiYElxNUHPpe+vxQmE2H1TEVunmaT
gUiOZj/Q1aFFXs9R64K6o9Y6tnFBEstxjIJSqIZMOtiCw1l2QkWtAGqYKAoHJGFv
ue6oUgmIcXG3ai9fAaunI8iZyOUc9r5opBzB/jl8/RwLnzOjYanM/5mFEzQqGnh6
Hbf+BlYMFF+SsGfB7f2tyWmwlwjW9HwtUwj8TPfpvEm5CMwBc2tRWdFFlbKjezEc
dJijEwUfUOSQLiiZgBhTKsJyKNPXTzaTgd8AzoFBr9Ztw5nPW539hT4aV1SZPQUT
IGs9DMLCXlJutB1TEQ4nBraQnDtMuuNqYDOhr85PDNWj3Q9aoz3mBJvQTFRf8MJ3
Iv4chSHupHcEDXE9fuWnyE7eSU73UIRWcP3gbnYVGI2Skw+XFI7/8XCSVecJcPqv
d/uN+H9GTwyep4SSPVq3bY3wPJpzvKgGf9TwcBveh49Nelq1876lgPWzmIWw+63L
JfUk8H2ot1w+lJns3FawFUwCTEhc0dCl2LgR6p8iIrSC6ZDaXFubDoKofimTxvsn
0cJtfuAzj+8YBCFrZXH3CVPxY/4SmoTkvGxU064VQDfxOs2ZxWCO6Klu3XU4qrIS
iUwSNLGmfikHOHKNrgg0Y8fh40HblI/tRT3PpZjt0Z4BX0nUIvYVIp9CC31VwsIs
ZKt4IBY3X1DItwNwbHXqKq2jRXjilK6te7y+D3yzkinRIfTl0aJLtb4hdaw/zG9u
ANugWRRKLr7vFpSnhUuoYX5Nszz2jKjdP8Cc4eXjvgDiJpBEH3y34fdHLidBIeo2
JSDCA4hsmu6zXprJJJla9tZlDXfMQN3RI6H3GguToounEg1tJtlcLWGXbqd+rS1G
Az3Tr6Vo64rD4ttfXFmsHm9cXeYblsQhzOlGD+eY4AER8ROMlT66L5vAVGoerFKg
dW9lNq7ww08Vg1cwLp2cqEJVauxO4AnuUqtI0YomZE8IxmiEzNCm+K1K4khIXYCK
gPZoYDqzElWU5yb7HFlihPT4oQqBPgz5rm1G5GnmNU84EZ3Bokgei3vk8Akhdb/Q
mw8r6DCv5Sa+RNxv+FCak2SnRl+mbmLzPGa5PeKq2tpitBOkA4takE4TYHf9Wtww
6oO8iCMzlsHIQA/BEh9T7RVvafKPa42OmEP17M38p0pdeupp6z77aXQc43QO9PM4
a2uLKoJDvxJpBxyXcZ2IxEti9muQ2CzTgTDXACQpHvKe7AqkD39r3z0dw1vvWPaj
ZRoffSzWmTwpumM++FcQyk0PKOOQ6cJ98oG8wMWECaV1bPsVfj1hWd2IyNxyHkgU
YMHZdY2pTTVLsQkRihqo6U0K4XDOODWezLJXdgZqttY4DTUB0/vZCo4eoY8KQfGv
bFWbBWQBFvGwz1KvsimGjQ+24aDiQzRzuX8/l8cuTO+QhRPjDN9ZdVE7hVlgRwY5
hr7JjUwEE9uhwL8UQ0EShO36KN9ai6ldL7t2W2VEdvYr0mTeJ+YKC07Sj9jSPW2r
vxCGRN5uRiP7UVYyr8z3EkZwwXn1kQ6NZgxTr7a+MoLGNOjcj93sLI6zxiqG31NN
mUUZ7VzzdaWFHKI4FmGRIVdUN25H4nGh1AW0usrYnXbKWGHjUkeT6aZD+tjN/Xh5
G3zlQLQtFCsioCPFhQC8Tb3Cvhr1g0FvKLQjQrDTcxuYYcfxk2p1bX09r+kSdXrt
4BWEtxu3wMCp5YQPidFAhDo/d8PIrNxOxvUl5acCLbPf5XwyEIy1wq9ozZ4hvhpt
lHc5AYPklcVGmF45VSW28uUtp+lnUkoJBw6qcc2xpPtS0BUVIA6E9W/p1gNSFsIK
0b7/k8S9t2GEN5Xw3v3COiohRrJfAjCeCfg1+TeM03GJCtsNoHXI2v8o+SuRUQrH
68hA3hqqm/v/Mw5gnP42/6zR2BR4lXPBDYmiXi1aZKPojTWxbm1Yyn0RX9fr9l83
FL89c9ZNJ1Sjju7F0QmuwJB4mAFGapmVv+nQrQFUhYwBwmMFc5a0Ovn6KiCkpFW3
Z3Si0yVmORctK6Er5Vt1T+1f2zQdtW1fHgbgfb7Uls+o8IDuUInIkGEju8p9gORA
jnoqEZmt+/y2lViLJj3ozHO+KUvAKvCsvRY+T0t5Liu/mYKWX4SW9GPiGLkUpLGL
bBsVbBRuhJclYbKLTSGhd3aecjk+9hZ05AOOzrfQHPTFI1IJJBnHUs5UR2qNxiBU
LDK1oMCWVmiVP3YszGmrRR9gWHYh4k0j8AvJ/Z8lSmBbL3UXODdMRjuXHcED6Sxa
i6zlBE5qViZSOroRa+pnCgaOKtnbI1N7zOy4QpJOBCZ1xT80XypjLaqd9qAvG5hc
nfbLMDHKdrU3lbfaBM23uDPV3FbybTPlRx2NSHPld/Pj7I26mFODMg0S2fEV04b2
jO0KyY9Qa52Zam174Uz8IXd5I47kI5KDAjhe7dra3HIujlaKVGFW5xsCq5szo+IE
uyv5+1USxwSkBtoqcpXHNz8Wbu6x86g43v3cqaYVTMN2PYC3PAgqt9S1j6Kk+hRc
0g5Uf/p/hfGez4x5njIACBg3kROJAb24F4yDR1pv8rc7DNpeQaHO6rwOaWTxX/eZ
R2yI9DftERXVymC60RK5TmN+uPzsJQ84QQV+v/KLYW0xDF7JiD5gksIIeb0OeXwa
/XmMlhGS21dNORB9iifEDg7lWHDH8QwuB34+pjg54KnprfKlKpiG1vKTL1caNS/8
CDqiGrjUz21nLIKhP70dMGvOxwiyPLgJgHayDpRmrBOfSmitnNeH8zZkTsGd7o+t
3XLp0Kxdyrqv0DCSlevEm8EOHtQWPpZ4kNlazWsHA4zqkdX5zsndIgfDpjRsIXOC
qh3N8gefIyJLHznZBUJxFCpsHZYyHb8s2uPlaxcX+LvYijol6eQs7mT20UxHDr6V
J9pRKbSqEsJpXBZB2Ao7It3CvSnTLSPs9NW/HbxBt7PmsftWrcsLPS6kcEhQG+dg
iVOdwDLM4KD0fczfI1fijio5uVhAozWePkf6RS9eSaJAjgwGG5LqXdhH0MKo0ZWV
TlVPOCfFHqHXov25nHexnrfdJwLQyxvZhCAhsAKJU72P1qVryYS1cq5dvOsvrNVz
LN/2jouGp0RGm/4xUrRvG3VAhTaW2MU9PSvL+BqvpgafL9jwej6SFD14bAnVK5RZ
8Wa7wnUsItwAPCgTVLOhyLNmjX7/Vnw20fm4z+kmwd843S5w66EUkg5UGxWTNe6v
af3iX3HYopcsfdE9ayn7p31Virndyx232z7clBAttYXJ+dFfWhcHrM/Le5YVmFw/
sfOrHRYmem7JCA1PAz4fGKGFWCQoESUlgIGiJolHVMM2RkzR631qvZo0CPt7xKQC
rogwszYBd3vdO0rpMhvWDprXTYnqGuJbfM4tvjS0ZDU0Qlk5bhioURAi//U9ChRj
jR/3jNDvc0NzysQRSs7Oe4zWRW8+dj2C3U1irYSzwNvqDv9qdGri6Nrar+uzJk6E
e96dGyDJUBy3alyYhYT8mfp1jB92BqUFHJdcIXpeq+dwdcBm11ICpAev9YlBURMg
/VPQhmWCoW8saO+rbmwYFmFOAOJwcHw+KrycbF9VJkmAQbae5xtSC5hOiGbyXc0/
PRzOtOhUbuBdvmj7fJ+FN90kVOhoi58GxKVvCiosQvLc2u4bgfij8CYENuc33crD
EFhCqcGisj49xhJI5umeXtWEwRJ1dQtqyWzdYSl/Czw0Y1XekcjEF7VKy7Z42EnY
TFCK6aws++M/8krdTK7iaqmegfos4TOChDIt2KTKGoACtcZS+arocWHT5X3SmFyN
a0MVa6MG7SmlfVDm1TcYQiRnjcHVYx+7fCRg7vTSNkdsSfyX1R8+wRlcJpkBK0hr
CkxgNmVj3/GtqlZ/xa/BuanFtgCO+UDw6gizjyJdkXoIDT8LV6kBL7p4r0T/LX7H
dZNrCmsaVUIMGR4MqpDV+DWNYzCzD6F8Q8/5HPeKIrZJdklQKf4hhAnb7uFUgdfZ
DBbhmRp1tSVV27DFFRxFk11k5RMHsrsC66ckh1vWRaK2WBGWE8UMdWtQxrCRAyCQ
DxNH+B7lSbk8Gp396DxTtRiyzkMcZjYzpY0YxitA6LJFPx0I3hg26S6CJB3/iz63
pISPouXsHrOskfyGrFFGQyCQ8yD+8kH9z4+5A6hE9I70eRMvVJnhLtbX4PPB5mBl
lalLCw2Bf4aiw9WHyro0zb4M9nFmMjxMW8dNtWRhTo9SBmDS7b5N4G2OzbzhT4pO
LkRbzoCSc1LXGoPtMPSKuw+UWUhyZsvBe39FZh6RFAmlZwe8W8y28FC4rmxzDzhD
aXMqGztoN3QuBhC/zMLc/NgKl9Bt3sAZEjaVShnozkwKEvCOOENzXzWEv+Uiadjl
xyfWX9IUG4uI/GObDRCYcLe2XY02CmRHWS7RCGLWgxaVL7fUDY2jY1HRydLGBZ2Q
ixjCE8p3hEZ8zPXsugXiQ+uKf29+UcUfo+LHl+Sq/iHlECHO4Ihfa5CdEFbB0Ism
TOAJVFzRNJ218Xlt6zDsyqxmmS4+hHfKVrE1Q4478xQTqVu/2Yn3WWBvA7YgNn95
yv2v3kvwiihdRyGMLseh9aGaoqEZPT5Kw5ZL0eMRWSVDv36Dev2zDBsArO9Jz8gV
0XgqeUCA58u1RcMA/v2G33e7IS8aKeZDNWAxytGk3MGb5TRLd6PmpO6UWHkxqVxd
LsBFvjm8Xc1lG6iTi3TnHHCK6nxlUTrlC4XdBwhobQx42IwB333q7plJGoTSWo53
Fim8QBaMooKOyAOPVJjI4KuctyiELsB+4kXLjYnZSrQmk8N69wmVlIBq5XFWRS3A
lMzLVm1ZQi4GE3XMPy0qq81dFe9j7nfCTIJzNjRlAu+9JKWtVREsQoX1DY7tS6Ug
lFuF+ZjAF0LWBoRBQSHfRUVSE2ztoW1kw6RcZJgLiKfrgwKXhA3HxglNzQr+uo5X
VFYi8Y+Sa/sgUvFWQhImqsw0/IO2TJ14XUEtWFrVJ/LxASOs5Q03ClY3Hxmx00U3
gt8kGT2Ogij9jeY5USsCKNzvBw+32AeeOm6O9swWedNj65PYGo2e7FRPpN/FhzBo
HdZBV8ymq6mSIkQB3ouHjZPkTpSfbSJLQnxtHiiQRjwe6WYczhi2w81OZgrwGbS5
h+pZk+IeJQO3eVNqyuleZ+gxRjSr7hORoj8BBCd3WCQwTWnu8gg9m2R42fwY1hqZ
Hr9A6STgiEjlXMcyJzyFgny/EaH3I6SS74xuNdZVHXsiuG7rafoykad2AdvqZqi3
QiTNHpc29AbvB5OVAOzsXN98jSABWsLbuuAf5jdOewWzN7b3KMSLRm9R9+Q4e2Rw
Bw1oLJ2nC3dtjaszAmmrWLy1AyQZYDbMIamTMkH1cI4HQwSKTCZFE1UG6J0XMAlZ
sh08JGfS6oFK63NcTjXRKE4PlhspM7d+FfvlJgqWzSS0DAMFnpmyHBkTWq8dSa21
pJd7kQGgBeUhneILKcULIlItCRVxPeGkbtzPybI0i+Gkt1iVf+pK/xto9XCHza/U
wH7GE2lZsfqMtAFy5imlduLSm8+Imfz93pc6DSpznddBCYE31HVnymI9HwNikVmk
bx+gf1eyBjf1iongSRjkM0sAF2oGnOEh5iFVGQACWGvQsF2nAjP1KXJYplJELoD3
oNqo70OlY9EsvndhctRIm3u2WTouJWMxP9nhe+GKFgtb3IihTbFP3GwGB229G/Um
zJHjrfd4aU1Na2719vCNNOwLwnYNq+gzdwCmD/AoJXAx2dBV1fGCABzy4Kf4+GeM
mbEV7lyG/RouZ4tqWbqEayGC5D7egaPMBdI5ky6enygq/OKGXrFhmbvz8o88dPwv
IVnEAlKchzlr++AI/giXvsofDYlL76q5LA7j7C0RE2nNxVLNzRPo5l/e/Q3j+qRK
cwLQrcyugEywoYlNgXDDu9ZO2gRUDCFWSAJMxuBxzuEpN2Md+fJq2HYv/bLYi98A
ByOvbi2/OwogzzMKIn4cfDn0n8BZxTGuKr33yiEh4MpopZWh2dkKuCRjfYFlsevj
Uzre8hsjLsS66BIb4WkUvMJci02CppqdfEgfUAd/bDGonrap9wQujTfbSahqyzHY
NoZ6+zXD4NiIah7R61nvNSgxkuk6hHgBZ4ciANgvENjicSdXi7M5x7/1da6sWSdX
9QBvxW8h4FNhlCHQJ7x5eZLpA7XxnbE14M84eTAyPCCBROZJia5M4jMKl80cXSvR
pCtclmzWnACsO6ESlUZ5zpAJ5aw0SzuFQrSK12HYLmymh57WeaARSV4ogmBuDF7b
Xa6z5rVV88NE2TYjSTRHWbaWEZ6ki8izmrkU/s4kUxFnsiyQHdMqXt7WNZ6BdlhQ
VKPpM6zMM9umTzKpY0XrC6piCScMYq0w2WRXfaoqWc9seVH30PehEUki670GBNws
E/RxRBu29N/QxUX3B5w25bx4oGe6IZSsaI6IBHWpdm4wdSwjz5/ewJDUwXO723x7
W7OYrgVhAYh00wPXPVY+drxGrPgSOqfrjoirCq7OhaIf0G33hQkNRJAosZ+TH1mo
rjKwTHUJIMmEU11kZVlJepOobn10GDLMU3ontWCqmpn/6aCqj+mPxWPnjf9szWPJ
ZjEuZSPy1801WENlJtreKpFtXRBR3kmWIvNIAKSj1CmNc73xn9yC0sVlIc5LtyUU
hzWem+/R2k1E2c+qmnnXMu/LrnWvxjZWLHYHP6lmQSfKaISJ0C41ySRV9D0tLr3E
6Jo/w+bDf4Tgytkq63yEKSM13gpu0TL0nkjKFxwNmetu5OvRefXO0velF0EEOkfY
QR4729IYCdwpaJrN68+fVEg+wI0FeLn069S8wv/s4PuAR9kK4PDAqlVks6//eApw
ZZZ4hRdNZyEWfUuzBepmQvmXWHEAuHmHBTtUrs4wKljm+34hEDia3PRj2og++y2q
LtU2saip/bMkyjBMeMLBOkF4kHv9n7+pkR52/03zzPc3/PAvWdStG7D9mJM5a0Xv
S6F7W7gHIG8HXbZ6H/cNsK36fMCPhiLo/hfnw0C8FJrsZa0sH64eA+77N1k5795W
apGLBj45tbUbWsMkiOzJmTHji2dNwUEA6FnG2hXNWG4NHmRJwQWSa33txlDygFDD
iV1hU3RpzCm8xEzhOqTtrv1aG8HuZBfk+GNc/M/tHXdOXT3jJGY8iWlQ6RUC+aXl
sE118QzyCEQHA9i+w2TDjciCwpJ/xFKCyktBzVbv6ipFJIfXw1X9WIErfls65nkD
reW5MkfltRfoYuakS+q16PczHRo48QH0BYsZvRtAbx/0G4hGtx39XTjuGAXqc8MG
6GXwiB9Q5Wka/6ZTktPkTd2iFI2WV4lIvX54QH+zoa68Xga9RVr+MjzaMYMC7Cc5
bnFXhzA5cVCARnWkffY/aZI0Sv3aYkQdwBjW2SwWsK5p2Q0o1eyZS6OFtNxI2QXZ
AeVZggrt+0DB1w6RrhSBb89odCZqbYiegzs7Xd1t+KoVRB7JR5eceGfj60i+DtHl
ixJ+AZiq4vNlIQdhNSjqOZcIOIO0nKao3KLJGLWFAo/jOmQmW1ccPo/obDfYWfPX
BwqFmvKlcPUrnSGmqdPDd/fRyoM4QtOmr6hgbgPNGRxtBvfulAUT664iY08vGsNI
nNLL68bKGPE4NXhYOrKwS0GTrt+FmueMBQjm8cjFvn7s+0vUoDc1Eeo3VzS9+VO4
ipbdogMyu79N8CjRle9z2i9sK2uqLjw2V02a0eZkPTyLwYoIYm4wAzVph1uMZ08s
MR2wt5ehAuffQ4/Q9k0IXbO86uBRpwVMB4gobdudURDDkN19htf7CkHK4SY+oc+4
fdCdO/8w0dKK8B3u0eh+rv2wWIpr1chnf+8JRTtZ7/94VQi0vfEbb4yG6b9BxEMb
qQYB2HeBj4OYHvRxxKJQKsDiOYuoG9ujPtfLupT9Rx8xSW1dfX/rVDmhBA36ogbU
QewYjL2oBm/+eti4VznXoo6j+g6pLGwgk04TNDcurOx3eYDEa4xw5b1wbrX0g7Mc
RCfadu/mve5iMHeAkTKClzE2VqDTTG5LR2rJAycQ1ryTbtMU9MFdWfc8BiWWU36i
+SspXFwQi+BP/AYMtwUz+jl1rb/jnhDz1sJ56uLr25Jzv4+5fRS1IohCHJs+jfPl
aJUInWiO3MMojmMsh3rcvBrIwdfyWj5d77adqZ3r98gcI+WzZspNjTKQvZSvnzz1
HdX89N3gjipQLsNlc2mdwDduJ6opa2+EVSp2eUvA4lJpxwv99S4Vlnxh64+pBYUh
za4hFhMmYGawzpQpoMf/Mwi/AAA4+oGlkqTPhepBBtnc+l8Z1XoPXrlvnABnkYXm
1a00MEoepI2pHNofJJvps8bUpfPVXHWDQXCd4XeDn/Bmz+pAVjV+31DAH69HYpHi
Fy/4bYRVNj1yKlUdKZKrtsWop/cpsdSvj7ac3ERIQM+Iz0bxSUChYgv+vk+UX0LE
378gCzvZ76mxHg5eHLxhsX3714AWcEJRYn2v/bN4kc5DZmo5V0AE7GNw2/Jypkf1
5vp+r4ae7aFztEFIsnMIrOY7vJWESUNGgvYVO70pzwvem4OGdeHj5NI0GIh92YYU
q8/4/jhm3YD91GBcYWiaIzCE1rNMtocVVRHeVx9I1ZjQhMWS4jk6zcD7GoZuoY59
D4uxFPftCCLL0rD7UfzV6xZs/VZvUCV2+EsaIqYWz3sU6zw2NOABnZcuGe9S7dAx
CliIv7+zyEZwRQy+azKdSgLomdxXV+MELv3BuI2OI3DkRv6JvJs9jkFUT1q06RMS
aIOdolVzzIlnuV9VW4+dKHX4miJAf3K1rHStyR+KunQdNTf7gKwUYj3hMAQs0Bij
05PTFYSIgKqRSGxi0p4bk2fosq1uJ7XBv5/VRfSdaRfwrDxRgQ/7yjv9W+NiIk+T
etvpt1Nl542bfA3R52qcYK97Mdvf822A/suvZxfnD8HOCJZzll73y68FQJNeeFmn
I0+VO82jj0ft2kM8UkvFmeB2hNSuYID/+II4nSeP80LNpBrXCoIes1Q0f4vokycJ
mZFRUih7gS5GQkcQAVdgHOQDlWi2Cjg4xK4U70Kz0mR0AStW+tNKg2tqy/YbbF/v
S8ADpbTuSXeEg4V3YARyE0dau5ljRJdImbRVv7AobeMa0AaT1ZsHo7/5lc9FQvrm
yOCx9y9Lyr1N+EQv6SIoqsW/bJbdnW30/Hl2FBR7CRi5iO4dl8KSHPmg7CeQ/hy1
YxRG6/yrmdzBIamjrj8Bn/tUpqcOcsixMD9hOkdLCnpJW+rmn/OllYGXk+zKWNBn
j/4zNL2xjpu4qGMKVz+FEzJ9/bx/hpuZoVwAKXf5RTLkKMbRYeTB5ruAVz+BtdNj
Uf69n6QD/oFRY7sZGUEH2WWDhqMXeRbxNESaO3l/Z/jHQzEh3QoUbdURIDQuKk+H
06S1I+h4zymzWEwHnfo/0eNxHIy1qDhz0vCuwtLyORj7fNK1XgV/0HRgLh1v/gGH
qxT09qtenPTRXt5XpEYi1bYJRJhuSXzMGP9KDsa2LvDDsv1jmYD21r0xeIY++vgv
4H1WcTc0sYU2aK9v+CevzpBzDDY6lg8Ct4jSuJ9wyZrL8mjYeA0VoSnf0fhaEb3g
FOpT6vVyO48COd3t8FxFW/NjBOdTBlHsHo5gJa3phfF6NvrndCthEFNwWqaDFt2i
E/GObzCtXSTm06lqV/vl+wBH5aadKLxhWe80+u9Wykh2JYSm80rIW0O++B0NBnlS
hl31WgaYGsQZBRinPte51SkuuLELAnHEszSzaSPe6UhMQlzHx0/b1v34UJyR582P
xT3B68mylihNyDM2qfe9D7PtCCFrqKtZPrd07uScvLrk6mLCR1/Y3uYILU40DvL6
lgsyFJIqSUUDP6WS6eG4lCJiafnR6/C4A1AsRDHE+9VIqjxKQCjmD+8b16s64bV1
EMDZn6srpm7v2jkigUpXAXT/HwNXpdYbW14INb1bG2HQtzmNwnukhHkeu3970qe4
N8DX9TIO+fzOZDcjOwYDfST5Y3P6BW32RFQsWiyMuSfx4K926TtMAWs2tr66HE6f
GCNYiMgilNdmxsPszJ3VTV2K3yK0KhtEeSmq68JMSCi4aMVvL3CxVGbjuGBpWwsa
1lorYfRupX1zQo0jyEjZxnj0LMM+iLo1+qus2t0hwyxQo30/j4HBKOnHLJ6fqNT1
jzyr0cLJRxSL5z6qReq7h4FG5s/ZEPujQggIl+eu0ZrEvjV+40OQ+Du7y7Sqs38f
KuY5Zoj9pORgffHjgec6ARydKP0om2x2oRpjeo2w+VSj31WcAdbcjuw8p7tikqO2
EsxQ93rvtgXPJythYzJfILZmqiR5blYtv1tjP447ADyTdWKrmeSTa99T2rMviNtG
60+1PuTpzn8n2GeJCe9qEeIWjj7+trWdDvLu28bA8Y7taCJvj0k8ViCOv5jnB4Tm
65er5Y9IOrbOMG3TBImFnDQFNs1PRIFc0HqmjC3amm+rhXSraQshou9+hRasSMIo
cfXf/cZ2Mf5n8eRA3qVk1QtqoZdLloINtJEGmHAH75TrXdvmOGQcbdYWkd0BR2Gg
2jr1X97FunPyAIhzdKNKmiV+xXJAcLIrGk5OlPNkZqXe7od39xu+I0c6/y8vw5W+
Q211stpSa58muCkdCWV6pK0dcNV2A6D1ggFDuAbFH0aRJ090LpK6/CS+hTKyV+4l
1r49Nsfl0jUxjkNGMixYT50zOU74hF5aGYutnEChY5x8RlO1ZILAQft9rnccok5B
Sv53TwdiVI67+m98PZTVRpgcaQEXpMIl12m7frqZ0P43QLpQW6bc/RIYwmgpal0O
n/uyWyl70wRyAURxFKKLeOVrq8Y/ZGMfYHMhgNPSm0GvBZkwXy6GqdPHHOThe5y4
y3VyMZ+BgWFuA66rYzJVbFBLcQNOr+e66aNJiVXSYZqvozSOA4HkS2g3VRwn1Vgp
Rdr8xQZVkTdAuIFiLEXEgR9slCcpM8v/vId1/fvYoVmlB6MYXADegbCqYoj4o57J
+oYflAIp0dUVPWWDabhJU6Y+nWLFUiySHmBmSMqEkWeHveGumZtdB19irOZ/3gvI
AH1umDHPKAHDgohseh1sDItn6eMRW4I3G/RtnNNTcu+wUAwirIwgFH2kvmONGhQB
1hgXsPKfcfcDJKaEUBUas6IxfrXgRwPFxYF+vhJ1Tkh8pKi57dJcUFDvwUpTF6/R
CrlqBFthmNUszsMsMokJM11NAaa1/ZIXnD360rNVgZyYZBk80A9ODq6IF5Riccku
TxuHIk20+tx2mNeZuS6IJTl40k0wfFXVw6OkqAVfEuicHDQQtLa0wEIjhpXYueQ/
XimGIe9a+ybljbroC3AJO63pvsDSblJizNbcyEVj2lp7AoYi35DHxAEfodwA/bng
1eALoM272herAWbztZ9Eb9H1oPmMGkj4HkW22vzHHLOZ5oA1eV22nh2mgr7y6Eh7
YonDpjJyy1Kj1KeWTulNh7yvrnx+IpMdHn41tii9qgtr9/Vk/r617msIDqeO/h1s
KuAP6ztYA4oXAW0QbzYsqyn42VSt05MhBUYEl4EVh7aYHsc/l4A/WunqD7JUyh37
ZuZG1Dv+ZjSGfgTAVWEZNAug66IPACO5/6p+WvYwqlZlOOc85+o+eCnr/H4ALsxo
kzTohdpU5LIUx1bkOTgO/ET24YtNI23S2DrSxfHR9vEc9vfCgpDKCtpZkBhFm8qK
lvIXGqsRH3/TFNvSo1g6NL0hYeHx+IlMK8B0g7cGncu59ycbgUUfJ3gLaGQ2c6gg
W41U5J+FCoYGoDRfdfjqP9nA7tjQnNA7vgEH99UteiqcKV/3oBpz8a3ctMRDvzfB
CWQefvAsg57j4ojcH9kMat8wPXtR4fxufwNE3xQ2o6tAtvtidVookY+eMP2n0W9V
ZggB5WMu/p1NPvmpoRIAi1NDRkaCKgZBg5lsYplfCdHaXlToh76KAYBw9Kva6ZWc
ckec8g0Eppu06LZtFlIB/0w4sb7IivsW7yd2Uy/35wtFMGqXvFHAtYTeS9CahnGV
9A09J+yB6EHkldidlmdgAjyxaOqXke/6od9vQwGXxK9mh7JbrGOXSHPoD8lTKmiK
E12cms85lTP9dH8gPd8Cn9NxowEO8J4YrZDflcGDxMpPOd31yGV4lGvmh7BH8Dz4
/0Xdawvqz0+Kw9EY+7wW+uCTtHUKIgNzNsdIaf9cxGzW46PFbdqjhnRsluvyC83h
KxtIUZoNCXjCJaaM/yddpdf/e35xjDaRrccH7foGTb/rR4CCxL8H7n826FzGxNYU
CB6tossjyAcBhQ0OQTeuTGQ9idOVDeDOLGFocbRIb9ixvQ5CUSQdpQhk7j5xZlPc
SeSDQC4Qt4r/SIGSOtbDiobdbMYA/oV+HOIkId1/nKK17zdesSm2qgkPMaKUhdc5
Y8cHDM04Ntz0txIpU0wx0DZFyaw2zMHbM+jLHszCxVnM9/j+PFFz1PeTO2thl19H
sLHgfVWb460pirr6nzJBLLaNcwHpSrJI92HASQCxF3Dgui0RNSVHwbvE1Fi1M0fo
ZX7NM+ZIwx7flvHOQ13jochHAubfWQ87YDig+H36YdOq/pzn7RaTyqDXAWvFKHQ1
HOuVTzaz82rcdHepbjBIkDjiSfSltFCon7fwe5VZ5Sc/7PUI9Sctof78nmdbcu/s
eKTejFAkCYoub6kSNR5gmGkaXXRkQjXcCpzeKZ9ArfM38DZc5pkTlh5EqJnhYBkU
CE1BvrWxeudZSSh9ntIqN28YDvjMIPkEIA+nLAfC9xfD1zFFJ9+GKI3s/PInstki
crPPSp0pac0O3J0ecWFyDnhTPTRQ0LNBFCFRDQgrIDK5RPDhrZFnWeZ67K1WpWQI
HgHoyidNFk0RDdA5GeX4GU8c2zKYCp65Spnw0vRck0Ps7okJIf1VjT1FluCQI3ou
XGdMtmqwKir+SZ65nE1Q8+p1b8DyRHRt6aB++V1HFJAOv4WETjLElp6R4HNrTrNR
QaRMLRmQ3xGluBjqOCHlPeEZLaFCm10IIcuHomUlPEl9LrQ5CVVzp3XIRxJHjYTk
pdLDQWDqXVtAWyuo00BxXgCWbw2AFgjGa9IhPQSrkrkcq96J+wTFHpbR+Mrbdigy
YTqR9Sa6LkE+6CSZYZj4VHp2tTEBQeTcueqNCUKTXS6XiNWX0dV4jRet6rPDzK7x
j36gr4cgPReiMdgZ68oSKmz0UyaKhvD/5cYa8DnMf8PPe79ABc/hXNjntf9oXPUS
zKouEwA/HhYGArcg+0XW4KUYS4NbJinQ+UDTiKmGx20qHt0LgBkw74/z4U96sUZD
KQy5QmK7zl0ShRg70Zk1VTejRUwKPm2z92nQbytdCA/ezwvPeFGT7pMgYn5IyOLO
ioafKjGrAJolhHaWz9z8VW8dOJPWH4zDD6AD41S9+mufCo7IpMwv81CQxbXOeadK
Rtw5wzLuXKe61pCL+z0Wc8yuvmWsZ9ja8xg33AIIE5TLfcQMl+S3IyHopQVa3gqh
GMppkNf3HoQxMyaZGP7/KhbJhYOYow/lwzj2tgTnY1U6oviWCSS3VrDrrNiVy9JG
f/wp3eQtAzfw+8dbZ8BbRlA6iS37BdP+qzIQOAMoWY6mDwy+ct54SGs8RqhbJAgv
9VxEA4lIpl4KDUK1Te73NnfwgnBtLxEWRcJRKil0duyk5oRiUhYz18hkf5YtqC1V
09I+Yden4URRQPiS9vWqsjiXyAAQbp7sB3eM+aHZeacsuczRkGswD+RBF+f3Ph00
2j1uEgMhQrl+nV7la4aNROpG04pItOEZDWWn8Ul7d9Y1f2wPP4+8MGx7w5OsxSIo
jIu+Atlk6aERVy/9w6j1SSZG2JA3TebRbB0rEM0mKuIGheGHdhhLR1zQIYy2IMKq
k8Db6m/1Sq9rCU/rOpkZX80+9Umgz/MTv4ixdijkwPU22qEaknzgYrCy58LFh5Xc
LCGVGZ6uCe4vufgElDlFpvURbXwMlGAyGIqHZqq3YvFZa7F/U5/oKcaZJgOlSSgn
gKefVSbWbSIDeQu4m9/rNkdNzfdO+VZSjeUZA+fLGiQb01sF1yRF6Cwyg0uvvdbu
ukTwtK8xd8Y8gujBUveg+pp3HRwxo9WqrWphwyRL72h/vrI/GuA2IFQhn+5UWwLc
UDos6QRVZema58HC5folU7qAYLYlwzSz44DbylDPieSVRP8gTHjnHz15feQVUxAx
dIJoPkNhmcTu0v+IHI66Yyy1bmSNpu8SjJRppA6ixPwOSNJz+55xcFXe3CINAafZ
XHLGAzNPfxrImV/GsUDAHPmMzKjPym3Zo9Rj74AijelzWxpUbwCqt0ZysZP1Msgv
hS/avxXG96gmS70WQXCJJ0k3U8ADNVsNRS6xRDLD+QM32EiIEbU9gJmg2OjCpdyk
Y8VpAksYJE500YlV3ECcfVhO4CD34GNnRTfYNWKrTw9cByd59wQ3Tpz0olRnzJ4H
hwZYyBpjwiM3d6Ho/XmQtHtNfqJJ/L7a6Ed1HtHWfZgyT3hsFrr2Bjn1nJ43CUVw
8/wiWGLvTCNKJQRo1ma+62nb9I6wnQ1Xn+RkgoVPGWF/klzHfwUt/5p4b2B1CUOr
V07P6M50GQb3V0kqpo0CwwzN2Iqinf63jMmocGR8LxNDi0ApbIwUEQmyKerPznpH
KQF/HIDy0yz8dY06Q6nrp7dR83AGXSHeeddunQ1zh7DUl1gO21+zs/9ur/aRhnLi
KmFD0jZri9ha7AJR5xTcN1af7C9teqM9h/C2sgmVagEol0ZKgOUdlxLQaArEUaWN
yR4nK+irJDVGQPPVzxiI2mj2EJuz7gIntnasxOGItqJWAM8wLR+caR8HDIIehwPk
e7AZZZg6+DTfZvzNr/cEgTG275aIWE2K38vYSUWYpjCrRMcmcK/nLcNmZyH8aKCn
dHGLPwYreprqGUI3+CeBb071dfoe+oFyD6dCfYn1LK3IeXE40L+nDT9EzBO/L/az
VuyGu96PCvXvhM717xXeToFGv+8Gm+VBe2wJYpyHuzvHC4sTKQBjMmmSDyQ91wKN
FEwK1ZKDBR79fwROOH6e3sZ8NjoZD8L9eAbqXkl1WJgxgo8TWSpQdALybXbS/9R6
dboUdlOEeY48HiZE3KjBiWQ3tl0zZTujDgEvnx9Dfazpf7ZW5EkGtDHxwYfSbyr/
Ll2a6c/NLqCp4b5w5W9T3vg6gZ9MCeI/Fwubb+g6jgV6jpmIa9dZtF9w+/wumDQl
ysjTQLNYeCvuRQREOCkV7knWBVXN/EdKzRbktwBoNvJGb3e0FA5KjvlAE5bLoE+K
yBId0W8n0RZW5dtYPcdgt+8J1yxywJA0PKOoej+HYvUh4gbpawmpuML5vyHYSM+G
0zO52QwPRVL8oxqy06tdUyBmje6y7EDWSaSnbLWVnKo/YWbdtlFgt6fSsfbgSLmv
XyDgT5Io7gweBkm+RL6jqkHJxCwIsA2iHh9Zx3S+xDQnfyt4Z9jmm9ByMw/7/PGf
94bInhsArQBld0qo+CAj+tN2y3Q4TjY10hQxQeMmqbNRc713YY5ENYzBqx5vsepE
rWC+gax8L/JRWPLM95oV54seHtKFqRGz8LCD0aO/HJEP8epmkA66xsXNsisdhYd+
vzh1m5pyN8pqvdReslvCyOUI8DSnannrIpath9qzr42gphUtlsuryABaEMwq1h0v
/4yHH7YbJjTzo4NHPxmRwc6de7Rw+Z+K0VYL7I1uM1wjdeL4bdR0dvaQLS4HMuVf
M9/GXiaqs6bnSSoLHE7t455A8GBpKsMHQ8e04unM7QAKl3SYJ05oCtOvb0wDg0IY
LK77lxaZctgnPshSGG6wabrWNZ9wPvBGUKqzbHI6+6X1rQxNp6iqN8AngdlW+lga
sfZpGTOcUGavW3IWbDX8RGDETU8pDq4s/7BVK1XSlUAAIeqRJdlnRtr6SJqkQgAh
oTNeTAXnGIC726q6Y5EyMeA8EM9COsjWqeNuQlqwCqpe81pOmGILq2Y6HSvn8ZJl
fmuS9PlRSAm/BMGazBUa4K+45YOpAc+rMI0mT8fJyhzzNx9rE4eOSQ2r4lOXSCyn
goXNsjRa9WAsyRdXtkOhQ2X52Y8VLYay8emKbfiIDbyY8eIhaU8RXz4/pzsejBzf
vKdD3zhl78x5HN6nkxYFKm3FCxEM50keEFFXYVwMJ6qq+o8/a3GXeyLK9+Ue6Dc5
ZvBeN/pKsZUlq/1tqcgUSmfON8ONg08T7kCn4cABkzPaFgG9x/cOg2kOC2ofgmlR
hZKREH+VmZ7lgRegTWvH3iJa216kXHw0v6xpAt0AY+RiK4u1vx6+JWC3vxJO1sop
0aDuJmEUQntIX/T3w66NnksoAMPWN1PQUY+O3tGpxRRsMeSz3UJd3YWUiGwEfzpH
+n6aM66LsFkD4dnOX/dyUx7PsAOFPIp40Lcr3WN20mvyE6Z090CPZ12UVVLy/HkB
Q9FRRnZGAqUyEL3sAbzXn2KjpWfrSyoGBJPo7891o27PzUpJXTTLxlGg9DbrtIr8
IWYdTWDSMUamNIL2dLpG40fvIdeEKb0dzUmttcehTF5vlUYg9SU29t11e8+Jb52D
E5zMqOkJRYuwQL6892DCqgpIW0rmtRVv/pd4qzWC9v7l2IxheFYIwZN9p3cWbcFe
XFmi0EwYAXjsGbdFd2PfSMF5KmyIomwRnkaZC1bTa95xjbkqFD3ppheCcghVTMdq
tyC/d2wGV9iKIFCeZgKvRfjGSadJxuPe1ha83MywDMKBHDinPWSapgKM6BiZGSN2
Xi11WaIEDvgSMj/xZmS2QGk/Q5ppUlRCxKU1VUm+bPCgA0iXhLhnkc3fLoStKpX4
eaPq/RiiAF9EKGyw/X+JeBtFkoHUq66brznDcjobUDn2h4Wh/4KLBh3fVLXq+Fbw
WA9+pgDI5/ZiNAujCuUXcEHI7YNyyP44Xm+f3MM/Kopj7lXzZHyp/pdWyJMmXOgH
VCJ/RehL7PM6WrtUygNIJ9JhZ0R+6AGvwbDSwmhMDLAAVsQO6/Vb9hce8KBxw88l
wr91bHY3o/kR5oaZ9oxB86OIEbAtSsJEdNbug8cND8+Mm6QO76iCuVGI30Ab9Cpj
3xfvYLwIIYL1C8kd8AUrd5zrpxkPtKqnnnuWkWnFBVcihIuNyq9v2xPlg5hfDMx6
WOFGofioGle9NsXXm80qYmjAeS9YeOTqRC/fnwJfML/3/unG8oFRihUjmWuYlKR3
aTk9aBhgavhQh2NxyW7kG73lkaq0J+OcqngxJRo/veU+ha1urKA0cC6mzLoFRzCG
L84MrSEMOWsUwI29dKHrsNzP3+dMw3/RxdtNsYj1PaxJkhqdmAaumCGNFbcmkHAy
CIIhCHNXLWUUqtFrAVGV7bldMgo+T9w/P7rOtjDF/UbKPlDAaxhFcEoGqzjMCS77
QFbM8LHoyLndFWxPJWEqTPGOBPMird20wXE//fZp1bpmWV03ngI8KliuylZY0uGu
2IX1CtnXzQmpusvZHyVXxq9ote0L8eg9Kd5LbHRBeJ5L857R6x2OOZ85mmcpI+KH
Y0IGk6hrW/StQt7nb37M1/rFNspHdkeD2JqbCKH8EpJK25YDk0dXrs1SL7yzN8hz
AyNA4LHOX77pbvbFyFAT4EJm+cun3p+qo2GPz3gfizw5jTH76UNDEvPoJouYAD+V
sYN9ZYHF0Zt2mhDwAIIVfdCSFSh/IMWpG+i7MncbHYtLH8926utG8EL560Lk09/J
LUxFpweeaypaDh4IfFDNN38hIc6QJrvRcRvlUuFR88sWh3BOHYhtK8ezl8mb87pC
Gep2tyuup2zqVPYYEvoYR2q7daWnw4/joxSsMpGpD+5vEk/r6MAbYtcta65TUShC
5t2krQLM2G7kAQpfbm3lsIeWXIbZCresCqLhQHwVo7ItzzP3cYyCPuFPBbqeUNI/
r+/dmtQJ+8zdzq/eAw3cckslo6iPTpKKfbaSAJ5IgZSizUptmswSjo6G9fllmqY0
X573qxgeiq1IfKojn0cLcx6cL13Jlar+VDzmXwuw0kf09ztaB3xEFM0wpmiXdVSR
2noSWpcXSmSl5J/cTrpkUJvn195wolHgTTXlYy03Q36PbqyJ7rZStRYK8cKkX4LG
QdFOT0F8Pe7X7KVMga2V3PVXmtkYrArDK9H5vDdcdlaBiqrPU2FWayJlCosrJN7c
CJdXuC+QbrgfofuSIhwKVHIu7EQGldMbXrr6RBGjF1OXmyopRqrTgzJlkBIUimYT
jHI8TLUyrBoZWEVQVzexrbd9QnlnyaMu94+nhPzAufhOFO2VSaZ0LsM2mPKOf6PB
WJIDdZiNC1S6JgOa5b/bNhdojPgrifxnzsrtARKleqBW5cluH+gm5hkRb2Dqx8BF
Vdm3vArnVr3V29vrhxJPCV6pfrXjDvg5dfTFER0NFdIC1MloLzkAwC7bVBCY4y+O
KMD40xiJE98DKeIz4yF5PScC78d2xLrWYMivgM97Xb5ms6Uvp0uubZnTepNx/qRp
ayGF22xX+NktjuAcLKhNBgIZXCgbn4PxR2HoxelxhdQWxWdrVZhxFqzrUWLPjTWD
MRuAQVN/nVmzrukA2DY7ShZnyA6n6SbDKJJPoxxMchdvlJY1KNDATZXjfSILRJsJ
2IdYlh1T2bPvn2jkXR/MujMl0x+Z8QPrj3/Jv2V9reiY7Maacy86cC+GRGhIwxTR
Y0cDUpHZrXvncIbm0ZF38hs6iKPzay4NIS/ht2XPlnwkWOm8T2gw6zbdUiT8hwHy
2fEQhe75kdnygLwpkoRMcgguY9fTPvZaHT9hiD+kERM294ekJPgP0tp0EQGzj5VM
Ww89BlgOHF1LZefoGnsbsnZdokg/j8ZJc3NpAEMrh00n7+8x+DkUZD/35GHURW0g
6uZEBM4vxc96orIIyspNt50DuzID0JYPU7fSSLMkFKY1kA6MlCxzYXW3dWaAqg/s
VdyEpdtjDgZqCdj+EdWKb2/a3M/qBbCqqEFjlOXVVjkryEjWskwW+4eA7h+YRocw
XqEntT91tbx3bQWuohvxBh6omOWDRLHMfRPtyKPW1oQpS77tKg0/h1j4Odpq8kri
CLzV1SrOJzYS8qJyCiS0c8Ur7/m/51Y6WJyfyMcSV3yEVJZeBVPEjAKey7cgf4pR
GQta8ArOTj5OkB055IABeO4H335wOz5lXQIvoJPmaJL59paYKFms8iswTqMUkexk
ny5ePCOCGHehphBoHJ7EmcFiDx2OIyY5JmDTnKfaYRQ15k4B1++5D1cp6/vQHR3P
x6DSCmM8QRYkZ0TdWhzhVJAvNvu2RF9PW7daN7JcJxZ4m9h2AY6cKYJBsYgGrqLZ
CcGEchPtMx0Y+Suf9RHd36W6bx6UZqb3mOEWxMI+pTApocCQ/DBpO+oXApaGyUSB
3f/ZsxrmpzjxbUJ+o+ddNA9zUbQ93jw4ilCSVpUL0ARtgasP2crWFWvPzSh0SbZP
3doFMvYtKhdgb6VQvqANxpHXy2Y2oJm1UY2rf3EhOFpW1uIwX/cYm9PAPWQzIuoM
yw6sMYiZS5DYIkAg68btnpm3N7uG5pJoOADjuKmrTm67moDSkMrGMA9pvTTzqeyG
hHcmjPzFQ9QHaKNLeMbu32pcEW1ofC/jXmV+w7E+3oLkwYYhf+rkW7MYtrgrSp4M
TXKxu/yuHqjyYKA00RpQgsUZnDiyghlj13FfL2fQVuzjlqUAKp8wzCO6wRPeWwxd
Q+DLyEHWqTXmjXlmafCsv/IrajoYzf3+3L7UPo2tSyiHl5ThCAwB6GJYLb+XCG6k
TXsCM1F27FOL2DPLJ60Q1yy8yKyhb85p9fFMKw9asA2+5NAquJR99550RefNAOxD
TaFsd1lm7OS3sNe8vGTS9F8Ru2BcrPcEhGg32YbM09humZs7o8kkMGyehxo1tHsr
MoRzsnt2sN6dHVYO2z2xFrBea+9CIdDVUfVVBOWbOWYhbS9b9GnVoIsD0JoP+iWb
LPt+D/953R0wc85wkkxrvR18P/wr6/FrgKx9GsJOSLw4ObxXPhvX6SV/XNW+HfzZ
gqLqaG9HneGbvE0tbsMoidhV66rR9I/ZEoPcLndGx7p/T4vE3Fq+G/18JjChOYyl
oK/pnXp0KMflwUv/ZVkOMx07LA0jePxsqOcIqkrnWFkjROQP1mMZFQrLo5sfCgqR
mPrPkCfIr06oDNgoYTcX0y6wWh7HstKU+SJiLIclwkwEecmp6fPv4RKgiZwW8F1/
LEKCnqqNz64/GkJVcwS5HlzCmpxk5jOnqu7y2qgt5PEzi4B1K/1q+2DpfL/pwoM9
VjcOoAjdfodfHfhjR3FSHfWEyHnIjaKvfS2GD9Aw7W8/iC9pOsMjHYIniwqq+OEj
fRVwGhDilmniBhBLIfqv/ZSA3w5yVyj9ebk2jR9DIzabP1bDsa8MbGgTeFRD3Hc9
TzaaMGv4QYiM8BP/pmaJY0bxYAXfGu8QIl5I5+mImxU72USH0j+n+vrmvL63lE7e
6fns1BBETH/iGJOv53ygAnS3BJXJCEslgS0+1SjhVpM1VV80UHG8cVaB50eRr9TN
1up39ORoWYOkdNL+LVEaCefICpi1bXTfzrr80jy91+EfUlC2DGQbMNZN0LDeX+xD
TsJpMAt2smZtvE4GXf5rrj+0CWGYdjNVXZZsZrva70W7/UXoCqyKb3niJx6Dbeop
PTbNMEodSUarvl9BXn0ndoOIgOf8QwrjUya+c8QAZ0UGtNYghGtKhU/9fgIkP+ve
RKlqUKGVJnGGL/4xBBpUwukduhOeufaCrUDDDPqg1/LE+7cwNNkqwVBmrEJbOoYO
nN0hV0TQmwAiAJ5mF7jIhcNxVtYhxGdA+e3A2giPZ7KoFHTgSmexeKYoEBQT9mv+
fLOj2kspbxyu9Jhq+3gF5JYhc2tFfnAaCEnknOier5T1BMC2mhgaZmf5vO+5v/Ew
5B4+cQoWJVhfrdJly12WHFkEl+jZILvX9cfNro1MGSpsrcXvUQzUoQRQocY7va0A
PJg2y2JQuYqNfGok38OethG2FlOTaOe1V4O79SZzQDT2PVQ216tPF+9eF0kYrGS3
nqGvd1Dz8QEyQv4WarywJKZTUcgNUDp2t7M/3cfhglqLICgq5/IVKelfDVyxqfsi
CYTLrZpmtq3IlS9+2pFdhOU/hYxzkOIDsRpFzI9/6nmSitSc4uHwS7PQDcTU1rcI
wPo3cXKgJVoHuXNRpgZzzFc3OYH1ZbgyEHVq6ZnD2EWb5nWKkRG67y9acldk0196
nN8C9ORY9EXXw6m9vnNqi1AfyIoTwroQ422XoiIN8GgP4f9FPzOIAftLeOtlwA5F
O90PDHA0t7YBmEebn34P6HJW+iPlyDJ6llbys9RFyhTIkXfL5JjOAW960HRWNVih
kLLRNvhhYLiZAM/ezKYTgPjufrEooGLqrgJ5g8czDTPXAWlKJky0EyFOkD1KdT/w
pjF+TrNfNw+s2CqvRTxFMgtYF0JoVcQZRmhTlx5qo+OyWLcEbAOjB/1ZxBB44I2Q
Idsd7yse7DUa1EeZaz8aCHUiDZJFU44HxhQg25wk3SCx97lPDzmQFsuUIqayBgbM
H40D2Pt+uC9CaZgIW2HpC6A8ADlGHMvVssi67OyyJPVsYuycpBjNGqmgcACXCBtC
jSqdVjOW0bKQVO3cODej+U6hVcoc/EzvxraK59DyY5WZfc2qK9MilIztdWF2+Sml
+4YH/6PTMFWu+OGrdTl0WldZalCULG5w3Tb+A4/dh6DVv+pH6wDA1a8AXXo0bfB5
EkHw+9n2DJIJGOdad8X8OTQGbBAkBGSdNMA6x/geDYvEcSSaK7/J4i8xMDoUIkTE
G0TkD/fX7NbBt862hKQeF9lAFSVUXqZU00rFRTHtT3q2z4Nfd/RWu2HToZPpn2+R
gbbHyhIkvpbXQTFB931jWimJJCRWr2yxZlRANn3d4cCQkB56mH+pWR154dzHt0HQ
qpsiV8+ulQcOcgiRCNwcz9izeloNiJSICARVqS5nkE5RrmURFI31ZQPfOu3yVF90
8sdRYx/CAn+8Zzb4nvcMwCNKkFJbtIL+JmseGca/jLMMfyXzMxVe4xMlHMOCduMT
k9pT7FacR3IM9//cfLfuWCo5khnTAYGsCtsDt+6/9xx+MatLQY34N/cX834YsqI7
L+gXI1qx9FioQrUH3iHik7Lq9tu/bj1pfhST75BTuHPuRShIMvkTlsa3Nj7Lumd7
ap8gsBjejPslqGYdGByBFmSir/23JkCoGMU/GgUwsswwuA5Hdz2TcuY2euk9qYjL
OwQjPq3tlej4eIBwnL6f9GaAfN/2rc/BGPa4Nk4FxrGUiEaIzmS/hnKTQM1gK9p1
Zyq0S1zCByLgTHq0k835v5wnZFzr4w3gAItkJQPd2yyy3123OcCQuxon006AK3nn
VqxYd/wEMCQzPdKmKGMING9sc93SLdK0ckYGj3OoT+qz9AlvyVpYh1O3mIYQcCXF
gB6jejsdSSF8rkC7wlKJLPWfkOCOQ6ITHbw7R18L1SfM5/r7UVNLZn3N4LP0t2eE
0SQXs6A0e+hZ+pg/RW/6+40jICZo9PRtKDq6NrNbMsVvb6TXU2T65H26ux406+WU
KdU4ihUN6/uM+8SKJp++xkOb8Sgb7cQuKPSlUi7dvW4FndM43BeaOpfILJify8AJ
DyExvN40OXOKoluA+FHGBJUWzAJBoiBbdn+JL30pnDZv5ABo+rMCcPciwAMxaq61
ssg6Jr2gQD03/LCbYnJ9qI1Rf21hPQN0hlA4JZdCUVz6Q5yh90SEUX3sdDbI/xb4
Pef1FBtQQgdcEnc4sBNxXn9/W1sVFRcjzZiPcINFgWFJCZ7t/nQ+D7JqT7wd2PJH
5W9c8HMXW2d6hd7h6WdIArh3KLXG88gpkFed35qguaKFARvt4QV8amjoogzLd8Em
SMC/cf5SM3zOW0pjvBMUlyWEdnkZ8GmjU967eNus9EuXb+wJ0e947HQo0SzT+VXc
w/1UjoNJ/zdNr75IQvzi6ROrJMGsMQPmfhdoU8lCYKoEh8nRQxGwP2jVvLAm37HH
16/yo/09TacH0MShyXPGOSuBaDYhlLuZ7oNZtVSd3y78xiInMkmmSB6cbklGURpl
tT/W8crjaeQnv671ua1VVuvVWndAHbVfwZTgle5AkSWZ6ibyHgzYh8sKhKmajcxs
7EjHsT+53Lk1Ksgi3lpsyNKo67krpIml3CBUcK5hzlzskjBY/tUf7pknpqs6zkI5
hfTVUR6/330xghtvhGKtOcQ5wBnq0TyDGeOWtBU1LoDoJ0D09fydYyAI7cN7OYk9
6hwfsqz4Pr7t71xqiZaxa9KzPj8FaIqXbnx5L4wIlL2wbUntF9AUT9G1XpUZ3k4t
dgX3WwK6kYMYKxJFLuFeMEzp1eV/cu31iaU79RNL+lsQnSxYrxoA+GcaQedgfOJ+
0aRsC7GGs+3L49y820pQHsqPlC/SXFHPDLL6ft0oZ6iDmXuLB+SBpNmT4JquyWfO
O1s7sPZlncaMppC0qIfolvGHm6ebE7DPoj6oXuudUXQm+OUdAvaj65UgQL/aEkci
dopln50CC9tyP4o+kXVECSnwgKaMdSMMa+YDoXnpwMgLPdmv+k7ItcQ/I/8dUe4M
NOMV5snU9iFaytewUmALPsyrvp9iDiUh7Leho9SWXE8s//BCriUmRo8HLJEr/tTb
oORm2aarPR/QPxEx4/v2/FNJI+Y7t5MbRYBX35hBi3zHV0thdaav+hUHH93wG2ZU
exmSiQ5cfHD7p6vUu1tfCmUbjHeLr8vTlGlWcCA/T1kjqEqbW+FdL1D6T22pylqr
wVPbThvk1t9qJXUENIIj+de+SIHk6UBzXBIdAeWmwd7B3u+vJ5VjcYUf/8DYvcKT
HMR0bYLH5B6LN3tW4qoSAW38oLMbuQ5Es2lgS4CdDUkulAkXxdaQex6QYyRTQC4e
+X7xOlFDm7nLhqyB0d2BmUiQk2xFXmbx02P+ErgRmCgKHIG00kUSmIp49c3euWYf
rt1XM4LJIk++fE3cVAV5/g1AAjQIi4P+A3JZ//unh33hXUAQi+L9GgSB7lCAU2R6
sKwZNy2k5yEwG1dJX+wLNJxNRKAJ39N0blWrkzeP7unp2NpGN5bpT4nh0fOgUJGk
PQUjxcaoTOo/mZPDAsxWg67CJG3m+pV1ak896sJRGcGpCtkX4sGeOlolElmKyk/6
FFURNwJOvzmFujgU+M7Gs29iumBWyYu8eRKnEjllB97mHD+jwfa/Kb9KMn46Owyr
ICH8BcH0DzHn5UpvA8x+hbCDJZnfkXLlAg9XzpxqnCB4iXFdShGKVCDtc6soM4Hb
sgq98LTOlUjtuSEwQgqiYeey+cNNCimnnyYApuKSCVn5QwImwvrLhBtROAEqaLaf
W+W6bfC9cY5frm84/N/v2QWX2AN9WraCxn2jxDgfaK82c50CGYmUi8gw3U1sAC1N
SjRoxILj2LVU/rXxHktPFVeHnedeS7U09khJew1MUPBi4KFTjD1GeFkYU/zmuD7v
ug1HcdwtwEDBqVs1BTLQRtAhHqZKms1PwTmSYQR9a8K0+2AzLCZTm8rfnlMOe6iP
0JaicWoCfGk8+XC+lcWDADwaqUUZVKTIKcr43oy89xjPj3Mw5e+0gtDzHNJptbqI
WOCPshUD7uj6JRNoEIlGF/1w31Fi2HCMFeIai7jApRb9P3DTgeunSGBgk5RklxB6
yqNEIfYiVkmkYuv6nb69QH5JIWEnZoM9iirK81qUP2YxCXLTILTMY1k5UK+HsFmq
S36bOzKIWSABt13/F/qzu3ic/YZdK8Ax7VQ8rdxIxYz9LdN3xJ+JkaRtaeZeHSWK
cgXrWdmdMnuqtwSzua8Sw9qzER1y2haCZfmflr49+yCmFkkvKQyQl0dC/9T3ffMp
IQWhQp+QaywTlJ0N1t/DCYHOc3q05/Nh9ZQkmtFmKzGpCUb1uLsqsb7cSYZXAlL9
TbeB/TOSJAg27CvZqnHFc67p6h27hO9DM7OLGOze7q0nb5c5fQ7so12PRMzNlqZ5
yVg91+5Kv6m1rkqjU5nZ6NJ/CUF0LtuTNllg6bEEyES9oxP//yt7g5+LJefnShzM
z1+KU/NkT2JawZGlkb0ubUNTZoIM383N/HB6sIDi/vu1qL2SNkkakR4+grRql4ZZ
Yuy/X/zJiauoiCvFrY8WPOwBjFkMrj6ePbYnSf9WP08edWyRmArc7XWkXrC06JhK
2O0LnzIQ6YrcW8OR3opeTNY3s4ie20r9XrwyR6Bl/aQqRDu9m3gv1nF4QhbGqO1K
mvwOVfLDHK4jevj3dVS/AWfKyPpamd5Sqk6+p0hRXNhNTbuJHLnFjDkJ1PdgC+5n
nMq5NzQhif5tsrfbwGwavYcMKCTSpkTSiknebDbTawFG4mNsh99YIUnylmhXaF9S
m1T+N6cNZ2CIbNDCFDuZK1ctoid01yJS2yDcK3t29KpJCikk5t1qkGb/nLnNivfF
aGwlv43hCSesQBmvyyrRKdFFENuNgDHpcbV8pqysDU2kKI3QdeZnUrkw8D5RFuDw
Pm54h5TtdVVt8HwXx77ZGZKNwY58pXhLJtcd6X8IodWzz01Hh72huWm+OhfJkdK6
OlvO+lawbOvGmubgebmu8HTumeqlgws9Mo8Yu/bD4R8PwmWZtq8jWIGafYD1Pz7z
vlheZ/xT497BLR6jW2sKbwLM7UtxMYTHP4sWQ52voVLyhzAry60gLQTKo/w5n9kq
14aWztyHg8sfCTxeqV4Xcnv7BX7X9wpkPivofq1UfD7EzHn+KHy5TVphWMnvoyfP
ok/fM0D8+qCcrULHHnrbjV6gplbusg+CiIsINs8oj8HEdGB0v/mU3a7+LH9wGxFR
ez8NZTafDZ0oNU/raV3Ilm6yYkjx1mr+YwYYR9nJoFOmKDc6rLYx6GfayonHH5GD
C8EcTYjzhNbIp/cRaLTP7+4Oo/xib1qJ+9coOU3zgfHbyaZdhUxEN3TOZkofwkyL
pCLGtEimg/4IdMD8ADOoYF47fvZXjRrJmXFkG7M07v9gS8Kj35MCczcBZ+KKvF37
uPMeEHWQb3fZnDRLDbgVdZgWKKHT4yA8scr06HitQG4Qs/1usrZpQZdP0UYFX9Ew
nEYpcmN5mBCRKjSSXUClKWMC8fsPB3/Ii5iFzNFDh8umGMG/dB0Z1AoznbIct/Xs
BstieXb9t/qQj1vdsWfhWAQSSVHMuZye/otAhW6469bugxtDRs6hvFRSag/otQ1R
IBM3GZUpPmvmkWCINqk3xdjtMTqcombFD0NwbNftPu1sy1H7F8ZP1rgeNojLDfMw
PSj9m1kliHFiqbyHkrpd1CvEvxEXdRqOPx5EKSTACw9BRKrxY/nGz6mjRKpmWK1h
C7Q42hCx+QAQVVTl0pi3VByK4BeSqfZw7TthFi97in8EC9OIKBVB8KOFJFaQ2bsG
t2JElXvp8s5Fvqc38KFFQfztHOQeD9yUnkX/hBz8fuzzv2trQOPfMBOxUoLQTmfX
kryL4+qxAv8pS1YzvO2JAvuX4jeGg54M9/0FZWRi87XWhssvwKabVm12cbmNuNSh
Wzr1IXSmHRm/A7SFVkrgK19v3xMh1oF+Q+trQJwF9G6bT76DmvXpoNGfqVaCrHo3
5ONYsTPutGPq5cdTBaZt+8sejq9Eb831snKcFjj0mZkmcYd93ByavurSkPLZFO83
QGzPAwHDKgQmPTVdAeJBaEeg8e+LiVdHYY+/vnyEOPeOgLXJWaVr7/7LwA2U5Srs
akIOiiCDqK3QnUUkQh4nffq936lTP+tzGnd+xcq7nNvMfRtP6ptaDK+8YnWs5lQg
dTobFn2Bgc2heyt6tzgSTZyxepu1vv+7xKQzC1CaExSc3qbPudggbUt3S6DNDC0X
YHaQckV1i7G3WcGFN4SehQdRXCr3QbegVic6ZdQVyYCpDTvnMEcQ0zwMtO0jPiDf
MnEf+ZkpMCZ9qw+em/y5730x6QFPGSFTGdrnrYFPvkR04XFMkcVqqDgEdK7iwGhm
7W9u4k185xKTXbdXaPSZ2Ukcm9X/WxkwQTv7ff6/uNC2UqCaYn4BmzRxu5n1MPqA
1rhAeBIDAYj8EHgtmOj1PnoVpS3rvfKHlRbGpUkVqJMLCNoyoO7CmYy0b852bfiY
kvcXuV7JfA1Ptpex/lr6KNZMzEsLiu+nH1VTG6n/iqTp3uIgZjIWmvFrEybofzNR
7wIS08bK46wNlH89bqWzIH25wOwHBaF00DjEVM2H/pPsh19JV5ecWPakRg0O2i6i
D5Cizq5ZG2bCv0/0SYuruAtMcIqftX+JL4wQuXYDJ4Hpz6QRxVKxA0wVA+MlEXWb
mXqVY4PcZCIqLoA9k+IpUtDzmEKN64sh0tle4+KcZBIYTDD4MW33WDswC6a0vI7K
ZcbYLGnn6GhoWc/tfPZ7dqeVPRqYDK6Us7evWJv9loyhnvpVGi7DtfuPNKB5P3aR
qLcGS5KXjYgihjV80V5+CDTxrMGKw1iangZ85PccOP1ea4MbFn41Wc+TsximHfO4
gh0fyoRTAw1ZKBdZMDERyAwrjRngtbiIfn8nI3VVDEgsttEtqjlT/+XFtd22aK7w
g7rnT242xCwVO9ohruV9vAPkmqRBUBmAbSzigv0FLmcs+y+ejQUc2hsQTfXbSGCD
WWU9xALEVHcmE7vT4Jus/W02vPq9nGovao1mqLKSaTX4yDYMh8786CGilZQNFiZy
WZbCsa3NlSgR9z5GrWg6oiINy1mjr/nxnSZStdUYz7EaknmrCO+8iJzQH0xo/BUk
RJbzvO8Mn1O2Wpbv48YZC/9g893gCs757RcOP/pS5RLpmgJCxvaDFsGINxAPgzHw
2tYVJWGEyh/XpOQE32ayaIlI69aRFw7+1o+LESgC9X31vW4FsuQBwR9zyCckjwwt
2FHIL9ArEfmKfja+ede25lct0ATpHdEWlJdCC1etGpaWxMkxtmhJdyQXtK9p0Jw3
9VTpuVCwGLPRI0fE7n2tiQ9VJNfnKk4keE52KNNX617XhL2hNZcjyPEUP9rkxgHQ
+1M1HYKaEny7pBLCQogCZxXzZ2FUp1FHoJ9GaSf0hiQEoVBCl6tookIOvlDE1zGE
DT1MtIOm9XszZEIlk0kd8b4iTJL/MBwDyF1hU7BC7CfFCdB5/Dqnw7PSTGPt0E74
mYYuB2nFeFGoYIHSS8PxoxJWd5tFjo7eyjUG/NjD/wuc6hAu/7797me4CNhnq2C8
oMrPd+G2FpIqx39g90FQ/TVc4Z4pbO9EGq2yk5Rcw7F+CDuoeaqzNg0qOCDhpdyu
6NxbRQB81NIWlOVIXEFDuS0p7PORBbkFAkvg91b5d6+SIGVfdlCOhlTqVKHRRKc6
7iCeZecZuemFOKPKCJvytJeKbdxGofZw66uFzaU8fEEdipbhma2EoO31S52SpCLn
1fibY5D6yBYrYcD8VmkOticbq/3ef4IeRuJYwuIze0S/l/7cW+GC3yJobiGUHEGJ
Xp6K2/pTy+w7v9pVhOkhpMz9xcvy5+OvOxhZuWi+mphvDuDpVKl5KTCY1NZqmXHV
pPAkEwitxsbAZxPDrVUBEpqYPzHdhCe/8gJmHtLkh9GFm3HjD+CldeeeXawsqm4A
NiUTkD1tNO31/o1P53jZxnPOT+8uJnAOvnfiuBzVvDtnwQAr2ib0v8mPFvpOCxZE
Q+6uNA0DWb5eLBeysHtUjF9hN1kfOELTx0up5nCZE48kuW6sKevvbPO0V9VJKoUV
`pragma protect end_protected
