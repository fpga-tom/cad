// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:22 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dvkRFB8KSfw6dGxk05NQXBXxFb9pfkjR6A+a+7Lyc/4oOluOOq9yO/ujk7RrjXLB
QLwlgMBgKa/xR1rSBK+bkWWzcS5FL5YRisDZvnf5juQeGH6RFileBEoLA99yTrCE
hzVNgUTOhpatHwYEHTM/ATyFQn71AkI39NAqIU/+zYI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15968)
/Jk2XxTi9kru7Iwt04/HqLn7Wti97OJdxDX3T3c7NEC3b8hCk5wIymcPKwn1oVHC
T3ZCsa5ByBpuUMSsX51baugG2ceZkj0hYagcqyIemGUNMZQslExLMUAFiR+K4QMb
DzaYlfzdrYzOmn3ndRGhxmxRfNX0CQn0ILQBfXYuR1Iarcf7+hlQBjDMRZWXbBt2
QCiPKnfSdrGLZFcufhynwjdmCFeKcrET/AEkkuUV1OH+C+qOxnHuQ7RHztNG2X6J
Y7Olo/GdzcOZNGdH0RsQH09UJASFBSL6hp35Yso7GRtGqxXUtGevBQtmoQYV2cOQ
Vl1o5bGAN3EbZFN+lyW9DRnfaTnnNxGd36w2PK1ROsnoZfOnuqKpXAM2Clx1+Qfk
9HgCw7a/mBAVuasSvuwLlTHf/Sd+F0FmRnYs+jJN/UGCZL+KETEoID2sHL/zy4dJ
dL+Gc9b75otwdX+mE7v5GyY8j6/4Z+KkxJZAooQarwiKurEAiaVDaRrxAD0jHA+P
ggplpShfihuxxqN4sMl+ABGh6KXvEaB6QA+mJM4+uceek27WFH2uEvdNg4JQ6B8d
lKfO8+6NFIAjG37IiOAHsrGa9f6REDWlwM9Fdi3BZ9+eUfrRf1gA17RnFfRJ3Tr5
xKroKjcIups6kBGIAE4DtG/F5zSu96/1gyhY4phNU2jYvhZaFiZ6lbbsVSbCUBib
GKvtxvJxEQwmfTkf1Sh88N6ntuGY2pSsDhDIIopwCNj5LvV1oRqlU41SeE0DgGtu
FEc4H3CLpQ+9sBkYDB71f3Jlz9Wnohq5oHF4TPLfbn+Nh4+ni6EN4ID0rgCKGGM1
Iyj0O1bDHMQJ+jno87sfpKOocPyOne7QUCx1LeIy3HqRWhPIdn0trZv4AFWohlV+
+I+9FTGtV/l1tXmN+aqD9gftP40Xx4XpSf49+F3TmIrc8VvpJT1RcLjMzzFOWFby
m0kfP+RoTMqTgV0C07dOLLo4YGsmCXAwbPb3yvFI12V3IoXonLIphXcJjzqionBj
T79DoDUuYlzr9GF63ENx6u4ELCSyIUh+ATIGmhtlgrRZRYrXur+fmKc/Z/QEDKyG
j2hbOBpA2MHUC3weeIIMi0AbNWVy2jPOO4dQcuOpLcNjJwQl+Apml66qL62RFhzQ
OGXiKMfy2X9gF7HLGi5OGTmQkewEP8lS9rwPucp1u3xRoEe2u23KZMlPzbLoo2u8
B/cw7v8ydGiWegy6t2kXwmGbuVVNZe4DESYn8MlEPKbr7Lsrd/Gju+4upiJHoGns
kEppGBy/eLmIOF0Hevo6rQoXgxN85pKc32L1xQ+nToLxRKBH7KJpBt51XZE451iY
qieHNiQqrXgGE9BpWjAjsjsWnEs5WKOp+rCvusRnWOgdQ7n3i3S5aQx/WFmcQtE4
72fxiOukJIA9vtgMQwd0OV8c6giXB+9gl3UcfxiCQwmKyB9AZnpWyYXJy2vFUbqG
a12qCWyjLZ7qhxmL59BfZa20SiUaRBho8oiS8GPJA5hfaAoSk6/eO78Fkvf05Zic
sfKbXAgLm2RtHEOKGcVlQlCP98OZGktHvqxrg/ISaSgVm4flMVz6/SzbpDpAhx3R
caWPXiyietFGHd0Vr/7YW2znnlxKTsd9g2jUt9PpVPkmFSR69NjrdgcplDZDrydH
NSV9ac0fnWLQK4GBsTQ8OBce5SZeADiyJA/ApKrtVSFK2IuDpjrYiDMgkHfCtW/x
vehFDHY/jLIIypuuyPL5F6GpEXAmXzWDkquyq1E2rjg9WVJRHQ1tGO9iQ0GNevVc
HdGP6moXniJ00FJm8ZhjUx5T7saQaPRsXhtXiis8IeyOqyqNqiS4bKW4mFrIi9fr
4e/VxSviDUZFfEcm1YXvYEIJll1yUt+DL4uGcE9px0NB7UNSwlpk7x3SL7v5ac3E
lXKR2kWq0qG1ihHIu5cqYlqwEM+jASSKw8UsGXJQq5/dBigtre7C2EV0Pp6BjfL7
N6qtCoGZBTZXGULMwVHHKw1JjXuUAlknh/M9GP/GhCkGKt9g/C4E+xlIg/3azs9I
rrlN5HWe4W4GvGORuSLbOhfXTcqk4a1Mw+F40Ew9SPNMGHRpLoOq4ojE9lxAzdnL
4EYilZHqtDjJEqwpJGd2rRJLEAFAxQbiFl7clymLEJr9aCy5fkOteg1K1F6bm1GP
cCA6Lepegnt4zZXDB9ihEEDs3G2ffbwwVIxyqHU/EgD2h+pqEYZlkqWm9mrKWRoc
mhZKCxyEsoOrlPSQkAQISeZDfkQrF0jY/mP2T22IYXPxkn8QYJ8RJrndAVHzh7uR
MHrD+rTuQ+zpacph3Wlhrgsya1Rv6IDg4yMEfMpDWCOyfI/3TDyukxqjBJ3b3xxR
hcst7TDM6EIcRNE6u3Ph4JlYe+abJSKgXUVJFxzxS9KodzqranWEL79i8rCWRNpR
Zhy5yRABXIhmyUXzYuMJwQ9FCu8HlEBEbHMEyp1foyfrg2qy5sxNMiYYuSI8lYtV
DRiCdIt8ju9s+V2wbn3cGKDxNiHpn46weM2vvv1dB4dPuyDG681vUwwnxdnbSRgi
eenwqzzSUmo+p0Pk0Yr+fN3CV0nf2VQiGBonrULtnfWCFg1lXTI2fkjiom+2ryw5
UXnlQfuubqkkr6Bi4uPy2nbEIKwSMFA0HCI0+IUJ04iPaWoJT7kRbPA1GPA/6D9Z
XQcTG4Qhqnc/iq29WQDPFB7lq0klmE5pLQMlHBnT6YxHuvgjIEOx0sqaLLWIqQSe
dXA2UAESmth6OjU4OON7Zsv/L04AoIqFCY5Hn7r8Jfd3JoI7V5anz002U8Rnl5rQ
M2UFhvapW4O1M/EP3Xiv4AUdtDHuUrhcPfdm0EXgpcXzqkVMJCBV4tO3yBp6J5O+
UTnNKSZBs8NSsgRYbyS9E5EhJXrbc3ZuNvoM2OWcdYyly+qfA1buyQ1fb8M9y7BG
MnO+YZWaIyrYE58kByxI/lgtsvVWwmmfvKh/EntPIFPodbmUW4HZIX7FW6J/iZ0b
D0WVZa9Gh8PuJ9RYPEu52Vj3FbYiKE+kkTGMs89e0wKaY0nJCb4209iUiINm3pJv
9aVWPE8yXLD9N+JufIc36LufwMZ5Vm/EBln2no8ojMmejpKUiwyuMqfRs/E4thV5
dD9q3/RZnk72BJaixQqpM/H7oalEUNAyTjIxfGuj7PATA3PCOfF8jXco3FkAUs/3
3N0B58NT/q/HC64hVji/FKtbm94qTG3wurqBe1aXSr21lJwrYxDYnZlZMZWQVxxF
y3Hcjl57fnWiDfTLlADm4wqgrxlHfadGBmKCthZI8C+3FMsADlDBLhVPeWjhuO36
u/OGJrkhNXgzr5R/jfOJU3gGvB6Cm1flspz4OpxNmMtCMZ4txoHtagH5edaQdhXA
qqsEapRn8sZQwkxnHMSujE9pvh+Bps2UKETrqXNLV8lSNH1l5+Hi1NJGhalp83qU
p3knhP091751w6wDV4lqTQtlNWSK7ui6+OzUpUxuMpPfLazaUFwZCzVlmMJF37+3
1DeNyXqKImJNzOU4daS5MALAeOQFKs/D8nttXk2eXy11B+x3SLwiW5H57/qcpoDs
tIw3MKY/sV5eYW/WrR56+/bEkm4vBd+IU0zExGgK5FdFTDnarUKCgp0d5iygSwYh
BCx60fZHrcS1pQIchDg8R4FMtFQDUOQR2THgDGur/uXMam0v4ifCOjcj6H/dQIbn
X2xjYTsYSuUladOzieVwwmJETT8Xptn/CxWzN7lSOTkJpBE8yYOBDgBVHBq+2seT
7OcsAreqyF7dMNZftg0CB8b9E9YqYSP/IqhMprg6R6grONdUhz0e+gYV6uCw9PoW
/J4fTHfXgY+MqjZ1SOuZAo8q9a9r3Q10J+L8e2OvVS5W4B0hp7XOkBdoXS+X9Uh1
AA+QXviZJE181A7QueoTJ3ZIYlD1+LKCe3QyzOCML+jj0xPZtc1OsRdGSvDYNRVn
UMUyV2z000AhV3O1on6GVnEbHjqY+R06qpZn2PizlEYk4/+h/ivs1IM52cJJKgG1
PWJdZUWVUwDQ8VgOWPj9Sj8Yc8+SmydhrpmDaGLCHUtoVl39kYr2Qzsn+1NqNFsX
RLyStv1HWqGR8wqn9wlHugK/VTCSNZ8Xs9nzJ/o+kxj+3O4f1aZ0AHOAPb0eoJ4m
/L2fzf8gLyJ1F/K2mmJMfbfeu7w/A1BUTXDn8poeqY7bwFs8bQ9BL4mb0JkF2Rj7
nJacdZHKx3uuqdQhLBbEYb5wJSUy3eGlvz2SG5oNZ60S9Hd+SbG6w2WIQV69oNI4
l3pXcrHdbBTY6gW2555J1Z60q8I2/2eV29qaEw2VGPTjmAwyK8tMa+abeyx8klB3
HGFbzc/ElGbS/0h8e0HrAiXY+D7K3XLVeURzLpwl41tkIKFovKD0jum3GgGpMTLm
KZRRtVIvzngBvRQeDGsZEZIUJKDbdWRIhTFvu/iM7lE+lUrxu0g0Yp6aczOIckcY
y+CZ1mr6PedpxoC9sis09ipK5O/pS4FinUTi0/Iv2MBVSVnHZ6VMVser/hoxCO4o
ipmjSiRAKOHFTtAKE7SLVdUSmIV3noWpjs2CU0euM6s0ydYlt9KHiX/WiOJGUo9k
lHK+X5s6EUpqldm3XQTsGPoa3Wq/mXmj4HhTFeg0+gk5v4Ct2rsuXIm5oc6ZYCJ1
sxGxdzDZ4aT7jLGzm4m812nQkM/ghD/CUD1WDc3urUb5Xji5DVGQAMsL95TCwlSa
x1xLjmgSe+xY8y5a7915yoByyyi+wKrSWD8Kbr5fRIuN9xVtK6p8T+wdah3TE04S
haCtb1iHihF6LpMyyBlPD8ZHhA2kuOzHbOZSrkgh2h2cJu3NLI0Y+Cc648cam3mE
yzF1jROUaOFGwBodItmf9g0YmOEaTIluzgv5y4BWsE7AJg4Zop1rU/+4AJmjlvpk
8DHGeVX/SdlGZVypmf2jJNFib1bmAF5G1SOGsozv0RSaol/dmwBNcHDAtZCVOIFM
WxKinpJUVVQvZUJC3pwBbHbrlibzn5NAObH+Jsh6rACjLhWLGjfGWf28ScZzHeby
TYKKYosdUUgp+yiYzBcJdNemWZOzl92T7CUY14dheRziqt5a4EzedeSWOOKdCAHS
MlZbJUfaPkyFEdqfNG29vgrL6myzr3ry4txWvzPDh9afZmerCO/kzNmF9MqLV2BW
H3uUINgwz/+75vytw5YV0wFiGfOqn8IJ/kNycDlEjbvs+/r1WdMV1XH+I2XOQ5xu
R3OYJfRq62WrZr+slBoBnmWx8fZJmd9KxREDVV+Pz4tDLSYW3RzKtZrbzSfYXjOw
6RPsAK7CQvBdNA1pFJ604e4omqZuuv/mI8t4OTW3dZpQOpWHXzkCJzulNq1p8IMM
y0TCaHInnbpI9TRIDfoyegsFDFTTdwTLZWakP5Y2iqUj8VHDBNYRWvPvmW5jNpEW
dfeKPtxZzSekCSTI6db6cVq8Eb2oEGvW7oZaL8yrKEuTkpbuACVe/1ueXY7Qd2Th
1GdAFXWOf9zqZDpsnuM9PnPUQHkWVclIk5TnUIn2mQ8q1tRtS78vEm3V4dfGunC+
/BM8k50i1mWcWTYAGg/dEs0I7EBdEWNInXbA2sAY6cMmebUszWkiR3Ut0/3d+JE/
mi/FhYaEyWG5POrGjAv+VfI2C/aY6I4XzJJOnm//lpXZYSskzX2w8zMpOCxUOPeg
ru/+xzS5CEEtWofLgL07ds5LtZLYPbXyjkfeC+0purXEYHKqgi3Ku/pzSzrStMGI
eDhZGc7SHk0W7T46XoVD8obamdLSpbeNtniGXY4xt6Cze4NYyo/B8/T38WZ6ej5M
cpLN1+dGCjYuz49mgtluH50G3QdzUz8CPQyRNBhI+5Sg4JC6JrE3jxhDfEQJX/0v
5p7KckB5pv6I+Z4NvtO+L9hXDkGmOiacUxstWWjeMQ/qag9IzB0eyAPNO/H3Hb/m
GxpPPOkp3EBoOiWC1qqEr///mFC8I0PYcoGKMMt+97RvCWBwzkbPQAyRbHtFve0N
DFNw0bZekwgwZbB3FRU2LQqT3OydvObPVSL/xwBTQCuS/xxOmXHqQ2zJNvkeBZwM
I4KwOLERuVMAFwFBWEBAbQ03MKelVHi08H3nhKd/+4gkXjeDYMTpfwuigGTnJcqz
C9OwySUEr9w/c0iSRiu2ru7lGuBr3ZzAqatGp+A2UZwozeD0yKqCj7S6QMnmX+sC
Dr9khpg1BmIbqIvLRYKpjwIW0Fkz8c8UUOgg+gmN2u+uKLPFN7Q25iqmw4rs6Lw0
vUZg/zydGk+42jZ9ZoSJEqsg4+Y52GLHjx4kLkX35aNmNyUr59Ax/e1PfCd6TY/V
ax4F6XQMIniGzJRFSD9NZSWXwgS6/ECvDNyXs4giJ8WegtBTG7+eMw2/Udig++3j
0+eQch/Uckbxsi8exfrZ1yRPnnpXV/ORjtNpIqGAZGAVLicWivLeENWXxQffa/JC
wsqHOUgY3JH74OWXMQr+fRCxV8vYD35nEF3Vp56i589v2GYByKa8lhhtWpTqWCFt
zKcYqWe9tP7NnIIEoqhnmuyZQqrae5m4/9pJs+nJwC1y5SEIzQ7HuCCFOpbBBgII
vKluwRFrhyRshlTpAEuJvFybX+XtqH2FkKfdzQCQsypLHPV+qDtxkeo2RL9HrG9V
1ZOvCbOR2jVqMWQ4wV9t53p4nxcdz8/U33KH64rJ+pxgqsQ1ErbwIhQDxLA1gKST
FYd+w/76KRSdO2rRkeCfBnBYlcDkV1X6W4QjcO03MhhGjz+VJED9dfBMxgv3SyIk
Sk6StUh4XihJLnHE2aNi/4TSy4D8eYLzobB0CG3Rzh/UC5dM3WqGr5PPq+fJeDN0
0STdoyy3aZLieUGVRAC8yYzWisMey14RuVvojNzsPZHX4FkRBbHAnqL/5uMOLxrt
gDH1F3h34esht9OnztkUE2SJKtrD+Da2TnXZWWXmiiXnijjA9AC3l76lH2KbG3+N
RkRvYIkJfaABXAD0ceLR2oS/tWWQ9jIPIpGwpDvTY3NEDOyJNOqc8jRYWG988XaJ
UDfFbkSycQT5mRgA6IP+gPiaw02qoeTMCHHPfyT19CuqFVQGUeT0C0kyRkCS0pAV
cOuBqb+mr318xWg5/oHcnNC6vYl3Ti4zLRgY9E0AegJahtPOG9lVop6AaYGk9ILm
K9jPO3uZrdYTSsAvUoJyyxiaieHlg8H6tyO8JtfFCkajmtcD66+RjZxv5Hzch0vZ
F+x8PkmeacISzhxd0c8n1wsy6F0kPMHEBR/7pIOdhJw4Eff8kLA114cttWwyQI6B
N1OOzCEzfRdTOb6xlU0I3J9jiJoiq/2uY8/41Im1HKbFYxEnAKUWpqrQ6M+QqCAe
FqH9zpaCxfTN21QsxVsvK7EDW7AisZKoz1AVKsWyxORzWZcld3EbBBHdTMPlsMBQ
5xroNZ0HvIOPkh49GT/WKUk/pIttoC8QZpf6nktH0ExjuCRqsEh0/fmcCIiw88bg
b5vR0Q9YSUhP0TB20Mm6Udq+FnagFej4NZflkb6SVNipRbc12CnIvQNoJuy0QZ/J
Rh+QD8HfYx8dLFjH69c0qNckrBBbzM1zD429g/OKv7Q32dc8gMFfJcCl4PuE7TAj
zKKA8opalX/+Vd634qQy85w9OPAKLD9Bx8Ie3MVku6Z7JPK1Sd6mmbIKsvE4QoZx
qWNKU4NknIVoOvZn0juzaGR9PUvNcooBzFO1IxRNE/ICJTARtXAHXyu5XhqX+i9X
hLGKYHia3dw7j4saf3HROrA5CmIikZHzylhAtGEBdLGcNfwuGbIxm2euWjzz2oVY
MNpWK4xro4a6ztzHsrIOgIyG+UQmpDucb/ASmgytF5M485iReYBlRoAgvJsoIKDs
r7r2eQi+Brnkx5tcZ3qjCjuUAb6mgPN3bGN2moe1jvjq5ymWdlpj5x592lWlzXxE
iz2yQfvlLC4BXrpxMJ/CnYvomPvW62Rk/yqiet/xwTq2ppUEGz1p/8r9s6LsPNzW
dqClBYhjQ9yaZ5uoFEEPxh39S8jn8eUMhV5CcEeWGX3nVSpjpJWgZXH7JsBJN3Ob
jlJBE01+tk2tn3aB/HsKnkmaND43L0WhqASnOIdpO9jae4t9qErEIKJVKAqAW8we
RDlL4U2wC9y+WXjg8iboYkBMvjYVVUgO1Bz0+EjiVmMk9zR8OG8SqJtCV5YxoFXK
wY6SGzrvhJ75n4Kh+68AWRp2Xrpu0rkKPaProwbqaKWqZPPzRqYyobVdArACBnz/
c4TW5Oy0bCniseUMU0CRSGj+BNfdd/qYyLAQ7kHXJquig7cFqM7RuDpmaygCvIcj
4Z9f30esrwekSbRG16KDl0rYe+DhHqBk3NJ9leFmSzT/1Fl4imw0kq8tz78xkRIW
lRooBP0St90jm2z6kdtelRazCiKOfuLCMN0mcq5tsNUGadCJAUig7EKeR8WHW116
yrn3JAtOkMeiMsgw7A/y7EFvmIOrZg2vJlpqRdJWAW9HVnIfeod7aBsuVJpggJ9/
O9C8LDgR8jN0GVQgPvUVSSdNYj6an7W/ucpM1Br5nbR97uUlWIRBM3AgwstHsSF2
FJBkIu/FmVcAH1B4tL4kANN1t0QzAVJtbyDYz1gxn7dGVwenx/xulxc1jCqhhpXT
k2CuF6GRVbUIYXchXSXZ6EBFosHWcDz7YMz6lqs2vnpV9LIC+iKEy3PYOTXZsehn
uNjY2saKusUvLPBoeUi4Jm0CZA6CXytop5/nMAgRu6k/LYSH6sfuQtA026Oc4nsK
+OouFY6iZY9hLUGVSDOQvaoR169DNb7wXJg8bxock8hw1rLQq/80CZGGf0fZwY8M
LGu761714rMuonegyLB3JBmwYu5qYJxEuw2qOH286AXSFYLGNBe0kEoaf9ztUA2J
Jn8JmSTWn1QTvG8AllBvvlYHZtEL2a5Yg6CB/ivdBvruGUigEpeOPjggAHqaNj8D
8PNSnZ1lW2qzTNQfdjc3OYsFoAtkAklRT7oXRfU2J9xEYeR+yBffxZa252cCh0CI
3XMalWtkHB/5ylxbGduRo5e25o2TsQeMHQMRQRszMOT+pqgQZLKFme7512efhPTe
mwJjD4dJmXjrQg6WsjlIIqVIFZQSfRF1uu15NZ63WO0BbrhSjVBdEuuoHkGplu0/
/x93HYd1DBxda4041VLiYizwu1N368Vl5oraeEacBUsrkxmLcQ5rF3wodPeN3NQD
g9wmFZAmMJlEjb8F6SDVYWVHvR5AD3Gpip8RkJjVUst76oSqAMW3yZ1x08zGvfv+
0InHL5g5xcKfnve8CjFvqLh31UaGhE2+LjGJcv1yHTDEP90wAzahVRquaiUnrRJW
uEBH4Nj0jSzldFoJerGSmv7hjIWra8JmNystu9YG6TST+1Dzzi6sLl0NNAdXsWkC
jnasU/RtZXTVvMZ8kqp+bUWgTrEX8Fw4WvI4dhYIA5Gj01UW52Ypv5OtXk9yPfrK
lMW7fkRVGcoHZTyCT8c8+0AiS/o0sOSR7hmUjIWImDglDqLw328zlAJBW0Mdm1II
g9tJwsPllywz0ScK3JQ1uN6wYxvjn2JV8GhsiQhiBHns7fICIw0MVHxkpztd/B9X
ETiPYb5yoR4lSpB2Jl+JFwojno2XYK9JM8aZ/+0vZeu5AUfgm+vdY2ICGFXiUp2R
lu4rQNC7NV0po9QZ8uJ3uGsWddKZlXPXsyEiKk4v3Ga691OWOIc9bnjmydtYd+YN
IyGjNG+H2YPVfafHeXMyVgf7JGOr8S2bazhCXJxO/9npcvU4JYCDBfjghq599Sc2
+v4mQWzA7oywTd5g8GbcIHHIVa6+F6hMnqcj3SYNheLT7nVt+kpA6DnK9kIDkxrS
0pWsI2/FJpr7rLDsuBMqNP/9dWxyebxsocDDpIVdDLDfca4WhaLUjFlLqm0/ara6
btXwj74JNTMpcJO+P5fn5g2CtArxMp87T/L1NkWnXRv0OBdKN/9MonZm8TNhCfIr
OQsC30XWUA9+6qBhSvwvDgIoUoadrpg/kgdrrTqdNaWKLmaxB7XoHF5ft04+5Pqf
xxNaH1YDyzlomDu38duDKdOXK1h/J70pPDs8fZa0hcoYmWSd/mb1KDkRInuzy16k
NYViWx5sw7dVDzPDhO8d6a7rBT2kxXz8A6pad4iBRZg3YzlMssP9CgKTMrTZznpU
WSN31LJwy8dlVV9ysBi8r/sAHLtS6VNTMe1NDNoYkp8hjzgkDBriCjem35D3zYyg
75oKRy64I/7cCpKa90DY1vtkZHaQzJ8uimlFDbIA0IBaZzc0d1vz2jv/SH3A2loN
RsqjEosy4pHFzSyibMSbHPSHvOrsOukKAz8OKtQtiQe7+oRQlNE2kh3wWHFjnzgQ
Hn31lpQolhxcxDLZLL077YUzoHMl8koMYKPGc8k6NjConq8zAWuGqXcEfth4siFg
JfGCZi1QD9PSRd7tABwX4NTAdoQ60oAD/OMUXs9yQ/bHNdLY6KSN5D9zDxPqKYj6
qy5DCsmlVlInzxwce6r5Kws4UX1YiXb81Tmm0v0fnGGkCCfPUWYX4bSyloWcAO+6
QEDZFZT9uZvTM8OlBUk4Z6CTIqzMeT7p1huZwwihz92qPqGZtSqnh5uO+uZQDgJY
AVn2GmdaBzcdTR998s7TuvQTrDorCaIkrK5Ebd1pTL6R72JgULkgtAdQMDLXYv7U
9erSHHWIzbLXdz4YEYzB9rOeeHM872ViFE+tNlUamz0VS3//mLSCxE0+COEJQg8b
TaOIvT283kIRoVUc4zHarp51M8ChTd+FejRsRkfAWBmxsSU20fid4C2vUy7TPdRg
QYk4aPSI87Lm5wwzWkTFeFiLNEehSkHhQMZ5yWj3IQ8O8sljmp880IV2cPUoE3tb
gaCdfw87EU2r+Ipibw4kNumjvOmu8J2NrPYYKybGIrmbRcctSoGOW0sYSrn+cH6N
SMj2F8C+PJVPSsZkYHDklsajelCaAy4H4UDzUWoget2UIrySQe3SCF2he4d8aiBa
wZdqWvUzWsltw9JP07acrV0+7WRl2HcrWSRPvU+O0q29UOfMgTj1HWDxpQaEBzdW
B20U8NHhq9DaNk5e8bVZuUAyIhTEwDvecRx05Cx292pwGG5JCz0kiH417F+SU7u/
aZeAM5pMV7e2AyDUKwqafBz3O7JkepEjmJ1TkBAHdf2KxeEuLH85hSeD6JK3DP7l
ysmheSQDWRlFqO3+H254B9N+lJPytY2kxJmmWQMSOtxw2HBIb3p3xflXoRuFo5ZE
158e8Gq9XK7Dyyx9X/SkWu/Y0Nb+4dT75QkmcFVLIMVgr9mjDlWSNvq2TAJnX9By
Q6VyIUk+zRzUit/CGwQU0Tsulb+Rs6NOEsp7q7LvyiXaJdUGQBGrO0VRoV4H87VL
GihiU9wQIoGZELRV6y/E0SIRpB6G1YCFReotqLYoPbmUASF8td3aesRmQJO47f+B
5XHKmfyD/oggIYBwyl+XlErUXOjmxH0LLaTUuZZ57FRydcE3pTeC/o3b4yENZ4+x
Pn6DT5GTywEtNZT3v23vLi6Lh32LRLRHaXs3nWuYSUNMqg/n6yYuYwBlXjHBv+d6
61ygrlN5rAqklSPMpswGWHr5J0Q2jHZiK4O8XzFOmXxnOt/6CvYiwZnQt7exURun
08Wq4oxTBWAkFCrZ76q5qI960WY1Mc0T9DfQUKnRQK28q+MmdeY5dwHaDgm3+YaX
ND4CKmA+h9Q1e+Q09TGln9oMXb5orOAQDJP0d1Lyp+nGrmBPneOdZnhgKyt2Sq99
Ay7n8vrJ97RZ3Jreea2jhPYCdy63gF0MCx+HiAFAwr2Xa0a2UT/np+hHamHKfsA7
4qjLlg39fV5R0stLMrVNahqtGQcwK2wW2VnVM9ay1zWWEU+1WMJl5fpn8lw6a1lx
E12xcb4OC5ZTPwbVm67xu0z/lMgBuDk/4Ky8Av/3aSxGzikWQsRlxUriCAoYbnwh
xMf7tM/6L+u6ms85QUmWAF/MXiIFavPRXvH7t7DRcM9c1asvjQw31mdVSNeIUfle
W4v3jFRFbCwe4CgAPBzfD9pYG+Hgbm2OATEGjeZJLiS25eTjuJPUwnaw/68gvOkl
5Jhk20bgNWvoGABL3JfVx5PR57WIrQU7uFYLnKrldRMDdmOBLd+0RxlP3y3TcGxB
cdQjd+QcJPRXOBHnaULTYg1Huc6qpDS3OUGEy08OUIAv158NKlSs863/VA6y8JJc
9LrFqSLWm+YGevchJpnkI07xjnmJz2rg+16INtOJ43xM1jGnWCWY0XJPqK4d9Zf1
L5E8Vl1BKEcx4jrqlnzevCwuxfq3WYNQ4NnyHhA0SiI3oDy6hI1o/NmSHVqKuBKc
mOmYkEMmLMRNzlAuz9E0HMmJI7thZJUc8t6rkSytOqkc6cfG6wodYaMXjuwPNJdB
4lf+LM8upcDPuV5eVhaBbR7en+ga7yNVF1bn+GneUi3c4eVsB4Mky+UJD7rVBjeu
10tIvHDUqwCySi3l9jKB4Yztbg4job8GlG6gxn/uKLY+NObNJpdTYJ9DELoZfEQg
fXu98pNI17zdqNWtkGA8niH3755HDYzNsV6KA1wJ1qvZqYnfOr1v49E1rBXK7+YL
Ns6e1R4804pZNRkeTlK8GymvVnk7g6I4NHYNErQg6i+3Z5wZhPRYxyfX1Ls9RhV9
dB2kgQo0mz3GcRcCdQzqoUgXbKApnBBNB2mm94/JJK3bPnw92QEyceiQY5TzM8RW
Tc5Z+95AT/02zZv/NYg/bXswtwdMsec6wM08nT5JTKgiHp+a+gYCZ95KhS7C33EM
xbY43muiNyhFVcuOFFmzqRmD7FeQa+wUxhhU/TpWwb59ykqUb45jcEabJP8MoZrF
vKwl+hFdGm5vzj6nBFaWDFN9nf6kjSmLGQqqH7BXvopI1bo8vsJFS5y+UNQlbuWB
cYG7wEZz3dVLMGG9hxAHPV87PXZjoCzOvk/KhMl4QaKEi1e2MiVveqKnqoZ9CprJ
HYUVKkxvGiaZ2hdfJeIpaI0YHfoQ1MloiN31HaJ2OykM4wGgEMaA4XXZk5bkvtdi
iNFCawBTt60WOR/3D9LMEfx9uLbHnd0cTUm3h8loJDZCX0BJbc1qRGSmRO7SY4ap
Rl5uN1j8f0V9boFavIXtTpp6K0pvh52DTuDlrVlYSJOluaG1gYbPth8Uo0E9ECjP
Tg2z4rCYkYuZyl1obBIw9EU90+RDd8BugI1K87vWDWDpt3INiV+/6vWUrceP8bfN
hZKlqDDCBtfKXIlZ+HdJi/rDeBlB4Gr10cUHTabANyQXcOKwkxVh1Ya8COvzS9/M
aUuJtxyyIr2cclvDZ5VmA2RHcLMcGUMtBAQtCdZRc6V9E5J6ZFGle1PVGDi4Ht4d
BDJLp2RgdLzrTmTPEE2cun9/V/l1Ms7XcEBUHHlKU5a/Bm/vw+4kdSqHjov7b4uy
sqcyZhmqVBiQ0Kg7Ac0u8vM8LN57Lh+EaxiJxgEufWoy72ycaG5TEFCHDYTncq9D
0YalmxwB8O3Sp9P61B+Ze7WkbIjw4Zs/HwT+XLSli2RhUvuIA31OA4rVYjxHhQZi
A/U+tN5pi75rZOFHleG5rEVf4ZfkerQ7haMouKtdektB8PwAy/Ku+aNJ4FTqlhHp
m0YQ9LmJz5R3kk77bm+S63yyoXC6ODwK9eUskv78XUDAL6gUjgVQ5diylz3O0E3S
rS0R82LHzg7MsGgjxbmLlz75bz6zjSlWhmOUsYrYN3IuzGvn09sF6H1ePKXCFQLb
XcxhlqFNPmdJyYLJvDXHPrJwANhk/TtKL75LUaPn9n00ixuNNIgkYKF34EDW978z
VhiBCGGbnBYjDbQmzo7OXmHBqyoTaZsHSoPlty4uMPmdIYEr1b2axAxmoSBnwPui
HVHLhITn22rS223aEcpVNDPQjdXK/w194q3oUP3gxvzLaMazL25JEElSxB/O712K
Zo6uMaURGueyruOMZywZ/7iisTZLp5iTPQiinus3W+mmJg2EpQ+nsvoNRLpcAQPb
rj4FDXKRQzNZmzKZiPxXMyu9ssw7hrzNmCm8ITBHe6Wrao8FMYUUa3KHy51GKrhG
Lv7Sr3c/ln6kO0tfM31202zwKiQeVbbpGPfLsGSk4P9qkzcFHXYzadx1jDe5JxHz
t2U3ITHwS+b+gYUs9GjqKbXWdtZp0aBGtwo+II/Es/DTbL1JJ1jJj0pQaa4iyRSh
eHwsbud5JF4IT1jw4qs+bhmcSmqNqc4elLTzj2+0s6OL3vgIWZOTAs93o3+owTTM
uAn/wEZOur7De8LUvhg4i99Cvg91ul9g7ClS6I1QBuZQWYW4MtyO/2cSGqFqF/Pc
ThJAqIbkxlTXGl63arpZVjTXJOC3WoQxB3jX5eHQYbH03LEuT3xBUANcQaQyOqG/
1yfqaXQfik1rW/8LUWQr/KjcLnyxPCLKm6XYzmbtgTUNlvi96paB8XTKApzJoa/W
X6v7oo8KyUCjGc1sU54RYfNL3oRYAZQqK0OGXbZVmxfiVgbnnFri58Kz86xa4cFo
RGQ1y7CQvwuBWybfLWNU8Qbb7buduTq+coUxwx1yPHydexErDeYUJQxEn4N04LP9
x2dKajFi3TMz70ChC1NZQjYOSO+9Z92KVIbA/lXEcc1AQL4n/HBBW/GjWhmjT5hU
XBRre8am1Vev1oQfgUez0+Otm2IhJKgpCb4sAudNMW0WIBmKv1iEpj63CqxmUWj3
qkgQ/n2IIweFPWyMOfe6IfD7S67b3Dxw+9eebsbwI42mdWRLHker9N+TE4u86whx
FGN68IjRU/2ct5F7XL4IDXDaCYB2VhGXIYTEiv3k1DP6XHzrXSVc+GZaqJh5f8Uq
0R9ZaP4UUGD8P1Y59+HKJ/jBh7picSmVL/X8IF1zvPGXC2nPMcrYa/VzvfYJFQR7
wNJRX4JZjYuENTJZKEHzcOUNUkRXXvphIxod/GbrswNlhrzFrOIlWfKx1D2hAuei
f1SJYtn23ZPUWtn/nYmOfIteg3IdJaFc27FzD1OjoATaSzGcMZnKgzmbIJ34gQT8
u4TK8hmuXpONZ1U9jVfnZKAMEnA8UtbKAJ4WPIwQOExbQ7Jyp6VdfkUNq2Cblh1K
auEqM1Y34wzlUYJblbtu+RWJSdg4VJePPGd+Jvpd8q5fJB4W9ACLti71KF17kucq
vlgRKwGb5jZocVnDYpggZh2/NFThRX4hVe6AhZmaFKTjposggFFkxvuL2A+z5Y1c
P93NP+yvij/FH2vAlc4RKOXNxQksSLlfKlDAQJypC4OVd7Bk7WPEQgcbeD9UVyq8
RW0czTiLVchJtnJ5IhSD3nezuN+CFGbPdWzJWrNrlYYnDAr8YwI7EvNfEcPva7y9
sIdEx2SGN9qp3XdKJyL/9CZLyzjI67FU9uJhFhqxPd86WragYg8CR+kxOdiJkCsD
1y70LOK0JIUOidLvpObz1O5LyqlK1Dz6ydPqkrsY6/fvQ2s2bSmRJz7M4CK6Omp1
8mMTk/i4om9gowPueOn12UmqgxkjE7sHeJrsa+Pc+oOnt2FMqC+gjJgGLWgr6UUC
4jS01GLwAM3KUmj0W108nEXOzSDh6QA+PvgHi1/M6w+tmFkmKNfiriKm1PiKMe3u
E4hB5x5k5ebCXzXEmngflGrt+AkfHXsu1Li2QSFbFt6/AsY36yZsvKeUcIQmWYrM
W9icrZ01w0faMV0INxUGxpi1PVMQypZiXXyCdDmXmKmtZZ97u/l4MTmrtWOMZ8X/
oetzBujlGWZh7jH4hztGP9m/dJUALeu8msGSo1ge8OiXOmEeVccjvMx/ChQe3/hr
o9lqWjeHdJMAUu4kvFGxGf1+U9LGfucyCS7v/cWklMRpAKC5yJQ++ZULZtFQGDus
7za7KnVUDvEOa3mVDPhyBu2igIwZ9Puvg+bNR5ZcCN8GtzLql32aq1Dy6NP5afoL
CvWOCR6NyV/Hd6nnzMoVvAePq/VcqWIMfKPs0zYYQV+dcwxI1Sokyyg2KpkahkKB
se8bdUAigBxr+fQRpRXlx+KTM5eAIHiZskhVQoeRU5iW0qUo4OAZUDx7CQ655Wmo
h7MdHpFay0bnZAKttuk1CoEeeAM0I8c2GkzQtYnp3yFQTJO1vQR/agWdoiupt3wT
NUUSNwC3DRydv1UlWs+yXH1vjMpBIea5URCeoDnkB1KJ4yz1Q+xJMvawCHJILMWp
xskvR2mq6ksB7plepWgsBbtcZQLsWHm8kPd5Y30NNAnrTa+wKQ088qluduLKKo/g
x+tjN9QPdday1wS2us6ArCRb944y6L7n75FNdDvhsFNVJlne8bHUYzJ6HNMYvi8j
W4NNc0/buup9kBa0PFvEx7umM+edyQKRTaeoCWvhAteb2LsBLqghi3EW6uZXYA9k
f2UeBGhvcUlbLdAv7TqPmsqCEETmD8atrvR7zzvVnTz3QdFzOc7YGlh9wDxEGESI
4K2r6coCJiiI7PD+FkkZ+faF3882OPKiY+Epl+kbGGpLEg4/sDUJxEBe26lgTfC5
5BYKl2Ee0bK8QgAy9hoC0LQCXCmzLZ5cj9TbuoHqaQBu/0ev+cOnmHQUmtYiJ+Tm
PRhekdyh4UIEy/I7Uazt46uVXrn9u8vb7jV+hGO5KX9xW2BZrMnO5kQByp/eAEC6
ZK5junHmHzWidG9V39HbbAfHFMJfXbZx9yVwQubyqTA8CxPk+nmBiDbw4mdQE2ZE
ALdbVy1CsIPGLGcmNHXsQJnlM2nqE71CNwPdmL1KWwyKq6zqfqaMq/bsq74BWIXB
7WyCXUVTci3poNOMxINBeszwCQJ7h/gF85AZ94AYNYX4RluOGbkGScImGiPzyWef
zA5zGkZnpCQj+BrHXxo79fiy6y1zkGxN7forSaxUMsrT5V6EF0JPk3d907QGGTi1
7VVMkrdN72m8YwAAzSoYKNHEVUuN/dShLW6CjQ5zMaPQ9kuMqNwYa44gEFFNoupr
hFu3RciENcsIq0LLOyiF/9nKWnahn755L88Si3SMiRaxv1zGG5BIAfJnBZJos5du
1xHv3gB8lQBiC233iI3atVze03aiMzK9EDFzER+b62eM9Kr2xXjAgH2MXfWtse5/
1fauymzDzatSOrKbc+2nQP2kn3F5ibSSwS/3FgAxm78UsuPgbIpDJteQVbVP/Sr9
aQgzZ2Zjq823oSEpXzYll7g+jrq22ex4gdHek2OJBLp02wUP54ptT+Wkd6yLof6u
2rspsSkRSHL5BcadAJWuKrtpDOr3YSOlpQc6CHTV5pykOqi8HN4l95NYUyArcUye
52f8EvvRHzAdZluInF9EfYdyNZcsJoZAff+YVqd4CnJdC7e6UEAmtRCO5HqZ1zii
e7oZ/4hKHYLc/M/LTE7fkySVOZ5TfX9sO91eiHtBwQ99EnUYyXn0zLN3vPFqpJfB
IlJ+ypVpe88SuDnhOH3We7Wd3fnncC8CazN5bExfNIeBh5K7EuWxeh0EFZ/rQ/v0
laOuxi23yldexHFIqPMLVtFnPvjjXw3QvJOdNw8tFhtT0TK9brWAtDgWKxSkoXZV
73yMJxJ8CLXcGJFid6emb6UYN2hwc0ZyoSKq7GaFJDnPVteSFIn8M6/D/fzOQSPP
zshTdawHJ2sbeSgzuPaxGvdvKmuRCJHNfOHWq6PS+M1LICU3FMsLl6f6pWyzeoCl
HXD4UU4eQva1mZIx5VOeca7tmao8Dt7fvwsw6vReStOrtcvT+6aZYZYy7HK92r+V
KpOw2nyWhdHVRCB+HMbe0r1sAYTm64vn50DfxwBFSbKk9aJtTCr9QY6TrKrfoNok
mY0JnWA8wXjNpStgKfOOJml0OnRK++05Opjihgl2wjBgfiKJB/pUEdRiMPRXs8Ae
MZZAyHV1j2VMmVRjlR1samOYQpuXcWrIdcIAaMnc0jW7QCVDmsxHfQvzmfUcbed9
yFpolgoIFT7r8kfzSIvk4rBhvOWdazks+zhLIycCQd732L4ocKGzLx0owGT2T3zF
d7UZ/AQkYYxUb6cRTNfg19N1BvSg0PJAWZocN0sYPJgQzDjceAKFMRGqN7B3RhCd
sjJw9zIrRGOWZhh7PMNjV3ovaMqNc7FSy0ar2KJa0zd5Y97fRMnFVHD9BjPY0QO9
Am/ttgh1ok1W12Reknp3EtRCVHXW2Ie36BeiGRxV+8X8RnImJAgsNEz57QzMvF2l
U0B638PbyK1G2jrGhrqpVvOv5EBHM8kxOUsJRIwdbvyZTREr1I5kdPCC4SdYR2fG
E72oWH+cPPDbwLTA3YZ2n9wrHh2wkNGCe1yN0JYIFfJ16mAL6UnezhLCVLJEB5lN
Kl6DTRxODoqXIshHHjs5+0EbA3fbyS6kmB3HhWaJHMj80wPVfJROA25XSAZY0T9g
D+J4F6RSAV2PelmIatmvnh6UqaAW+fBpCl9RKo/mHHtX00iYNwTRb7m/rxsrPlI4
xiDeODHS2zYc2jXptsmyA7IEvtROwxJneSuLCTilPTBLKrJva3YMKd94DqSI1JHS
/3lgDLVtlSfy/ulZ0+kK7QREfelNgF6fp/tjCMZwnYxri3WCaVph8+e1YvhMkmg7
R83aHAumcneJDxzPee+quCbnA3+ZIHLjlHvXWt09b7mrsyCHbPe344Y3gH4BKGPW
EcDa6++VoErq5U0o4EAvx9OUILu+RZcVyR4ESJKGMeleUkEk1t3SAoKtRcxSvZOr
yaw3/p0e+R/vRTLiVUvGyJdBhXANF3lnct33kjY4Ai9nngQ6R21TPQPWjkpUsYsz
ow09MOMLbUcLcPEQA+sRu/tgEsS5wDjuqCs0wDHSAeyDHymJByu9nbTK0OACvtQm
gtoZcjLWepOqV0JcWK7Cfcdjx1KW9XYzPfDQs3K4BoCA98Hix6zpDaCTZrwiYkSw
3dK+IWW3xEZbzjSfJQQ1fIQvyXF2SaFfo8VvgFLl7Dn8dCRYlkCSCfFZ6JiFopYd
J84NNKpHKPtzglT24qlDGjikV0Z2E7+MKDshEBBFOUc+bZKppFtw0yuC42DPmRky
e4jmeYZ75XLaAsOMCKu7vLYo0DoHH365bKaKLcKy3I7VEfhBoo7bzPkDk0F7XFCV
HUQTsMpxV5WGAWpHwUeFN7Kfz7b+SQFAydJEnz2JMWqJawXl7af6DoIuW43zPemk
xSvEMQ9alH/WxGXpkjyXXQyr4T4UZyd7voEVG2yoTPn2bWfyg0a4dz5XFS/G+ayB
W7s47OsjWCXZy/G7nTS8pi+v8RrhEDf6D6xclZVn/v4BCg1vWS8uucLXsCEz8goj
h5bbCtCxPlPByt7xS4/wRw0IhWRp/wc6dbV3hIJFX076Xoba82QvyqKg14rPTTCg
xvB4QPJ+wpU3/bjize2AvUq9fBtP0GvmC75EQJPV3ZLVLr8ru2i3cKDdBU7l3Bfj
bspixJ6aI8iUxRot0VLhy9/t14rJjVwcNkXR80x55HyH/L3wM26P2BkiVQqOzMW2
36GMhfm7IF2lBT5wpZ00Bxe1pu39czlawtYm8kimNJSxA3dWNjCojLKwBSL09fst
2TSWjuMBir5FVevOaF7UH1Mj258nclslSM+498eoCp/n2JIhaLqQ6/AJzBrAsCd2
8HIMUafPcZStxkRB2I62bFBk+UR+AMubGhWwyNg2VBZP1K9bwba1XqJMX6yYhNv2
SsalsBRAQN/oqnqeArAkscyJqKuMaIDQWEsgO5hzgLc6w6QgGQj2TwIJYpkRU0Rx
aeAPPIrSkIUSLkd8LzJhA+BBNz9ejQ2DHhPklZv4WdsLWdH4bW4cINF9HpuPpRm7
pF7ewa00iMBktqBdX3rbiwPEIvNIQxkboxp2QI3wzP+yLWUe+5naaZy8DuzYG6E/
5J/R5n6SoW8kLW6B+BE5/pbaw96LYaxX1mxCzAWa++fe0htIz4mOofy1q+KDrSwS
OEbEaLnFV4G+H0uTVwjLD5Qf0AYoliRBF/mTbnXEs+R5+FIG+8Vc5b7CgVrg16z/
yFDrPOzYDTvf3or8CcbMUKwAFMKtlncz8ZVGPzdplE4JKY2zLGZfgVdr9AsY0Fg0
7PXYYrsu+yDcSOJT/wpF8inHc3MWqLssdDayC6kVOfyIhxGUxyMn+GTJNTsCvnWg
sPkYbBT0zxyQCUHlAylS/UcKcNDyP/86ZIuTZ2SvqZ96jvCcQfHGwX6YB8epP75g
PkZ4Is6nZXXUSuxUVtXyaEeW1sULORCeskz5IamGmO0y5fja792oPAtxYJVlzEma
tBbCxIK45I4Kr+doUTi/i2oiZgBjTU0uBKMRNyqQ5BGX41JV+a+eOWHIFrs7G9pz
4oiu5JqzPgTQHwob4mlaFQ64AE29sSM9+5WufJtyhZ07w3dt8jU+Mp49B6lMnHZp
nd0BgwaiszrxOsHx49cp4ZjvrBSX9r9HftQqnM1SNhCxE4a4d2hqJcE9h+3M9dAz
cleL8ygtfdg+wcT1FYtEcdUYhOW1eGKK/HLL4Exrx2Fd8USRgEP9Ro3bb1bTDCD8
z6eyJwAMhvwepZeqNmZ2w04kunF+7awUOYgdZglPbxmsl4mYZX6hNolhPAu24avW
nsAcS3k64IMHOd/DSGlUi24c03agXiJ8twab2AYf3rOOqqi7apxipeO5Vxf3/eZn
ZfMuccciOeUv+HEBkAu/WWTiuOhsj6+zG/vJTlkl6TM3D04f9ED3VGM6OZxxu/u5
uTkjKZc5xi33GGYIliEq95ta38jXNcOME+4oUI+YPmG3PVi0OiGOCTQVgZdFSoP9
krU1sclwViABT02DcC/cCxsPc8k8JgFMU1z5f+OnA2s2Q7/HG6kG5qS/KNHn4U74
nwPNo64to/TUOsCGderlyIDoF7akNZy1BMeS0nZo6+QPVDa4bASrbtJZzO8iiqIQ
uTflZ54vzLANo0UWLMkQJL1z1OW7/XqKjaMlIWwvnaz6u+SQ/+SXD/u3D3KpOPNq
wlestjvQ8q6PxkDIo6BBYjNr10lGYj80wSQunybFTMuUJ2roHqD1RIkVRO22whWD
LpSslxFVoVwnDMjLeOvitFlaq8FMB0ljf2O6kzDlmX0fwUZK58uY7p0v+wHd2RAR
reLJdCKBeNrT0xsfKitMfZ37wvxm0h74VxxvOODeHkQZfr0TNun86mUFNbye4EYG
wVRaA2aTcmm+QUTQjj/iOWWHYW1UX6/jqRYrJM1+I6dMgvnSpzL6H+PrJMqzVTtX
oCWoI2/BX/n/icjb/XBFlk+3vmNgFnx5jw+J6hhQjDasXGhS0EuioNIQj8ynCdDf
hlnLcm+6yp8qks9dazZqaqCXEKdMrzORnSwlolAa1LU=
`pragma protect end_protected
