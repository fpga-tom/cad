-- megafunction wizard: %FIR II v15.1%
-- GENERATION: XML
-- dup_fir2.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity dup_fir2 is
	port (
		clk              : in  std_logic                     := '0';             --                     clk.clk
		reset_n          : in  std_logic                     := '0';             --                     rst.reset_n
		ast_sink_data    : in  std_logic_vector(20 downto 0) := (others => '0'); --   avalon_streaming_sink.data
		ast_sink_valid   : in  std_logic                     := '0';             --                        .valid
		ast_sink_error   : in  std_logic_vector(1 downto 0)  := (others => '0'); --                        .error
		ast_source_data  : out std_logic_vector(29 downto 0);                    -- avalon_streaming_source.data
		ast_source_valid : out std_logic;                                        --                        .valid
		ast_source_error : out std_logic_vector(1 downto 0)                      --                        .error
	);
end entity dup_fir2;

architecture rtl of dup_fir2 is
	component dup_fir2_0002 is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset_n          : in  std_logic                     := 'X';             -- reset_n
			ast_sink_data    : in  std_logic_vector(20 downto 0) := (others => 'X'); -- data
			ast_sink_valid   : in  std_logic                     := 'X';             -- valid
			ast_sink_error   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			ast_source_data  : out std_logic_vector(29 downto 0);                    -- data
			ast_source_valid : out std_logic;                                        -- valid
			ast_source_error : out std_logic_vector(1 downto 0)                      -- error
		);
	end component dup_fir2_0002;

begin

	dup_fir2_inst : component dup_fir2_0002
		port map (
			clk              => clk,              --                     clk.clk
			reset_n          => reset_n,          --                     rst.reset_n
			ast_sink_data    => ast_sink_data,    --   avalon_streaming_sink.data
			ast_sink_valid   => ast_sink_valid,   --                        .valid
			ast_sink_error   => ast_sink_error,   --                        .error
			ast_source_data  => ast_source_data,  -- avalon_streaming_source.data
			ast_source_valid => ast_source_valid, --                        .valid
			ast_source_error => ast_source_error  --                        .error
		);

end architecture rtl; -- of dup_fir2
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2016 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="15.1" >
-- Retrieval info: 	<generic name="filterType" value="interp" />
-- Retrieval info: 	<generic name="interpFactor" value="25" />
-- Retrieval info: 	<generic name="decimFactor" value="1" />
-- Retrieval info: 	<generic name="symmetryMode" value="nsym" />
-- Retrieval info: 	<generic name="L_bandsFilter" value="1" />
-- Retrieval info: 	<generic name="inputChannelNum" value="1" />
-- Retrieval info: 	<generic name="clockRate" value="125" />
-- Retrieval info: 	<generic name="clockSlack" value="0" />
-- Retrieval info: 	<generic name="inputRate" value=".25" />
-- Retrieval info: 	<generic name="coeffReload" value="false" />
-- Retrieval info: 	<generic name="baseAddress" value="0" />
-- Retrieval info: 	<generic name="readWriteMode" value="read_write" />
-- Retrieval info: 	<generic name="backPressure" value="false" />
-- Retrieval info: 	<generic name="deviceFamily" value="Cyclone V" />
-- Retrieval info: 	<generic name="speedGrade" value="medium" />
-- Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
-- Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
-- Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
-- Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
-- Retrieval info: 	<generic name="reconfigurable" value="false" />
-- Retrieval info: 	<generic name="num_modes" value="2" />
-- Retrieval info: 	<generic name="reconfigurable_list" value="0" />
-- Retrieval info: 	<generic name="MODE_STRING" value="None Set" />
-- Retrieval info: 	<generic name="channelModes" value="0,1,2,3" />
-- Retrieval info: 	<generic name="inputType" value="int" />
-- Retrieval info: 	<generic name="inputBitWidth" value="21" />
-- Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
-- Retrieval info: 	<generic name="coeffSetRealValue" value="0.011459181505378719,0.006662559453172948,0.008441885586611384,0.010405392494141283,0.012535742680276057,0.014799889271815258,0.01717004967250996,0.019606469859767797,0.022073648142220164,0.024514249717149376,0.026886111105804966,0.02914864878504396,0.031258423590992936,0.033150766468678636,0.03480833182241072,0.03617518372488565,0.037230261211738405,0.03794659522867296,0.038306233934559,0.038306233934559,0.03794659522867296,0.037230261211738405,0.03617518372488565,0.03480833182241072,0.033150766468678636,0.031258423590992936,0.02914864878504396,0.026886111105804966,0.024514249717149376,0.022073648142220164,0.019606469859767797,0.01717004967250996,0.014799889271815258,0.012535742680276057,0.010405392494141283,0.008441885586611384,0.006662559453172948,0.011459181505378719" />
-- Retrieval info: 	<generic name="coeffScaling" value="auto" />
-- Retrieval info: 	<generic name="coeffType" value="int" />
-- Retrieval info: 	<generic name="coeffBitWidth" value="8" />
-- Retrieval info: 	<generic name="coeffFracBitWidth" value="0" />
-- Retrieval info: 	<generic name="outType" value="int" />
-- Retrieval info: 	<generic name="outMSBRound" value="trunc" />
-- Retrieval info: 	<generic name="outMsbBitRem" value="0" />
-- Retrieval info: 	<generic name="outLSBRound" value="trunc" />
-- Retrieval info: 	<generic name="outLsbBitRem" value="0" />
-- Retrieval info: 	<generic name="bankCount" value="1" />
-- Retrieval info: 	<generic name="bankDisplay" value="0" />
-- Retrieval info: </instance>
-- IPFS_FILES : NONE
