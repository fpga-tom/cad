// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sBxI+6IjzmdqOmQQlwPwfd5hZTajXNscRSoNOiHl+gZe52GDgM1WI9Q4BtV+yYmz
0n/e+ZuL4hjTFe+eNwjSYdYyT1Mj6Ba9pOJil0xOI7dgcxNmuXb0UyxvKRZcDUDx
Je7KqZzjskSz3+ftKkmNJua/CamKt7tAj/0+/ZBtmZQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20480)
PRNPmhRPSEtVNS8rVeKDVT0EhVMbIAAwNMQwax3XEfZlBAwujWoSeWBaS7oFgawp
ZN4q+rnahSbH5ORAFWX/IAGKfXM8c2V6406kGsFUGZ/BFCJn4k1fMeKnE1m2KLfZ
nLu1pKbHBkYBtZqagk2wGQAjbqndMoc0TSnOEh4T81Ie335gfJXr3rjZir8vY1gS
Ogs+sFmHeFf8GOLXRSRvX2O2vqiIwDA7HQ9wRKz0ZxQSQfS7IahcxQbQ54/QO7VV
9C0J1ak8Tl6TslZyYy9mGps2Ce0ocfj8fpjWu4T68jN0AFcx669mJcQ5aGaPAQf1
p3ibxGV+LvQRpwWdzAFBNaJ+p/KcvMF7LW4rwDigjV78UgJcCgIig3gQSoNoozLF
UbaRHFXfDK8/+ZJcBNqGVtxfxjW/hydBQLWcsaVZRqdqqYoTeyuoj6AcLOOgnvDh
MgLLp3Sr5SyxjJx7NK7JNHPaT6vVnFqpyUWcUQvM15Wd/01RtRMvID06P21/Maod
sWf6rEM+7ViZU2W94zlvlBBUhXzVuQBtA4UkP7LpM0HdvmEcK9zNNTphohJGNBXc
KmtGBEwz86d74TMAlXbM6LJugobMY0O8TSwQTGWbfAlY+glmDqLPPId4/IEyGWdE
FtKwdm78XM5guYTD6gLh4r628NeAEFlqwbIVNICE8qqURADU/+/Wxzp6Jrl8l2M3
vFIPW7F5OmHgV2fkpbTEfRmrgWj3ALKVKHj8CM7dHEzsm+Eq8zJ4gDWD0d8JY+Ol
9n8kofXxHk2HTk0Ep9erhQTmoNw+Z7L8jgvHpBP0r3yeElBDP1aYQWhFZ/o0D84z
R3owvAnVoeiF8yEdUtg4FH0gFZZOTA/FMndAUr7hd7lPhSA/hV9O6yYrXv3YByTn
HivAc1teOgcVG2hvHkL3DBDObtvXT66VO2umMoRN8VVx9ICY2DWv+2H2qG+V8mPB
5EyTf8qN/f3PusWWxOBho/4PMubjM9XyjNqNxXcOWNkPiByjiLCotHZ3pYZsPdkp
uZeLHlGlYigZUr8p+G+0fNSw7wiDm+/zSnUk6Qw1zkSpnxgp6RqD6s/xbfDVdoV/
Grx9lu8SFhgGIJ70kxnd83V+3pulIkrhJwoyxLCBfdmIfaziW4WI86cX/uwagz7A
jklTz76kSZzYbpThxBHGYSQIUZ2LO2RsmhXhpF2VhuCAxP4jUpl2qZIV+TmefTst
URPY7UiTmzb5tbevZUPClYOD6hcx/My7cgyHyyUg5eKj2fWJtZynatP/6LOQm3E0
HUNS/HlWRWy41npPHU4Oc4x893hQ3Ax59N8sAm5CfsIqBl/8Cc9qkFh0Wj+AnmZK
2zMuq86uavCsObRHo/DZryN6oMbwdwPHmp0f1DIHEHhkeFgCQBgnqAvMjgSrI8Lv
Hre0gzEkcsnsx2b66oiad7ECaiL5PIXP6Fi8imSdo5sj1AByDOZ/CPLspdu7s1Nr
tLuQ5Z09/3TGCaK/5cHR5q8qCeReA4N7ZunAUX/uk/RStJszvSsoPWCMq3sSok4e
C4hpnIGDKVz1O2KEIQC1tvFNV0MHtlxeO0PD8Hbtf2QnnlIrjWV2hhw8+64nhMi0
ZdE4hPrhEvrRqCJuBLlDLhuX5AATJkPvd4v4zNoCXzgU5TStWi0S+pYPKcMzuOhI
rSZUm81hLET2s/1okt2NuvDiR0G3F3pCK0WBoit1mZ0jzhQQ0dKJmS2Hp2KqNP82
vEzBhCvGrQZioZ+d03mRM6p3VgKtefTnP9E0w/RCx1GuV4xqRAQCSBUgGBwDSsKW
ESSIjCdm/uc+Fvk3Z5d4JyUSuZbC/NpyPy/ZdPCiQmtw4no8cl7RnMaZzeoQDTX4
HQMkmoswcBq68AJG/HHTy3GmHywJh1LTePsAHpJ8LSJIq/TWyVdwY1dlsJGxsvdQ
2VKoZsBdFECO7IkLmReshN+i6mjQo+FzR6jtZb2BIItmSsVFLKdux89LV/ELHeRC
FRWJ0dznv/Fw2Mj5vdAH96UIY5p+vpp4kVzEAWcmgRzoMuQaYNBwOMZWgZVkrpZA
MCuTRbugiLj4dW3ygzwMgmhP8G9srbiLzMTwrKODlKpz+Kx6xGULjNLkNC1/jsgZ
jqJYmGOQ8NmCF/05UiRuX6c32droG/uI7aKvB6l8ZYRzBjiQLVUacklp3sdYUh1N
tYMBQPBRh8wdMWkOqZIMnsL0tk9CEn4H/m4kejKN4PUx4zt7SHr8Ri3W0rivJTmZ
/11rV8W8pP4MpQ1NhozRqtaOMzO2breqGXoAka/aq7z53H+DL3UsKBkauBbnpfV0
SnpQHUKoEAT+9DsDDEiV5Tu6HobgQTfePFlSo2vIm7mLKi3bGFGuXLSnGsJMnA4l
05CQzlf7X5xIuPDHILBT0Mu05rM9sLEH9WLbvz74ziRITkhte/KqwXdZCCu88vcy
VxvVa25DEeKjE+PBm0zwMqaRDA7r8EC7dQT1bVJY7eIdr/nveRGPpLpvqS1RwSyg
yXqvvqtGdydMqqm4VSfkGtcqiyY5tr1IVp4wUNVdrY11EcCcAyJoPG/FVTb595jC
tFt/LvsZ2tLAgeyGhfO/8bu6tpdDMBXOpTDXAqa22iZTrFYwTkzpn5TwnOqIrD1I
ckSxxu1W5ebcme1iYGxRk3IUznu9cQuIOzOJJBWwoQJHDl4qlywfj1PsLlcr+H+t
VffVrlicWkgDWasZSOd02bkEjsXQ0F/COPfrzTfaRLXQpb5+WbpvytXfvXc0Revq
85NXu8WtY3pdJkxNInJHKhIOLdqchRxVqFH+LfZdM6+ZMydy77amnryEc7n3TXXI
QIcdg6XVyhccSVacmRs35hZyYgYun1j/gP1TpYqVcNHdf5L1MjxU4fACFZgMkqDj
dXIkY2P7Zmr65afaRbm8a64tuOS1iFouvWX/odozAdG+wlVQwXVkDmSPo3/cWLeu
QhGmWuzqIshDOR50dVWShvddqUTSeTTQxNGhC9wuVEppR47kw2ZPSaOXevJXt4rC
gmUqEn0qTeioX4s/HGVyHBCpa7suj9jNRjS9+H20TaxVulXuDaniLFkrh6Toe6XD
h2XGS2pOX0mcSC6DSdEaRes4rMenrhg5OeD7eE6pT54Vs/MAe9DanOWIg9yK9Y8X
p/8WqBquKPLcFw0LQMbeh9xqi4ipv/Nh07TA7aoYW8GdcpPMuheQ6xYxKoAKOBT3
HaQpEDzjUCBlm3tSUI9ycQRYAw/UNu8oL8KpAzJnkslGwIGMGO93rpZnWD4FSC/W
3LGwcrhIIquVXjqCMBFCR44WeGfj3vsX+2jVuLie9BXu8dr7AEpAqwTRmInnMSgK
hrYf9vrzP+fmXK4nr3PQ6ErLu8UuhocJqDImLcQvcOV7FPySBfc4ySW5Wg+0A7pm
HM/ouP9zL6euLxX2UNcThiArEAqfdXepFh4Eke3zpwt58mmosfaabMK1qQH8zczL
o6Oa8dGY1fIDC7St156nru4lgzG9Aml/X4nCviCNp6wNhc5q4n0oj2U+AOVjKpsO
LbJFdfieh2f9sIRkUqG544Sd6eEmFrmv92Btn4XOiZ3mVDZzQ6Gk66UzF6uzra0D
AEFOw3x9/n/BWp9NWhg0E6Zo9H12mMwjCYIyxadbX2LAEqAFLGnlGdQbLOZUj8Ov
ihEhV5xKWDcmvHqNHjbhlTpRnflTrbl7oHQxixFxrwNPl7TbexEo7RONH5pWCkeZ
fiBzPapqCte4RDQRR1RWCsxSNgAIpLf629F6XPcz8uidtYwqy1W1PVcslfLFOyjf
0roEd1cdJdhq+p0lp75QsFiznahhdxQT5Oy07Ip5AGZrwxFol2bbfDAE7v8kI2c1
mL9FqPOakTfSE37TXzBv5KMy7MZn01fiwA/G5LHPsucSDmMHee2qUTsXfnl9DwNN
2GJHEDB3Hez7BKA3eAl/FtOMuY297PPH30fuUYxL5WB1DIx2SF/YknfIV05Wi1tl
Hpc3i9o7zCWyTbM5y7UnyG3WpV6Wlq9MkgJntQTXO0LEQe37GleePIBT4LexOkCM
0RnnK51qOJvyDgYNrfnJH59VCBCbnFzD5hpD8OESb5mUIKBHPYFuoHtqJV78g5vV
VjOSIlAWN1+08fkBDq5Dddm9BfvQAHE6hFDTLGHe7VNDVZgt42kQBXx0hxdUBsNN
rgiiHUcBti3p1mCeGGXTN66Rvf4bcQPeoIEs1tdkdxZvujf26/w71fKYBmlFsdK8
iX9eI9EzF2HFhrmERYdi4O/+icTbcu55PG/R+77E7RZ5dvHb5kHNBV+W2exQKL5I
19rQr89JHSvAMt23hoV0PErz20IlkbaQl8oiiUtmFJ/xk707Y0fs86/lXkAbDeVA
dvFREqAl6D27BKP8qs/mFTJvwEv6BCRYSYSQGzvyNQRsdpzW2aexT1bFtXTFnKMB
InZ+uqWjE0U7ANCFisUUsFQFZC19+V2rde8KOM7Az5wRBtKrot+lxWDgxIi5NDwR
bPbJOV9zJFwCFoYvUCezSfY25bpJcSf2/o1/dVuS142YPfkpUcob9198N2UFMV6X
BBxMfgiLDzBZyh5oIbjuyCYH5aCRIOdTRyHsRxg/i/0ytm8JE0jF/vqp6/4rIhVH
tKD4wCaz8PlAejNqg44/BSaDeZBEyCtcbNZGit0OypQ7BTAudbDv2nv/lLQTtaYx
g2ycIA8+geZxprWz3MRPWo052csbxPyun/1hm91HJop6+vyqkZ/o9C9K53ZPXcyZ
XCP4x8RAGAIngHaE71AKW5hQOG+rkgN95oRHNjqEuwRlWhMVo+CdPfO5au6PfMKd
+ZXPGxAWA5U/GWV89vBO713TKaWJW865A7STS8BDgEMftkCRdFgWWqGWe4M6PMqi
Eqp/QSqSTyFDTMSM7x8vp5LgwvudniatiOefFcEB14/wFUPJsXdSHlY9rUYB6q/j
J8yjsvro+vHQeMuVLW45fiYMXF1GUYHq3jlEw5fSDSspgGMJBaWbFjm9wQT2MbTs
r+KX6A7nN5L2q6g3Vy8dXndgrAEuBu3l3SOlYr0Bn7lrqvZfGLirFKlMZJR8yBJR
Fr/AOLe5xCjAx8mmIetIErJ/a/9RGGXlmfan4CvSW7asT/ZlV6HJkqylm8eQ0aAO
XMWmOzHFFWiVYwvc4o2+rXjPR76ukMsMv/2wuZMiagSyPeay3HiEGlV0F3N4Hyu5
m/iB7DRVea2PfPZ3T/sTqSM1l5TmUPGaYcIQ7mTilRJjRz32euEvoa+hZ3xAX2Az
QfT1XqG06jIrpFeX2zL6CBhKnyXYjvNPX2h5JVyUZcN5i42qyW1zcNkhHiwU6KC2
2sMJpC1kAnxRAL4WqQvZM1VfKJK2ZWtgsANbgGy1ivYHV1JbEgQTe/Gc0nbx9Iy6
TuvYx2HDtA3bfeJt/aqTHC3Z+AEnjwUnLKgxo4E0t06bPolNQBq3c3I6vOIIxOJc
zs/e/zop7KFk7bRJz13/Skrq534J+AAPMaV6FKNwFutDdukib6om7WzM6hrziVSV
iMHzbbly9DC9BiHOOv07bR84MKxOriO5h8qttekXDIDQYEWiN2alzh8iNEBd/ITC
2UkTT5A72BM/IEIyIptsaiaBe3WnXQ1217Qfl4SHPnCi3I/1q6ejflAn2twTgzdu
VmzLCiHiAhJjjF2rLjwR2kSJECYbFDIFbcxTItgxd3mK6V6dIYtHqeQ5AYXHsApC
ryfFDCc3o+cjqKOvxl/vzgwhl8CjV4ttTM80P5LU18VTl7BPesRJGkKPz3ArFGSF
u/u+oOvMMDXVAqlXnMVv3ntlQIj5t1gvroZClHKFi2ilDnxkcbw9yg02iy0xqKsV
46oFmwlJaC0MWphJWMK1e6hUICnjLoDoxQR00/5bm0U4ydOzw1G7WzqJhPlZb42Y
/GrvG3ZXJNPOV4UQXchSuraifDhXD0gBtiUIUBqqiPzzEyjiNETAz1/en4uaYTCI
G5Qfacqq3OUQrbwXLl3veQJeZ8/mEsHIiu0qNgEnhhmU2YdFiVUDjbVdGbQ4NcXz
k7eslOdmHFqGQSpUMcN29mZvfgZtvMwte8QO7uIuigWzr5PZKv0C1/8E7k/yIDrH
SmdP74BRHAVZt/azPyGnhqQ2fZrsGKqF/iDYr+3FNeCNwkau0huvugCTaoXGVzC8
E5FApSUPf08muudn/crm8ufFsjUwSC8QdL1Z8fCcAFY7QQcrhltM3ObRL516z8U7
JTf+sLg+txG8O6QSWxMnTwMQqrfZ6A0JV5LiPgDRjnv+a9zrNQ5jLFPsgoKNZ5qy
sOrD/RuGOcfC3bzoV79wyJN7NTrDzcuyEx59t1W6QbIwoIz3M8D7BizCAIvflyYK
HaJ56QsDQ+o0Hb+6yj+yL51Galvh6mfXtqKS2iyjeMqHTqOhAYsvtijbKJ/N46cS
ug5T/VbVr7Mrt4AAXZn8TS53XWsspdIOa1BEtSibeknoZobwMbrfWbV2GKWVPdVf
yagrg5AQIRwgdF++b5bwKg5vevlfrUGVT1XM+OI35oPXL6dUwITQUGd3EgbpXS/Y
jQ/f6n9gRwRe8F7Jra2ByX2q2NDsuw5YOQq/jVyALdn90HTB98KpMxzwRuEPgCcS
em5fikK2/w7tV4KVJlJnm4y+UIuaBGSC8dyjXLTpbJSy3+faII5iEpz+PpxDE8Cp
YDmrM1140PmQsapwbLJJjzecRd6hlJSASEXAQv5JpSedQON703qINeEnB40yEPPQ
15TSFFnopCPniwWJG5uTDYPzLF796ye5DS+oghbJIUOghLDr/ag2HRzpqz42Akzp
NjOqva2yfl3GrfT+utSK5VxrukF9oWaa0nbeYLxocxlk1MzeIve6Jwcx/jMoY7R1
E/cX8fVY85Qkt0vryVUIVhN2ianjxmU0W1PF5VQs18ODQx+ZyM1k6aMmsidFQ0I0
8YE3IDXWBmz4p1KTXzYRNPAamB9FzlTxRByIa4mzOFvQYTdGk7e1Irj+YUL2hJN3
ZX5zkyU2EWS75fh7wBl7VO7pZcXzN+TfSSK67QspW0ILkzbSNgBHr+0C4bLhcpRh
cbt3D7vHqYdOuOrDWV2lPQcNo0rjTRz/aLzsWx8Bu/Lxav2e5gqSx3zzFmq89vum
9TrifypjmXYIJ4FQev1t30Idl8PsvC+ADKpCEPoOe+zUl5dvELIoOjSDhMVE4AM+
0TLjFD2X7GOQdzcSsy2Kh8prlS9V5UKB3vZyjsAd4SFVFxVz36YaOL71/sgRRBlM
tZ5z0X8mz8DP4TykMhcVgkSJWo2MONvOh8G/l5VouEEfzpf6/u7+ExCmka7/yoNT
yH8L8+TmPPVM0btCux0oFkZ/+CC23eZRIfX6iC4Ir0jv80Y0VDkDdo0eFxRZbmKt
d6eLknFaCoyioVNxNEELgK7Xn8NpkzVirNxP6dBqiTIouDK8U0ohra98h4NsWF5X
1olwFg+I0V9Zo8YgqzImRZwQ94QbaI8o5AF3rzppszKM9grK7RVJpA/lppzVZV9R
BV+Ic3SJ6KVN1ymCMW4/oARzgL9a2c9EDxMCsqFPdS8iKdHCF/rhT5c9UhN8DTRu
TpuMDAbQt54QOFgUToJg3p/ifKmLy3Q+vMtKaLkBHL+7Pvflx02Ct3+1IJ2C0a+S
WCmdfCkGbXFiFBAXFOpqmml86VQgSWp81OD2pj2g/brb39Vvkc76qMB3HfILSwx/
kxzH0geu4GjhQj0T1sWSxtAejY19Gpg8zcAGI3pOuBhmFmndZwiVFe3mhapb5m8j
SEifELunZaAs/WyziW82qpJs05xNSXUoYpI/5qDzz2UO478FpAT6MMMbhT7c2ZrV
6MrNpKSvuw8D4xZKSvTujnhP70S0mcYHNpMCifiDWORDxdWyoaJttESaXX0YT+35
dvDBmR1Ht/7C+U5qRrNIDSfMUgLxhpQqdJ4h89tpUbq9EKEMrt4s7OsWqfkkp9p5
oXZrrfttkhWdqoy3/WDNkc4io5mqj7KhU/l6Cafv/DR1JOe7cZZkpygrP9bntkXg
p92JvMzyV3LaWFEbm8vS0Cg9NduOSdIOBECagYCZVrq8CRjzzMStL+tCWWvumtmo
RHVL6Jq44+hSlsMT2vyj7jjIanVjSwqwXa7iTduihYPDEtqrqRzb8S0hUBx0IqiH
eYRfc/TDtdDmpoil7NSvBetYtVb0dvtXTuvxPj+RSeIiLh5uZw/+3GGln1nUB4/X
aTdzt6L2YFrf+tDi1SD3KZ/4xbKPG6seEB4Wr/baPTl8Q9B4Gzm+oTw++L299dbE
SCjE1XY52z2hXomtoIm3ypxm/YycU/jTof50fQ7Lp6GwhiOmjGk1pM9ThEfV+eNH
I++jjcemlRaf1dO4TsBVcVenxz9BvSpqe5Qp7oRTXOaeiH0HHMKHMR5o7GG9THAQ
9J0nMDuBnYJCwaJtyX7yYtlPiiuY1TZflbzJH9jGuJ15EgfVyvajluYuRVwZEGqg
2iZza9Y3FUJwnCxt+nI9blwjuE+StJJZl0Jmn1yb4UWf6I+5aehCs4y0OgZkUYn6
ao9SRNdt8uc5ctolBdgZPm52KWVWpyWKwNItT0gaTzH+kCwGePJQVtJBekm2sCna
BsXAd2YTY/peQ5nQylF/AEObX0Owfmh/GWMVPnis57gs4HGI+hoiklj4kGn1eK66
g2tvBpDzhcvXouNW9igBMaMFGrMqGs/mIG2SKTKWhJSb51a9S6c7QdApoT7Z/aWF
+Ejz8IuSiVgs1cdxEgExmK+uybzEROucyNWk+YowZund/R4ZG3JhRQj/HQLPUHHw
WAX/hyNCDIvcpQBnrEAWIFAEBbhvsFGfME70GLqXu4HmWIq+3NQghYa5PlbNbWGK
FNBwei2XMjPf+m2hWOcdZeH4Gh1I1oN8bDALDf4ju/F/iLNXZCLbzPY1x7AGkb2e
7IalGmVrjHFiG0JMXf022msDCYEqcWbSogkzsaF/K06ew+/oL3SDdALYtwrNGB1i
aotB1IAlXzPJXu2GgVTtjCuRfJDxAGxKfQi6WJCCuMoS5UJk23CSmcKteQ0EDm0J
M+yUskalNuk+aDOIeIlhEN80fKAjKmmVBQnyhOr76Xj4CUehqWcH4fPhrvXeMIk6
l8dGbv3JdTUqlaY0L6OjLCYQb5s1S8lPNogW1AbNxe6nVC9LT+cJyYeOhFYCbxZY
JrlIf3HufZ3WAdefRO/gxNunMZp1eQv6cr7eVh3oxsvpL548Ogi6nEIqmHfRPM4I
SBA4okRxV9TZtrvJ8jDVXcHF6naJ9MlAUqRedqQPfMWzUl6SEzrpOITe4e7Pu1Oj
F7L2Lnb7qSNsezqC9wbcxDQO00prpaTShYc+ridz82fkezgPU8uodXM+KW9KVuVP
2bGGO2lTSWXmcdASv3oORyjw4dBvLM/wqymi4uzh2EFEMRb8/TDrS5DJEZQzsSKk
E/sAgCbzc++dnhoynmJtD1FiwrALqfXTOicGcXcSVWmTC+BKdMHUKqASDqOCxUOU
3wPPIJ8fb3pZoxGHveF5i2sD7O4AO+kc4RMyyjYtEOpmyROqQ1t++Y+28jvmCggA
xziJnKcoOGjdg/k0ID5PwQtj8utnlshyyRiRmdECwTh/XodjmUT191m92V5sugLm
Q96DGjFFg7vKdAIeya9RkIuNGdWT5k3Ax/qxTnHUcnRPktnn/GvcqtapRlT6q9q/
wyUj8/NiydXblrdd6TgmMJ0MFQnF++tukXFecvdA1VRzL9q3WoXtbyiPMMAPcBw/
yIjsRG/Dv4llPZB9bOyyjS+jouOEtiI+ZTJO5FEAnOfDVnUnOGW573EkHr4jf7Pj
AKsGUCf8vVRqnQlaDYhb/IPA/n7bGfCbpWAHHe5euKtKXGOKi1Q/lcn1IWWRBKtE
DIIPb+PLXV7zfsFWXdTK+TfVg9YIydADNkrx9TM+hg+3ZJrzm0C8+7+u0027QMpx
x58T/NYJ6zkFH5E6hl07uAOaNz97KslHyRsDV/fwuTf5C1B9ZpAwtJc30kXKsVe7
XQxKy404aR0QsvayhRYagtVGIpfPJ/q2vYsGEbirWO1bj4Kao0L8S5Vu2RiDoIOW
/jqU78Lpk4b6S27rWsFRm4ELjP2mIL4n37cckpGW8XfDLrL+iVQyj15cluam/dWX
XFIXtc5bQWa/WOQrqmBoHIEDQic9gOPd16gttKhK8yJjtfMX+QJP2BfDkOeRXOPv
Gk9ygT4gmVLd4xQJGdTxSy0v+kXpg1ZgKM/JIYPEPhGJBYOJx9K9/YeLEcdvJjL+
UiBrvqm3Yq0fPXp426liYIDdj39ZpdWtxnlW37ecw6IHH1gGxBy13r8ygTYsw0hW
I3UwqU/Dn/UiZysWKzMC+lTx//e9bmaRp+hZGVnozTw5uD02WZfaGhe20vNhalmO
Sbz0EeC2nXJZNVeN/zXtj+l2LFFmMc04ZrHJrZMQcFvmmohp/C0WyAvdXqH9Ka6O
SEjrIUdutXaqrlD51P4OynKm0pRM5hopxBy2yZ4Sg2LY/h9sDARp7dDiOoE5m7OV
5TgG7JkaC8Js8fvj2zTnVJNRP9cj3Sw3PgMLFYtd6o3abLoi1T/XsruoJLGZi+HX
dyh5oNnBJrdy60iRiQWboMfmWT6a071h7aCNl0tZtZRMc6fyqLgvxeUBOuPYS780
PEX+uyZpstGDHSxLlcmibq+HFazq7HpUUF4kE5pQEjNtSxvCB5TnWwDft2E1hfb2
9+mzs5xzcB3tEpVREKUjZfUAqfKDN0pYRWSnVOoGxrkav1C92tVSIFrUg5CxFT/Y
WemyvIZG/FifM7VF5UEHxUUugLh59HUrJ40PmVHWhUZawpMn+GHCRVuVnNPnUXQq
qp8yoOC1ENmT8FtjyMwZ5By9w36EVFUYBuvogMQ97anhiOrSDry3fC0WsaLMn0tW
QThvqwxC/j856Mjdovh4ER0isfMzuv+hzWzDJyLTK2/bITwOnfWRdw0F93ZB9jtT
0aefnmj+MFj7aNvAQnXvycCAKN48YlrWlyxs+HwdCzFhoz9X77LRy63h9fo1rL2I
3Dxslz6cMC3tkCwNns1rUvLewq42OrWM2LZI/x+fzWuhlQZ8rGTG0J75zDPgTxDs
zoZ5oBZTFgy/ilIy5s3S3A5uTTBwg+huBzCOaz2y9hem6B+rIZKviRWlaBgPUE3+
jZc3O1yPGlaXsqE+GOBGtZoQ0lY21jUz6ua4ivfOPCWKfaM+/hf1kKLI/uiJEEhY
aiHxIzQZ0Ij/TZ/5FcFq6Lw4/1lk7ip/YnIZChl6N2qIYKRbXtW15fZHuh91Z7z4
MGrc022VDmbB+EgmIel9QPHYFN/YX3bdBreE2i8lErHTB1ZqoZf3F8/N7sg4+Wen
lAkAh/9vQRIdw2dr0LQrjRWVSiIID7x/Xj+d1h6Sl2FH6CwFsrCGR4IipF0Ydp/N
j4Oec5AdgW3L2ydOMaOhfeoenPV0/LmcDBHa8EaOKnC9NHxfw6sY+IAZt5gZpahT
j9i9YK0vswyUZOdppEkIvPnHSIcDi1iOyfreRWoulfe/huksIKzg5jYqJNZIuMDe
qZfGhVWWZoB2ZC6w8xLmHqeUg/4t03fHA+JLrYJcoI6ojh6xfkVlhPUVcmjvuZXG
DPKM6J1bt33McMQfKB8Ie073LgbKdhv0yMkf3cJO1ucNvHNhDzn0HttuLQHPbvzx
Sb8hBdnAvNcqGvMhYdp8k99e0wkq2LSdo5r5UPZ43rK8W/rATBJYvvLtCq+PoTWe
lT5R29xA8gKylr5MIriClIDdCOsOLX1md0MUrebQDFdH64LdHUeJFFUzffp4yZ6k
MNXIdFuV9/MDwRvxb2NBFbJ/ruNTfIxQtZqYxtdCm3pTAbxXrzR5zkacIDBnt22I
YSTbkp2MCHRL1upjc78omVbws7W+UJLeaGEERjI69dHCEDVKSG5HTH488lXrBgE6
qoZ8urBUXuiokemP3ygZdwt663b6MXgNASNr8WV6TPWUGaeilgyGsVKlS6vV7Nst
GmRLi5dbD7dKgK9b8BaJ0gLexKV6YqgXzU2rJd/jT3Bo+8Y8rahgHh0Qivtkx6gb
tSYonTpPYKss2XFVLob9UO7rBM2AOdwQzuQQqYRfLoFJmZRePj4ZktBq1/5O7xht
6EeL6/9PDi2iYiyKkRPSlJRKfNRtzNg6YSySEfXaVf+ynlQaWp2+RLh9+dd4n/+t
hODf/+Az+AJL8ipTrt1SnMdHEdnaD1A0nwPomcy7P2NIMy8Yf79UTgBhKiJ6ActQ
wjQeLCpF9YuO+pZWBnxFLcuE1xDYX7ERSkvkoyydS2sHL/5CwaHEaFDcK+4tZcAn
zdSCztP0GEnTcF3pH4JliOhdnBq/E5aE/pzlURpO+WK20U+CGOX2YONBEroP8Utd
EYPGu7MGkLqOc86jChK79lZRklwz6ZVJPoz/i7IfFt2yPB6LifCzgocP2EN3Yn17
8t3yNTx+fzEBoftZjAJz/bm4mgWeXy5qE0K2gLy6svtj0UDFRDXu2kgRIYPqxsQz
9uXsiziTQLrdtSdxn3I3iVlqLwxvp9iU/ULyGUSbTrgvqtJymbSgiqTv1SC+5juU
mTJiVcHPac2oBMQ+eRWBt0u+pv50l9uDOsNjT9JEwTF1kAqjDYa8eh7la2SeiyXh
uAUi+u6SkTmqO53lYivshPGkZ2pwLZZU7/kOv3SR7mzoEdQ4mZqE/UaFpYRlsRxa
n54KP9o4xbY6NEdwcO7rGrmlX1zjCVoBMNWFEWOwJGIvy39bv756GnC9kva/13MH
Mm6bYrj4+j55MSVOGRmvcn0rtkF0e+vgxzLFAojBXYGWZqjidWBj8nBqzUBEkICr
pywMUnlZIYQTdGOuoB70taIGGrF8zHhp+fSGVp4OTtX0kSf0QXvC+hlqBAC3V/3B
cRV24yDljR3EOyycPcpth/w6bbolqHohICTLScpyeghSqffSB0m+ExDpptTKJ4A5
FsRrj6OiM1uD4+qw/CF1542izaX+kknJB9REkhdrPWUzsMH0tiHSUI3Jp/3yVgKE
OwqO9LQYbWlOK8ZQmrCMPvUx+8ySbq/x5QL5bPGeB71WvUKdWbO2rRHdIQ7S6wVa
1HmYZkrfOrrkcNW1tcZNfzJX6TgK0+Id08HstBTbR1v98IxUaR1V/IQi816qSsXy
3PTNuJW5vbS5K8NmS6td6TT9XqsBfvfxeb82hMIM000UY7v2P93Bo+oZCNUvMrPj
ZOacjbE4KgNmRjZqT2KyliySAVRDGb0P/KfZ+Ed6VXLlHA7/4cFaj26IKCjUXqNX
zzwT1tbMFnD/XJAjsTJN3zTixyRLisRSXgjCY60fgrZMoqYQQ5+9B5q+oaOc3Scx
tFmBXQ3YZAQbRfmOPyhU0sHUojQ0Th9ivGDY8Co+JZFGReAs6/jsri6dftEcIZK3
nK3ugk+O9MF1kbDterEtNsz9bUkvGhtexoKQMmpL86hRdO4L4f8MWNmuzQhyTrUR
PVbyQPjKSVf5MJraqwJN0MPAuZmAe5dcn/+leSOjL5opxtL5xtEJIfFCkv8VeHX5
OCwIU4dcKeLh9QAUTG07wxu+6+9BJFjTZa92eu+IW+6UI9oLyEN436BdpHLV+xjy
qMQ71RsxEM94pt4SNFL4NsSz1MzfiaqVtxI+GGzIbUI25Kyj6y3MMzuNh2EBNiDq
WPMZBpiQN1vQrOAepfK39LtXhsFiRPf/QuYBO8/aIuVKcAT/Vq8KeBpRGke5L3Y6
I2xTu8V6u9i8SGUoK23tUQ8zZEnoM6Jjmy7iKYCGqDUn4Jslu4VHNAkRqkCb53uZ
7geehZDFCTC/Xv1lmxpapxgRCjKgHuwnokbaFA+EOLM1qs1uEk9q37ogwf7y/+zE
J3A7kD9Ivm8ueEUyJYRqlPcV/5WCO35ojUHQT70X23UOn7sAEGx4f+bgK6NKBCOk
c7hvM9e3eGv5lW/04M1C6y+z4bAlT/BBI9OG9WcnWjBKOfCGYbiKsv+ZjPxooa6Q
wadshkGNcO8+/aQJuOCqFGrtDu2hd1DALEXGjewEhEbagcfHw/r9bQqpjVv1e3V5
bWy2XafTJQHK59bD0bE67QDc7Yt4iOw4nRfid8JUbXY516y+YO2RS+yZLZqUl9h5
7ybgC1UJVeKacH0nr2/NYOm7S5k+oorPEFSOst863q2kBMuAqrBYM1EJLbNm8ys8
OhT1s98G/E/z3WNDLPEV8vm2Yd3ymDW4Q8hCXyehkrqnDKNrcDR1g5TrVPmiVs2i
p8Jcw8PtpbIgXLEkjZXrEPDKtBT4o+amnbRma+rOFvcL739DvPrsCzsee1WBOk4V
2HArUBdXVxZ+qEV0OiAQlExtaZ9tNOFiOdv7DwfiCDLaRla7dw21WZrWT76gQ6gP
VmjshRNA/8CX6mUVtqjEJfS73QOZ6tgRu1lHcsopLMsih6qGoESFbsRvgY+p+osY
skRSAs2gUeJNJnWor6MTw4LOtzOJqmh8Art6Hrqedpm0+QiAcGO/ia6GhM9RKbsw
y/R+mTn2LQ+WKNDWKD2Qj50nSnSXSLnFMsZgG/HcEL8hE8QDy57l3ll+qC5pNntT
4ZbfrpoTDY6r+keuSSqAFbeqLkD+pWTgnwlvceFK1x90vBZgp0gdbj6VuZY5DJpY
XEFeBM58HclIPs/9T0HaajLdN6ZU3ma5/tb1GsjhREFzmn5oH0GgtMuAyuaSAwPi
uPfza2suC0mLYJpEnjTJLF1yVNn5fbJCj6s7eCy98O0nw/bqUnemTNFNK34XHRrS
mUyAcMP1XptEgpMOfqVxhMRv+sxA2xx+mev+2YqEiSU++tovQzF+gwfM0ZJZ8hoK
I0pY+gU4O6Q3kBr/DGuhELNIWSLqdFzPDnXgqFJEEUo/iXQAvbGnSMOGnPUAObgG
ZHJztbgOJDeBAN5K3CBviYLbsYCGgV3xbkItk9KZsHG/Wx+ujYf3v+GbTDoPpRG0
f0Ku9KNmlQOErQgHsxFlMb7AFEaG5KHpQ8amfEnM4g/bnSNwkZTo1WqBALuiLO1u
l6OddYLSberBVwUOeKDXIP8iub4JZXxecuIRLNYpNAROIYgjVsJF1IHDq7NginW3
RA18TDeAzuBa8NZCLhr3V3rIkRMWfXD9Cj7hRZyTe3KgL3w74AIrxPukUR0BgFxw
JDc4NLoypmhfxpQ4fJQxoJg9kuMZK/07cKZj676JhRh2ixsTOuC4CLDmGhQLm+ho
7sk3fbUHVf5mtow16TBU+piv8BY5pJnWuGM5Tri9w9DOY+7ECxlxkrFPqW47BJAz
S01/FQgCgXNHGHBgbo4dMF+ft/wEkvOVck9XuBwi64PUXGcuQBUAj5tqYHWdiApf
FhJRQPmwSSjbJsdTl81mmcnbRIrxpXYEhrFIJuPDGhX7tyKUIweOBh5R744RNaUY
jXN0ri2wqBII9ak0iri77kSeDT8fjtE4g0IE+E2uoPfBGXdagd4rgmOakjoJAck4
e6U+/FnfJdj2Al2xoaRMXDASbX4StukipEK/f0CpDcmSlpFgMXW84CclLWXS6bcx
9I/2r0Lp7JLuulqogp37frrScKZW660rKxBzBtKfqkXPmYqjx8rTRj8WuXXxJI98
RWMgewBVAON7UeRgl6WujJhZ6XsJiMYcQ2wfGOyG15BjoyWTO4Dfy7x3gi+teGXi
qTzLdASieyvG3m71VD/BM2YnAlPqHfakZ0CJm6KOPkCCosCCXqSUTN6Bq7eU6ej1
R5i3oxSWlmvICDSuKQQTa3yDPqyEWH0gSlgXduBwRbtU6AwbckuKserAWkRSVjaB
X7oJ0yexo8isxq9rFI2NF7fyvffIxkLO26OMaO2GDyxPbhCWJQZk686Ur1kBEaHq
MrLHPBdjEgo9MO8fTJlkBWOHuPa3BV0tHhDEyph///FzVTVpQpIShOTu3gF9nuub
/2+8ooXyzbdGfxIZqMYXWsxQNFOXwOWyBeFRxyUvUbrnqjiEWivU0q37zQ5RNDGb
xY0t9mcOC7PHAuFrPLbF6NPjXwQYKZU2k3Ld29QFPhNJujeRDeafeTVwDP+2eQav
QB/TuvFmIA2FApJfitJMSZDMU5Z//i2hq0jpJgX26eIYSGeM//dT67vR8dWCXBnk
rw29bYIfu5iewUNwDNjlrH9I1MwaSUdmVASQtntc9fzlELGlpf9lkeCXAK4aux4k
0D9dzHvyuuN44Jz0npJO8sOMYKOLCXV1PtZC2PlZOvNtpbq8U7byvJMzYXrf4vV4
Sxn4y081QQsrPX9quEbczKTzzK8XvcilJex1osy9atQXzzzGflKgkzUeQ0zEE2lu
t5HcW7BpF+BRV3MEZ6nnWfv12+VBMtv0dbk2l7ZBYb/riYeQv1ujeClYb1K6BIrL
ZuuIKWuOg1l2qjvgIkGxf9SpYyJIFXIR63Xknskjpss94By/AIX3ZS1+/cSZ8vtN
fTjmhkh4+TbWfGeZEjakZkzlXGQ1Q2cmhHsKDUp72feNYuT5ZfpxwBZbGeOLL8sT
4v8RlNsqvyiiw6sKbKh1wFV/IslcTUUuCQ1Pg5NNX2Z8+i8ly73wtZqWiIzZax6c
L8OqdMkxa6RBwoy4Wx35M/YXLrd8mMIm8mZ/0XMgp/fiYY6QRFaJ6wEml/HAx64U
2kw6Z4n6Y5E3N4hTV14E1je0Ei4uVv0rcSdwzWIcmKTtMiS9amTwF11ttTRTT9xj
JeKdawMjTzmnDBieruR81+tq8adEzorulR9pEoEUzUgNpHei8HGyRormSyK2PymD
GxtF99lCKp8JOHIZfIHRdzAO7PiV3Tuq8gNyDtSj2ffZAljA4v119NwNmoJCyHNs
jcUUyjzl0cO33m5P6khZfy6Bzi1NHClRwLp0es+lavVIJGeACDFfpgKY3eawhVOo
88oELtAddDigpzXCa8kw9bidFq4CVPuWdTby9LY+XPlYzaqzCtLHjUb8mEZABnZn
EM+iEbjgs8z4dK6WPd2cL3J+Kp4dmTm0C30AtcKx3KbGalv0GQIo2SjibOX0JBsv
6ahqCVYDYtwp0WzbfUBnrG60pQ7Vb7ysuexH0xduqJG0uFSXK99d9fuHWHXqFJtN
PsmBTfdCCGKIG9aPWliEi9J+MKtLl6vMH78mZDDBZFSyTPv07Gxuoo/6phLvZSv1
idrTkE4dzw4rV5gAEG8Yj9Cw6Vmk992scF5M6BpQgsp+QyzPwj41gEVwjOsktKHz
WFbUpnBAmknwn3TuVqmKIzUMvC9fs1ZVt2sJ+WGiZLovZWsrk7P/zBJKVM/Xm55+
Y4pIDpIO/3qugWrr6tN2PWuaU9x+eTDG665sYUQHTXQHFEl/KHE54pR5ezq7+TCp
yEg6BpRbj2kZBhgaCvHEnOQefnX1URtFiWTYcFxLN2KYVsAfI5OTooGNNkb9kgbT
jKgCLCDVAP75WdNgcL2PCX2NkFbT36ew38t4Th26inI2c6fbsb6/S5r/bOF0uz9O
DDwLxYVFYyW0K9dc0300AtkXWNHy09HX9i6G8gRNFGr/v7rTSV/SevNvSfFsmUgQ
uMYFmSyyK4HDciX3yEr8rC1OW53NBKGvoKBNc7Z6dCi6kScALxktImiUUFHfcl/G
Apv6TtMnajoZatv0XQOdNc5qX7mmRKDGT++jlZ+Zt+VJFJanhNqvXSD0VgKHp0Fn
gvjg6b2vhUQ1oiZDN+JcrEdhE5hG8qMrM//UmQIT6B40QJcBzlFe6cDdsrYYbg1V
h5EUOv+lH3dzReNZTK1GrJzDEbXkC53Ieu1yimLd0fQ/diw/1xZiVlb7QwHebOAT
06e4B3sRc30gKNSz5nYgaWER79NXHwBoK6OoESwxJLxVbxzhTdqgAMGjbEtnVwY9
uxkDxBmoQWTFvqOyoHqNTqxtYgu4oyEWZUNhk9XzGxezJsekE3dc9jkdzmeMXgjY
/EGYASUDOHXfvAPCA4YZTi2QkdFW48kRKRmtTvzx3rZVXVklmVTLiGNMWrZ2bmzF
ErqBWa8oP/OeXmx5aFR3RIESXUeXWrNNFZaSw6qHDyhhh94AtwFOHw97Ue5k+2zB
cmRa8PgcHjEjhP3c8VO6TU2EsKYO4IzIOZQkws1SnJy1GHSeYczohucBA1CQeQz1
gm3lU6cn9EATSXBxc0xKSUROOZqTAy2AWzcxLlEGxhN9EgfI9hSbu8BlrkKsVa85
KOwQ8q4+CCWxbt3v+2DrUk8CdM5qOoWMNYoiZoMh5AJZQH4bo37zK+505cvoJwY+
Mx22/CW6hLREmFEHerS7fYAcpagt6eRsuRxCUKFSjL/Ny9fsMVIliT6MEBtOWLhi
Hnwy9OQotOCAck5E7pik/BvPcqgzE7Q6G1wARUAz1t/kXoSPZVZZqTPriTXx6zVL
NZP2mDdOKeT142ug3o089TN+2mdZ28ssOodtZ4stB0vbunQhhDYsVGQXc/KZZEoG
5PtndW1v/sZC6p+CXfZ6Wg2eZWokZvGNthmtYaUWB0ts1MgtYe6lpTIrjUqKyMmS
UQ/dIvORC1PjxikJZ6r6fX4zsycpEbGBku0A4q2qMWa6lzOQWvVtWMhSDXYBAVLd
UCMHQLh8AUWpDaROIbOK57VPhFvRfVB3P4wOw8nauwc4w/Pu2Y4EdWJZ6neYNPui
wvDavdwF5TE/imU6qG3XzY47lzG5H/jnNJfOAN9LhyUvlFpS1tOt8gmlsZoU4nUA
uSZJDrgv9txW4MywXXDTuCpoEm8GQYYoZQcyZ08CfbC7bMhjHj90R4CpEXSye0cF
ZxKT5qCuhXwb4KZs6ir0fNv90SbwCSYCZRwD5jysOCByccFHhQ4eHza+aHA9/N0j
SuC+VJeZUdBJ/k0obRTIA/ERvTAhjnJcQWW16rHBu4YPqaFGpJSrR8Hk4hF+xypb
Ks+HwD8d5w7vIjrhSMea/YvJ/eaCIdt5yPHZZCEPLuYjXB+vKsTtiBjj4GIB9rn5
/D5fqEsS17/WEU0Y8uIn6ZImlJkniMNZs8h1VU7+Gt/VL+HdMuQZMTE44XEqZK+j
U2FsNdgAIVbZvsx1BX9qUPFML8g3MGTFT+At9vpKspAqGzI7L1pzqfls/rLdS/ZA
bXXXzfl0Fnyscip2RSZxGBNQmd7NH2e38ARh1kgcyTXL6gbKKENHeuGzpDixZ8c4
azPE9p5y2IW0IvoLTVNoGpITmILZHZlODswwip2QNMeLb3N7iLgkMhXfy/k/yHT0
3ujOCCJsoWRRAVSvx+6DjCw8Z2MpNl/1XtLYXlBFlibfg5xTNmpTrH4sZYnZ6W0u
TYJJiEF/NdTUKL3Pu2cMiZr1B2lCIMOTlMtOiYk8eYVFrappcCIvxpq5TmbQdySt
5297wCz5TDWCo6xOVBiJFnF5KJfCDAKFuvmlnKg5V4Yz6ia2G8zL9iL3u0KZDD+4
EYkSBFYHs1w71ci/YKSbM3ZmYh/ppEQrVjLyPw1R2GbWE+Qk7eONDZL2TDrk/P3q
0Tf4/MOVpCZLYWNa9AQmQwI+m5/qMFSiCWxxXkWXXT7ugg6xG2oSqQWGw8tPuF38
6DF46yrMp+uikcEPdZamBySBBnjcktfm3n7y6QpBgB3zrU/nkyLjS96++dcxdzvk
WyzxD1jwSu8i75q7Vt+T/sAMEE3uZRmxs938bral4uRt362X+5OhvZe38WQGkJzQ
a/W1LQU9A2/i9KU+HRKezLB/D/o2ACD0UtUsUTfchiFtvD0WlgnzeUhY5366eWXc
dze1w4Ei0yOfI/vsf6OLTUQYKPGdWc5TI53kTV2svDWzyPsujrkr4pC3JXPkmoqR
2Avs6bxS9/DPO1VZsAUCyLPkhXmTY0N4gtwx6nOJZXm/FgyiLARU11fRgwfIjKn6
MI4itT8pPcIHhKOTSqAd0o5CcoCnmWgqUsOZabw0Zj/ZRhwIqKE6OSqeEp1lDzx4
7W7EAU82gnRGtG3Rf5PXGEp4KMXH+59aI7rNM68+LAKQPBLGcFQ8AjCJajSCDhhr
nHdFnp/kWBJiMIyQzm2kntnhowh7NkclvCWFB0GXREEwOYj3izjzh3am5qXb949P
JGSfTx60MMoAEpQVznw4U5D9xdXU+9ns6dQ+795kgfCca3ORiP8gEKY+uNMgfTIS
eaLCag81Oqm7HPj0DQ/rAXEDDjNOPISZBLXEyL3goW2XFx2Af4h/DsRHnWSoV/hv
vQRue+XncowfIYcqaLqcY/DS3tpCQWwj+G000hnIn4R/WUZZka9BBzKLr8bpoqYB
xxilYmZbIgF6g8S9lNYkufdfdG+q1mEuixXK9Q/yP8tC1ICeZ5fyeWtWmlrKEsFz
teua+VekmyrQ2EoZ2jfwnSJ6FUYvcRcQneVafeN4DPcTKo29+uHZ8CrN+RXseYMF
djapSRaJKjdBEh8ex2AsXMaI/svZIrRmaCsy72tve2ExVCv+krJHGGpvoR+0+TuH
9yEUr8jtuEKxWYnijzfys21sXn/Z9FmJB0RAdtU7hOYOuKVBp0Ox6Km4OCU4wd4J
c9j2dQU25RHJ6bKUI7DpgtoAXsQgeIg4wLUYHQGvPseJDYpjWTOSy8mJpvjwPqop
7FG4w/cX3/LZ5gesDhn0RDn3yU2woJ1irJsw+crT4eFk6MZEgDjtFxpL3fnRAh8P
hFu2GTiYKGtZqRiyeqS2djJosrBBpeZkrRPvIVxrnw71FB/NpdHTc1yNkGpE/7z+
PS/NOy8Vvto6SqM5vJfwAy7N2dO056A+T0nOUnEa2EWK+TC6/e8hiXoi8SbVj8sy
ipk8iUXdpxR4G+bfFSZOMm7YntzZvkfpLAPMoTITm3RK/cU5taAhDncahV/YT0K/
9jw1ROFCYMeisv7JA8odymZu9wBAGGk19KOIKUFRbb2ETHuf0wa4qOc+74odcIkn
Lgin3z4c7EK0/0x/yx67s9UAKr2nq6yKxRabN32gJL08unLe2pbktt87OluMrYv2
id0UaatDQ3XidT6LS/+YBZvhHImj2n6yIdZRLyrmokRIH4r04Nc0JEmSF8ty8WT2
9Nl1lBTbPV2Rt/1sCNiAR2sDEWjMPumMd6CynZP9T/haQulQfLw2i0bpqM2Q7Ple
5CTPRpwOGDdfpa29yQHQIrK9KZAgEjy/oWAvoEsPfS3HM2eoVdd3KMz15JUpVxji
51tiKvS7qfnpUUsD20ks5ukDFNSQezWh+Vz3f4CXqzdIwPEvymPyay8n16jpcR87
3x4mEBvQAeBDBDx2p8qI9IURZbToA4YX9VMZG5zNpDtmTbj27OqFQhc412jpUvIT
X8Ig9Za3zZs1tFc3a3zmZvmXPfxcRggNmdmpWaaJemLhptihZ5xwVY9coxpaF9PW
zjjzWgILl8hKOAIE5Fj9wdIi4+6o12ohnctMQiGNaZavvNfPuAcXZRN8Kekd8YmK
zExvkDkn4016CZz0xV04PR0RlXN3aNdCc1X6ISrv4cDG2e1glmhLide3f/L9g5+v
E4V8djgtMDGgC3P7ClAlzpk39lXU4s9dfKsSl62KvTFxYvh+mO24j0AYaOn3cN35
O09sYNCzECVoMlix0xuCKPfcImqk6shwtIEL3VnDKAvK6dGLMtIIc1RX26yexT/Z
FIaxnySDtfOXCIeFFruPKi33tpINzddnR5RX8aidcOeJwKnvo5CyXAi97i/AC4fg
9PzMfe0QQ0xv2BWqJgmiVO/H0NVMcrlhMmouKbOP5UUnErTO+CKzRDSp+rN6cJ/a
JZJG2uMEZAvHPWXh/66ZEhu6/39BsSNkubgSl0f2sVxJUoMEmUT3vnXAcX8nv9Wo
mQ06ULIEV61Li0FwJR64G/WGnPwGLVaWcmr3WivlbNm1JVByUdyN1CORbkFk/DMl
o3BwjtNlTtWYx6MxAOmhAauwv2iLtBTHCLhzGiNdC021nDJPvH0YDWvwKDPNQp01
xx7ju98zWjIEEmQ3H0IXqgIun7gN53kkfX39tRrZPgTgA5xUC11YbAoZF7TyU1Vk
IVX6cVZ/joqk1P6zLQtIxHbHZ2fLVrKHm/SdnojzmAOqq+j+EnIWlSVi+pxHbAle
QuXbv0DIeJrUyWiW2UzgVyhge9jAMUro891itLOupEoMWFzTAZAK7e8+auLfgPaY
txiauFMRN/vmgU1QLTi7leygIOx54ATKE1HmqgsaUZ/aMnvnsxgrZxBr4mJeZWCZ
elrtBOoAzRgPJDtAc/XrcUHZQaaqRZ97DgkeyToxGcK4ZvkblkvYEB2xAO4AD8zN
bLwiFtkLKR4euxSkboNh2eaf/wKpW20PkCs9fj6cXFqSZgx4zcKfuadrmcvi19xY
xGWnUgwZnR9rvhoqMEDiO7o6PiGDNphI+Jac52FeLDSWpHENXrC91wSZnQIs3Wn8
cva7MJYzaVoDYtAiATa+bZCzDryH3io5ojfPrvxNdlpxGfkcF5VFipdpdunSVFTq
0ciJpoG/4BjVIfQI1a6SX2QsAG8Oo37rbZ/wQ689Y8buF74IpU0Ufa6b07ElDKRW
szEr/Yw5f5mnX/XGi6Cv07nju8eD8LV9YoVrt1kjKlsFnlqcUfzsexWcoI0znNGH
dyFnx+f3CvWnp20mz5BFqM9+YP4r8inqez4TUuZ742ZPNZNUWPgQWjV9c0o51RWh
Aqi23UnKXyEXQ+n/nN4t7tsyrlVwtLlcPYMDf447hSOqdIbuCUus7iKM9EivfreS
r61CX5WKdXf3RmIH4kO+Pb4w3M4cNWmU1Ch9vX7QAJtvMnif475sQTmzvgboWx1Q
xgyz3QUZghDl8FRdNH3HGjlNIWszGKwXI0gH+vKYtpds3IkIdX8f9m4UzIVlFeoy
9kBJLpQWZAOKHRtkozK4P4jKqfwqljIVXGpCbl4Zk6OQsFtaI2+WRPKcR9Ji+sAa
ZV0zKQsUiaA0LecfUt+1eeW4f3g/rWSYDL1CbJ0Fp9auU5kJlMZzq666pNa8bjD5
0SKGZwladqf+VNV3d0tuN+W7Q4q0FQPOFmClHemiDTGGRslyU0q6dLOupJogtM2E
8ClwgjcknOVdEJ1RDU7czNtDaAiJPgme6IbGrPx3QeI0AWKicGBbz/kDsRcPUWp2
2DCfC1EOcrx39zLp1SvMBdKkTK447cH4/H5SBkKiWujHk/Ou6L47GbQjB6cx1d8I
MsWiBu6QgS192U7XYN2Ceuml8xUzM2y+/g+bs4KwLQb9fCRHQnOIZXbFTxOMxBUW
F+/KhSMKT+QuEpa2tSiOsu5Wfvc4cqj7cS14OnGDnmNI/YSUnwuuLIT7Ppqk9QgW
afZ2tKOpKrhmKSwpEgObPf2hWhJxMhaFgjM2Qgi7NNIF4vR9cQf2ajSbpy3u1qnu
/c4bFzJAYhOAcAE6MLyUbaJZZzVvQmLBebDJ4WPr6JzOMiFg8AkqCbid414LIkKI
b5EBLmGyLAFRE9o34Aknhe6hZqITQuSLU/aCZCu5lepnNlCRWa9+OtUI1Otl/o/2
UQK6tgWPJHNH+S2EsThZUYNGWgPkPCS0TIL8f0e8Nrng/lUy+1sJ5esI1pJsJZ5C
TA8BsZkUOLrjTDzjDIOR1UqkkNY4FGsYnbJeH0uBJojaljzZ6HetJIDhR41Pe3It
AkCjB3hGQSHHw6ZqUE9YHM8PyYzGkGRco2GZYha768lojojnXUHUIS0mMI5u+0vL
FAlMEyLbGq54+zp7LidclUVCwmcNwT4onD4D1nfqmlN35dCuHZD/iLWo2K2cX8TA
Xv1nTGW/OIfe5Ker5WYRzj43SXLFhOLVf6TIzng5997FuMc8WFE/xEXaUewobRFs
Z+kO13zaCBMqZFfUFp9CX3qbL7Zw4DZzWAIkdw8IjSU+dQBtLYoioop4ISpIQ6Mo
CHIspp8RrEZPCeBbItULCp4l9MnEqXb5ro/4iXanvUL3bjEzfwqAEmhhHtZ776Tr
khqz7nMJc2Rc5jr+pjnDeFO6CTjf4MjVYVZkjFHaMyORSqvm5GZb2nriecwkykpN
c3CNGT9vjm+2MtwlneBYHqVWhw0568/wUdp979z8EbZG2ZE7xuIMcQ3YFnLXjVHX
VFfNRaqtdvQe/zyt+6/dGTAkBFJR43QH0hg0qy5atzzwwbcCm6Pf7uXuadUak79+
xBmOmTzYVwX/sNGmtSRQ8vnKwRBdxCQTIdfeF1szZDI5wmaYc9kDqQzxHdtUeVJh
25mi+utcBZR8ZNw6tgzS36DeymHZUP/AkiILtoZX5RRSVwA3sJSNxPubL/+e2OpE
3RRFI8YKF/JQaurpsrnChfa3bLhKSL7n/SJa0ptKP3i99vbwWROyirYIQtAqbvDL
xiAHUiVb1vk9V3FXDfZABxLi9Bqih/ZQy6PpmFNN6bJTr+qw+gncdiJ3+jM6cgzE
cXjZhm+tsaVfQuOShkynC3e464zv7Rc2U4Mj1jw8g9oD2tMUKnH0qqu0Ni9pNstI
a0LaFM7YGUfgCMaKiyD7GNLX6bMVVQlCuYUhN0vaVwpUa8nT06b36eLSrzkX1WiA
Q0fuTheJ+Lsbw+lfeu4au6iRJtp6GTdanTcQe02CHWxXQ7Oe/L1BSiEwhSOMHVcd
FNstVrgRdn60tLaGBhYa70YTC2UdjBKfjv0mzczrI0daLT3uOQFH4k4s/vncCwN4
84b+NNm9BKkzeopDKvlvdDIsAZiOC1XtwwtsunXzpzstLdHnekmQSWDKo0EAMeaO
qdF7D6e0WRgSOVMBIJ6Ny3tWS1vztRw6q7DpJMpi6hXcxzzgWILu0toriE/MSgsO
/sYxXebyl0x48PIwurDQ9egJwNZsOfWCxgphs1mk7qGEpQ0tS1I1UNSgZFpq2Q4h
0qzAUUkk42PbAmEoZMkE0yxb62Byn8tKVf6cIPOThtBzfrp+DAOwYb6waCL/Hm03
d08wIVfO7rh3Xb2h8DUXdfMnCoqJv56lmm6mDt/uurnkAmsjj0neBvTiiGmf6K8X
adlcLxrlVUHhOoEH5i1pvefcqGySCGE8Lap5RVvbkhlf9L530ndsODTjBnT7c0P0
bnStIwY2dcOl6RdIixD63w0Y28CbgPDTxKTRzhJpsZbgHhW8xOHO6k7vqnfXRi+3
9gtby8Tk3MsPqMIdj/DovxaWxjTiLS0EJ3YPceQF6ZFkllPUETxsYPYMCBVk3RSm
PYK4ud3hdNaNkEyHLt7lO5wi0bsj9n4lmoRXByw23QGh3+5OyPD+u27xkUGh+hgn
ANqy1553SQrRrQggD6+Z1ISHz4Wl9/UpsSGZntcHyWr6igA+v/ngelAd+rtdDPje
sQrMr1OU3J1KOcxh25UAnoNosb8M4NS2hTMGe+LpljN4EKMOuzkokuhWMXqkaKXm
BKE7i7Ed1yyDve1Y0p5I21BnaTSALVoufVaX6UBEX3XxGHoIb75lz6WT7tCQNkSZ
HG/ouCUUsb01i5xYc4XPLTftBbdgWo8nVVV6wgg+EHs4S8PWXuxQiIwtpjIlhwna
nEAmmOLiC/bnYThAjwoCg/agu/A6AqbU6GKVU5klMMkx56JdYQ8NSp2U13xYWPij
SHFF/cM2cWUodS8hbz5Ssdngr67TAP6vw2w+GwQ+lV2EZu3oKYNbRkRVETXmgGGV
Vp8TTZJHBHRpOapb5Jofk24KUvUol7WpSbV7tteAcGiW96lorOBmBWRmukUVpjmy
JO5RxBY1x6APsVEtmCGMj5hNtfbKz8ug/haQXup6eTyfTPSp2GOB2zBb9mfytNUI
TRlVMSO8wcOMCfjTMx6jrkQ2aR++bu30aoUR2lnasO4haVSjAzYsVAAfV//Z2NEz
zGyqle76gxk+9kexvXcezhDiFtxK7yQQCrZ1qP9H3OY46bNZMQQZjChEK4pt0BdC
vfER30kSZwZrupx3WFnxrgnxHoYo7kk7ixMzgiDiWld9B4IHa4D3cKVknr7fkxNu
nmbTToBpnQBPpOB+GWaVyHQL99XFn4yeFgNHs9JP0nvLvBFEf9DwGfkpUTWDZ7he
i1SXmo2d8Jjo+ixZ4DYC0aWROXkGPJvO2p1TcRg2htDslTvRKxIR0EEM9NKFSgOl
hwl99tKNyj1vERbzxJy1EA1c909qkkN1frHqy0CrybIl9d7OQftj7ro5k5dnch3v
Bajziw40JIJ7+k35WVT+hkKB4xhzdu4p+YHVEWM4U2Xdht8oZNjRZbE9tbIecxEe
FaxKR8uzmg5EhpJq/3KWMOmo6DbBGumBeSSVx25MoDkxsaxvGPtZJ5jFgNJITCMZ
vKU7DhrDmyMAW173Jzk70DO9MV9d5kdT8nLm7UHqLH/C1D/HgqZgtozME6fyHS2P
0y2Nb/XrrSQnv717O6m6CbLi5Fz5UItR/HpUe3YZ0TOyN0bU5k4jM8ltVSADJeDG
DZm/g1cBxxbAtbvYZc7ZOUAN8HtcUTIq0sVg071RxBF7vzMcCoIFN0fGnpSBRiAV
vm6di4XonW+xoBQZR6YW++a83DDRVidtoHVYcyYYHUNRQSZpjsI7v1T1wTaEXkzO
jDVx1DeTUxZwePmff1C1Nn/EANdmr8pV/ij+Lzwp23q7Rvb6p73oPnYU3/HZyVx2
KK5BpDp6/rotArR+qgCU7UWOoMUyEsS/2MEBEBE0FGjiujd6ojjcjIVpI/jng07b
Ih8W1JdsFZxE/QJyFm55yZHqnNlcdA+qS70RYu6QWyVp00NopnFxDHfoJCrAB5M/
XY+bsASeZqFWF2QT7vACLQnrPLkYkJaaEDaZZbs13/srMYLjsLemUHAAKWtR4RNr
/U1SoLG7qsZ08VTSfhXB470NtDT6QkoJNof3VBfgE5/7oxZ/QS6pJEHkRHs0uZ2+
pA0E6QDjmYRkRwxkwRRBf5vVC+MH0yci1egNbu4HfbX04JUPbg8gAahUoX05U5Ge
WVulJ1UfUtiEwpOZhtUX5jSVRxJrRGzi8hjzJCNymnx+BumqUdfZOq+RO66DL+Pf
Zo0/694lIaj3GWBL56k/W2zTjLThbrUzEHhweWRYi8MqvaYSZ0kwRhvNuGnVGK0I
3LCFdlTVdHHcxQOiboBBZPpMm+7wEaY/QJEXg1UQzyorvLOnxjzMmoYMz1wteM5X
h3V0/A5D654D+CD+lUeCztlXRnLz8mVMnYLydqcb6ejVKlAlhYGYDAVSTv6t1ksm
pP/g7vaG+fbRY6ZhF/C0umghA3EpQ3t9RxgnHh/AV3ynASlygucv9h+yayvxXNVn
pMIfNEbGwB5GjbPrUtOL+CzOdXTMCgUm6DDvmrhmm8zec+EpvBy23JZwbjfAKRd1
HbsZfwSm4YYx3L/UUgRwvnhIQd4ouYfNKZWHu6WSyEEo4wdlTKueVbYLHXsMgYzN
vpgE/BLcNRfEqRXCsEIXGZQPzKvAwH6cIhcvyI267kZT8VTAHK15wDbOgShpJ9cG
ef43ZrF+n+yGipbq1YRLjIJDCa25Xhj9s7LYh9UNuzA=
`pragma protect end_protected
