// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:33 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IRmGUILz4TAIBkbAL0Jtks97R9KPUrXY7yenI6dFBfvUmxwxGkSmG5OK/Dtlw4o+
lh2F5yWmyZM9JAZViQ5FrO5O/DvbmB2nyRFnDuO30LMym7/QIyx28WIOpUhRKjWG
4NjD4OeXlzfXOWU0NPvaCE/6hCuvl2q9CrwJNh6W+f4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25664)
bNWpA1c6tZiYyeJ5MynFXhJZWhcHc+DgTAaPFK7mA/g3qL1AcZHEean4EUjhlNIM
sZE3VHC2mOa6L4tayEBM2QWZoyOy5Q8qWw+ylFYDsHeXEtvV3MEqywyQIkF8Bj4T
p838BdX9VTlnZ5zlO7hmEupAIxfLjNqRqRfbvIPD6B1v7sw/svwa4L2reP739IKp
SGsLtmFzO+uELMubpj0YErvaTIalh/lrCqKuTzlrTqPAHCKRmc5Gho4EeYktPtWR
BNnher8wJMQbmLSdP4bqF/ys78hxrBYo48jzjK5fyttUwsJFKUZwIgrgsefdsGJy
1qB2mZQt6xWME8G5hkp65YxSEy8x5Ib/zWYdec2Q1j0nK1tCy6DJKKPIdCE+8gt9
Fbd9O2ZHLULR2t1f4fQ8jaL4jC3Tz/3kiclUx69/sFYhlXflFaIYmFSgXTGlpkJs
HKtDq5my5blDx9FuZnUHNyupmGBqBrdigeNiyUgTE/BUQmiw9kjKqU1MSmTWKGtW
rat9xt5M3kjIenQxCejl/XW4wdJXt0aTsNGRH5ey20SO29KrWd1OvBOytOubof2I
g27xsomlhD7ANQvHg4QxBMSsBGB2bvmwYnyxVND/wIcgZudvTcKWzGE+z90APC0g
jpwZRoKpOast1JR8Vpr4bbj77E7/MGX713X9w+cuqLGGYG4/8fFYH2vpK0Ztc3UH
AjiGf7ootQ+xX/YbFsRRTJY1Vd/7/vGN7hn4GZmoPHXmkuIzTsPbXPE8GW7ZkVE7
p8v+ajzrdNxRfzYAlAaNXkcc0C30DnHrAt7lp9pp0/QEgT+CLFINxmLuMdbhJ6Ur
CriTmQ9rIgTJci4b0NGdJXYh2WesNjDuonHn+xXNhvtStu/fPxhnvRC1nJL8Mvpz
NBfPEyW8x9AEi8agPEnXpYbp5s33PeRjNz27sBXkm7wKubq86qS7dx9RWHkuV6//
gbqJUcyVBobcEjt499kef1B6g7CUKTu+Mqcc0dwcfNNNgqxIhyKZx2Z5iNMygi95
NDBoX6wyONGODmnOvejW3M1KNglyKPg+PWqLCSfi9sBC1N5xOQD+3KBHjdK2dCYD
pSJ9+LkSXRFNN0rf/I/YAjRqryt3RyQV73L0xmpcesaO1Az6jIR+Bb7h3aDuSKpj
zQ/SNgyuGaJOxDEKuogFjAwfBcEBF8mHyJNBRrTgdR77LJps5nSbCjh2iyDB6nhc
UTJVW/4xJietZoB+MlG+lo1CFnRgxsW1PawHJQNUTrLQe8/8V+rH2bM3Vcvb8L98
yQQllFGpt/a4WBDMjzUvlj/HwixU9W+fN6bEaYmfuXI8MPadxmRe+BuR+26tsH56
CpmD4JApv/h98HT/4kIiHaHv+7IL9E/B89uG46QQwqjMO1hq0URCKT09JD9GYntk
nvGboO6FYtGvDsX6mAd1PhT2cvGFn5SYTJIllUhpPURX+cEuNyQQQyqSiHz2OX/A
P9kp9fWYbkKB8aG/wRQHAqG6M5iiFFOYLdc3SlvvuMCz2IoWAij8e84PTPD13Yv0
HhJi8jcCmeIlDF3rMBCFtsZ1sy/0LH7TER9UMKBWoOwt8ZCPXM7zM777SU1b629D
mgW/B348cDxEscf6rm01fzm7nLbz9Nn9BD6/FDf0geHvy57N55lAo3+jgVjex/cT
FuZAEjbjrXedq1ISrDy9SrQZJgwVYhMIhSCrmQqli852Y8mh/dJTa1JiW4ErfE6o
RlY50CbLCuVmn/+73QiD+Fdk4sc5DYIZSQLutEcnXSwRTLKvAHgbLWghu8TlPxWD
hrayz/N2Vl4GplLJ9uSSb3HLavrVn2Ex8AzLFpW00B+boOMgM0C9/Ci5SXt8Vw7V
9wKoUz3rx0zVHY6+eGxZaqSAoYJmMchFlIoG+h3AG9NvsarpbwsqpxgEvOVueAER
hlGa+m0cQ6KVoisz0Pdb38662LzuC8Flsc2HH+u05Epgpmkqgr/h55hmj6uRppjL
xovuq90vJAogqnWAdmq9Ukh5qZFcwI9fc99dahrg2D5+DoUZXOM1Z23PkirbEY9I
iZBMllXISHTjc2g/Y/g8yAf05Ji6W8BSiOFCjBNc+rK1XUC8Bj43D4z4nybpbBWa
6gTIZkAtRnGWU7zQ2PTBU6DumTUT4k73XbyiCV88pS30ZFtZO4dB4uO8r4Z+UMjp
i8B2RFhT9T+BbtpsQn/Nl9TVQPgIVWEvHyI5Wzs4bgSaIGZoV0iFb4QxpMNsVsAG
yF62PPR/9psOBg+8/aan6G5MJUerigkVvaMK9G46t+zowdqxf1ZmtnEwO4KXF2LJ
CwCaHsdVafF999bLB86QrKvJQen4YN4wy26jui6fluTdrRO+HnMdllC8JUMNw5UC
ph1dspxeEwiNpcTEIEtIAUN2jjG+p/P+mH9vvdRw7OjJsYi6G6p7J57sMrQvS0tF
7LYLq07mvnfE3Ihod+WvvfwHV7n2IrbyGE6gHrNo9GF+KTfj9hJZBnAZzrgGFM6I
HNAhr8oCmcyucGaQbfT6/maFUNEXS2xGs2WqdPgZcPdMLTtaWj8Gr05ROpRNxFgr
Sxsbo5I0YATzGsiNNO/rKG1Jm7cxyCD6M4ZvvoEna/HxsvMcOaf2zsYscHbwaiYS
Sz72naXVWaXilh+lhx8tvJ2iKlymX+1HHjDW47HfN5Do2bWS3uWBlntKzzHB08BI
GcHvcFGbx9GBRMGO80AdeFqkjyu+vvsV3KYqgphblhxgePuuQvRJsS7mNtyqBf9H
T1Tkf6X2gfMSTuHXIiwpaN/tvQOxC3eJy6fFVPv60/jvovkRsmSUpsuTYHBFvC15
qArYpNdN6hWHr5GH5GHlbhKPgd5ETON/hXPoWjIXzrAauwEOrFe2dJzNBFYt3hYe
lpV+TRMCm2tUzFtwN4mQldsvespXJhynvq0hz+twoKo081o5wXW0JxA5zK1t5swA
N6xnxbqLKePnsZsa+hAN8vPvcHbIzUMfW+EFLEMRPdwaaQIlZ9xzHgYtxk5nJK9D
yqo/78zzLOepzA+4/2aJo5oDTyx//RsSc0bbVDDHaJleyaezkFESPzxou00Ue4Nn
zrYrC0+AiDDAJXnc6xvB9ZJv2DS7hoYnbV7r8dgKLv7fh6MwkmVcxNUYROkvtdUk
16PQTnnlv13vyHysQqrkPHxVVqPufpWhvTPjFm8ePi2ViWZljsJL7pbbBcf0RStA
uu65LjIP240gsCOFbXAI9QsE3i2kzZfQUc9Oth7C2jU8X7QxmVI9BRKMJvT/P/Dl
N3lho+vuMF/JMhUu24Cy/dYmWc6uwih+FItUVALr04O9TFLTyQ0msvO8ficd1W45
0o9fnbJta4jhXtQHod7tVQPTrc5iJ7eaKNN5ee5pCC4VM6AMsdkA2JZAuIF/5Lbc
L1Df64zS36Pzo6wgjbxZ7h45dWq8yn9/FUFSWF9GxP/2jheHe3JQDslxRvit4ahp
hyFwXxh73FmBBCXI2Qn4BJXrRT9E5xn+/sGRhSrfq+rhjeCWVTkfUSdGpwlaxYif
eWgKBzoPxlU2LhNZAvSSWXJy1lNzrCIx7Xd2x2MNFACtmbY2eaRAMY786CxNZoZp
N9/XH9LOEIxBjJLwKy2Dq2He2Pd/ewpyUgNy4gnCn0Y9e3Jl+9KY4wI1morFi1oH
LZ/Cx1fkO7iQskcmX3ZUsFCA5xJDSI5VUDlVZYVixJGaDijOGxK1AwruWbg+xGS6
wY+LG7ilKyCZZmdZ0EeJvjj3OUsABkrhkAM2uka1WOvhrRiFxKECZZ8YL5b+i6Qe
DATb+GzVBvCidrVXTYXLaYfEjwW9XTRn/GsjWG/BNapowY8Z5Z/43CVCUvJQG64B
5w+rBoJdqY3kxzqcBcRg+1+zpT0VzYc4ZIql7GciFbz1OaDx7oqWXNn9cLV8koE+
go6og/kgH1Id7nqLsfWuOAz9ibnY1Agt4+OKp59LhLDRW3382JQHS4YrfOztdPzf
LOdINgmVmG2A6r1P2tRlxrDiBw/W3Em2LJlUUla33/HmYOBjtrFfgTfE4tt/011S
UTc0coVt+2NInQG6wSARcTNZgnlHU8g1AldvhhIENgu94Cq96lDQKpkSEhH3zXxU
LqHjRLZ0SJIxOFK9ZBPSliDpI0Q9r+uxsL4GRGyL5EtZ7OJeuFr27InsxmqcscOH
yPEaeZAfNYLvDIFfVZ8/pt2toAHEhw/pXOgq3MPIywUROkFMDqF9aKZnoCEIyfdL
4Dgli/eHLXmsdlIj0IT4J4Nr9NgyabRiQh0HuBrMzDSAEm7LEpPr7g3qGZhahsCV
Slzp1dy4o1zU0OXN20zR34Jn1MJIC6W1iWO92duJv0+tgeoPKIbbNTf1KYtxnKfL
6f5XJTjMjnpIMCUN8HGzxN6oBdnjP15hgiMs2kmjz4lfkX1q3vstk4fjVEsSIBCP
xRJ8qSfQ/DiNjFMflTBsYlc7CJytt+Ax9E81IC38nxEy0DAX4ALZX5CeWrbAykwr
zjcUlUuMP6uqVY3bqndtU2puwSW6fi4qNADuCryknojouWOjzXn/50yLg3wIFsGP
BmZhxP82Tk7GsbfZkPmZGhD3zoXcoBtcDsxeYnTcebJ9Zd77ggi1wg3Ec4f3PxH2
V6xrJym+Zh4ADBgx4raPh8JMyoR6RB7SLUXjTeseB5LeQMI90lcEGGRU5PPwCgeo
f9XA0AuwZyJqeEFYGXGhNofGCBzNF1DYvrF8ku2c4tPCXOxlWlHh3ZCGj9WcEKS5
mJVKMJfUvseOdXWLX6UsRUvvOXGpHbprQxHCJYOHnAuGOh44TYh1K7jxvm2f/4U3
DcPN3Cge9zWLsqCXoVjG3O4I1Ki2GfOESNz4BbMvb7+intL4nFeUuCIM1jvGaA8l
0HXbc7TGgkAmIiICzXbLA1u8HZNDhfEPETbhXasoWZrngQnsbiPsSjNqC1DwjuNx
m2RrjmIvmV+4p0JHFUXh+b0kEW+gyRtWyXJK/mOJvXKdXAl5ePuNr//CDvCcj18z
ZevGIbV8QfoUSClcbAhhh92DzIqncvnIGekp0EIgtynGlYyFUn6KKBLJktURYL0r
EN/M87ghUSgwfKtyxvyby8Frq4FqP4iPVBj+VjJiy41N+D4DkIDGpnoxjEsR7g//
phb0PvMAFUuarNQWPJYRdB1b37gHisJ9fZ9qGD1abwcFExhWYUVxr6HAAjoT/wM9
QjcvIgAO7DMIyCBs48wX+EGooAnkNr/eT1PNl1RSfa9XmJ+qeVYTiJ68z1iljfNm
dk1LvJL9vyRu8fgPn0Cob9PlzfsP10pYS9VVl4f82zMUb49NtEW2sIjV9lh1y3pJ
/42dmUTOl5f1LuVgsOIvfhzgsc2XNx4MerhPSqKSl10F8dqTs3yPt7iUBxmehwM7
7m1xLLcMyCilXO1PozpHUWv5aO8/o7IKJ/Szq+Qv8HYbaozj/djhDVUh1XmsBIAJ
PAFIK6blSwCq9Y62OMAHssxlH5Vj0h4hg5ibNEY3nmUPiivHf3/o8iKwb9ENwqYX
kA0Opjey8vAYBWzfOB3zY1yCQdUvYKTSuG9m08E186tG/gocds9XTJ7nSolBg3XG
ad+Kp4kcId2QRv+3By8FoMMGWrYx9CHTlA0R7Ugkvx53m/+vS+yCHaCn1V6A8jw/
fYx/QMfmMGDYsOIOhPUlmM9n//AYP9xaG3dKbOfcv/oVZKBUpcGWGf0PYUkYN0eZ
uNfPmONbtVWcabfeTQJPXLZufqF1bZkdOxfC4kLsXGqLundL+0b2CAAGNn7Bgdgi
GFqpjuQ7RplOH9iM2i0uug5it7A1qZ9mery0v5wH+BQfBw/5Ra+RJs/+9H6m3aMU
Ze3zJ34ChPfReG7vn0MC0jQIrF52on9NqBA76oiB/p5f3cxJnbAqV4SzKmBuxWZx
Vo39jt3JQe//UVnv4fZleZOt22MxTCnRsKY4r0VQYIX6MuCASsr+aMwiZMYJbvvH
SIqdTUwcCGV198dHl/B9sEWdbKc+Yj0WXhKoZCqYkIuQXDpmk76rwRGT9vqQMCHe
BIuz4JMHR8K+l5/6P39GBipqIDGtwPIbogBAmnJ7LpOEm8dU6bTCAlKBg46bfH9L
2SryFbfNZbnZdyPaksRgkIuLDxi9uF6i+dttn1zYF0wc3X0HX2WYRQwD+pYNhmni
fP7dAQsZ+LyOaNVu5b7WFKcnVV6z/NMHcY0mMUC29FR2B7S65A/RNTTZ6DuCQGDw
MSITGwwfe3Z+27itOKOB4wD+3GKo2UAE8njjKbbJlRZZIiZB3ZvfK1PwRAjC+SJr
YhU4OGuZB75uqf0V4H5LiG2ET9ETTKDoHk+zyTTFidU9JBtUCZ0Aoy9KWictVnpd
SmlVwOkne6ETPMJFHARZYSrYNNcbKHUNhSVmMQEEbtJ5QaazsS/AOYwcEt2So7Nf
S9ErHr3zVn9wJNTevteFSedZShjF0gmP6zkwuA7YEfiMJyQNjLvamPls7n3KSBNo
b5agUVkWZQbVjL/hA1wCuEFc0OQnD6haMyTSb569EWtWxMS2mh8Z7kTZLgYUv7bk
ncIisIolT59q5r+e+QSHlLrwFVOpC3Yy/lteyYEZTW1FjpIBYwvvsMaOAbJ+hBvX
ImdZ6yn8zWm4HOQoSrPR3A+IisfJi+Ug3KbI3hX+7REwBVQLX+8BJ8YhyElbBT6m
T2xWMub5akQrBmxJ1sCaQuVQnlBfCPQo8zM1IxgWYTa9ouiINVU2Mo5mX3ShT4s6
oJNxS6GtHSktO/umxV3JQbtmw1sDdJvacbcmEBiIltgYaNYliVwZexckW1u60N0j
Sv7qqof0BnmaVA3rbIqktW8aHNUJhegywgFgYhERtfSs+peyS3BHWafPB9XN4pgN
NnELkS23bMa8poSQcPTGEQH7wVVK74X4VNoRM+tvozCUbrWpD3klz5uHG894VdY6
UOBKEZUdhQ46LZwo1Rs1Wc7Pez03iWpswnjdAs074cpg0Sc0vaK+Favf73tI79n5
Eqw0KhVP9aA0BFyCGPPGDNn9P2f6NRwzVMvwKppq89NJ5TbOhJ+evhlOJLyhBled
mEJiKJfHXrMPKc8hNng5dx6RMgBy7LQfQRy3LbbrdCjNLqAZN9LccesMToIoW8F9
RltkBsaVeoDnr/eyJuhGYM9bhGP0UYUyolv982/XBlCP2DU8k6LZFfydudVQZtOS
sXjVBHMhb1CLc35yJmlyd+xt52vqUP1YzlMDuzbEqV/Rgoa4Fe2FosgtKNp8t8Gq
Knlr0Bt8CN6uROZFwVLe92z9KZGtlYNApHF/pSJ51+LM7GXkEAGFptjoO+ztnLF+
khQBdHXzf0mczGXid0TTNwHsFqaL3R6EzuvFCEPpib9vWDChNz70/qVcQEpIZ1PE
WC6C0bKTPnzOMfnYOBfA6d2Aaps8UAvgvVKKCwUjxIOJZk4hFWv6FW3oxrmiIobm
2G8XLu3rg3Xa1+TeAMIYhFU6fVWgTJcaHvsk18HfXblhe+ci3n5wO+jIugHF6PRU
XCgSXjI6APNyH2vgRbIrEGwEDPC5cM3lZicmkxP+kkzy0hsi0qU1DKtVOGvDBFvb
YokcUjEiDoKEYVEWON+BXhHeBn1ymA7yVeVi9MR7TvXjVnkzS3BltnlTAEy0nimM
zegi2gSJT2uA3gQqwMcZunPck38PZ+2f+yJtQ8JE5nOfjjoN9jOOKw3iEQ7CkN2h
F6G7BVejhIhM09N3JIrv8XeYmZbZRuz87N50Muc9Jv58rwye3fOx8HI++4SB8yqE
LmZZnTP4Zhy+yzq+vWT+GCPuwWw8drFRUfevgWzWLBSxQDOJOKBJERa37/JlnFBY
OMsPpo3/10hkcQQ3pgqRIvEmr8HP7EX7Yg9la5ushDIPMaxce436ALMJiQxgFa38
c4pkz/rRXXtseH5oATXGTZpdsVpoq15Kq/5fn0i+E+Z3SFSaWvRw19liqX95p334
yXEj1NKTx0sgJdWecG68HnPihQ0JInaYF58ilWvXeQM5g7peajkl/vPds+QO8drS
QfOZLACBw17NEq/C4BQt51HotlBmBebN6RBIsQlAm6WuICgEiuKoJiiovX48/3f7
I9nXDEGqSsqorMu9Ti+VafGLp0n0iVWRpFprLXPcVm78PmKXvexB2TIxAVvsySJ0
VPIKhbqUT94ZpZ4f2RcPlE0pSHtJ4tuFs2ZK6GSkgy6AxVMG4kZIug2ZXZHa3//d
/oUWEuDmr1LYqDQSJE0+VXDZFH0poBR5pIILSvyimeTqschRPmRHMRmuIFcpglzm
uOv+Wn8a76njdR+4/Jr5ElsZNgCHxNB3+lkRvg9ZlWbHyoIfHHjCnGkoCddiOETV
PwLvSggTr/agzN1PWdq0YsrPMMfx4UAu9yhpfx82VvAaX1VB92FYi+Y2o2xsta9/
wje3mhCVxYaI+8xTwWUEbm2XnzzeUTROXHMtuMVUrBJO3ifpkrEhQ6FlQDwspP4r
1GFlwGWEdF8dvAPfAAEi+aeLkXIwwLuGp58i9DnTZlf0dzX6iilRjC7Hm+yKyVcX
e0dBq/bbYK1WiR8L7qG7npwUXrpWvNAVVbQa1FOtls1SXByQ0atzUGAEmybZ15Cr
qbEch/k+39VIep5GCbbtPLuWFGCAKAquqEusWPkUqrE8SvReU446nSpw27UoWLD3
0qPcjN3u+83j5iqkPEzbAn0EnC2djYskX/NCc2gjPcriOzxOQPjzu5U92kQcs1cq
TH4fRrsdl3Xn1NESvTmpnuVm6TUAPpRwtUL21rmM+m2iivFGyRcMjcnwl7X/OONF
DE6935yWa1rtkwAnxVA9mioOZzzCg1QNr4gqP1B3Te5U5gOUmIWh2VUxgyzxzwI2
BDkZTebkj11NV+wf/XBAZqn0KAvxMPLk5WCmTHAmlr31ARg85bZ7niQ7WSA1izzJ
7g34dfd4EMWOc+8LB9t8bEa1qAFx3EvVDz3jYeCCgmiBzJo7EyLN2rGRN07rh8mi
jTmNICSGSlqhfVKjSjM+Og2bQr4kyJNpz12ouoGtZdHzNtHZjuWwJ2TyelE1aJ2A
/e3tXEAANL3nbfIr7QO8l+c4eqmbiTWDqEStCZnj1Dp2hZtgqNT+sFQkbdIblHkd
BUAxsFmHlPqEOSJ1f2RT8W+vAAzuPsEkXTLpNN780sYzbkNttvP6sy9H5Wr6PqFx
q5nQWB+ZXFgWw5DaTtaurva71hfawtDOVkKds0pIn5gl0PB6Ef57nbZEiB42eUL9
qIhKF8FcZ8Ym6xhMyBc6wf1w/5Zym53cKyuZMfAZd4nESyohcvuDZUPDjje13Y7S
w0pnz8JK0SRdFx9pGaiz/RvpRPSM1Vbca2Y9WxJ/3mnHw4mbHAUvXtzGlFJURIex
961NJpoxcNDsopR4gnrXmM7SK0hIJOtigLNEjxKJ1gmUNHuVQEPuiT3jguVRSWS4
F6+c6EZjSrkj0cl/8PMWY3A3J64GiFQLDnt0BgK9IeJIUogM06Y3lxajTk3cAnen
zNeX4/6Z6NBAeaDL6NlaQmuu8S11Q9dVBblHbvmVNdF9EluOuVwq2NcY+7v1YDK9
e1FqKvaYFTvnZ0QvZJ9pB9xIX19isw01k6Z7JTYhd3+bFBC4DMf6t++J9I5zfTI9
JA43URy2Zu3iWmK9U4vWZlM+UxWWmnm1kgPU6V5FNfn0wQpie7lZMdqTV/EbfTc2
RkG5NB5ajLMSR+e0lvgXetT6K/gWBDnGX4FTV+emgh2yfxUHDynhxvdGa5rjAoeW
kKs9hSiymt4PuJRQkkwGbBNe8WsBe8MZHxWYpDtZDrTPcm8Ysh0qmCk95cLUqyvj
eNCHvmS8F2EHzzrCJgIpUl8hb1DQBvAD0T6WXaS8AAE7ynGbq+VZ+oStl3osjjAV
RdGSYFJ6j7qaTVvj6a+EGtAt/tVfCaJN+4RAJScV/OMyKsiNFMsbrg8h04eFQI5r
WOdvc9F361IM8GBj6Ccvk1CpdFkmF8eoK/vJnH4KTFsYaObN6HcSATbaSd5vEaHN
sRjbrehSTKvMJJLKUJd7nQ+oJ02UG09fQFTIIDEWn6t60juO0nuf9UhJ8u8CdTNc
5iGNAR02MpX7+5L6HXchjlzZGzlzjF5ZBgIFzUiRw1Z9iXDzm8E1BgnnZ/KfoJve
lueE8TUBAj4lvV7tBXQZ2xEOwV7kClZ5F645Ytu/Y3Rk9fERWeEiSZUNHbuqsjtF
Yxdim9QhSofJF1BFL3tqbjZhk0LlmtNf40CzdXLfPuzXDTNGZHwt0NyiUWJW9gBw
69n6P3kG4aHLjRotb+y/J8kl/gca0ivVXDMrodDpjTv5+35F9uUXXNHfc9+q0UhY
yN1FxduD/HZ3nsrcbJBYXjbrLWQ3KRq9TjHWsfssaahwfzUdDdAgOGQyrtEfHK04
0ksLuuXRgt4z5jsV/Wk6WAZiJwLaMIZDRt4JB0Rau1k5xVCdQO1/VCamJJEJ1t7C
Jk+etoyIbQ0BS+IoW2XFy6T+xCuxiG34DFwOagA/cK43vVszyvsdwuUMJJRsjUFd
fpP+mzhMONb0Z+OY24QRZD+Nmm7u2gBULUfyE9g317cPykFixjUjj3kFq9DccUyj
dsyWoY67NTg6DORpaiXlK7NAlwn7NZKQUpu1qd0Tzxx7q8gu6hXalCZHzQRvz24t
T/E363OUP1Ax0WcOHSajuMhTY5keX5rSdt/wq3KP5qHTjYPpdiIgfuOZGpu6BtMz
zHtX+9DAMMvBmEBY05zI8P9YBgs1yUi6km7AUEPcCWxmmeNHCsZ1z0IV+YWsdscr
Fu97WWWKqCKSVC/++aWrYy93EP+tbrrx/RLeoNoI91Z4bp6nmhOufRETM61fVQu6
zom56LlW8E93ohBQVoRIcFjYL505w7aEY9W7LOKoJ5WmDZMkcQYnUQBLNF0f0v9g
cd71zd29wN8ZVzzWI0IJql3I2bADqU4oxkfz7pbDFUF803tiQtFsk0RMzM6LEohz
Eo0tU4IjfEjjZea6dh37phIIzJfQQnpKON0O27XE2dNUxsJSY1ZIbLpTiIxsgwpq
1LjtAbaM0lM1CHbkr584j+DLFMRTmPZaJhEd6Y3QACU2tqDZGXPwYSkaODIpwzy2
g4wZ2EbfnhfY7qg8aDGTIc9lBVmDsNJ5Tj+1taNQmP9thNVat0Y3f9A3b1b3K51u
R9pf/zkguAw08ikwdbHQooqb+G3as+PqRheFQialqRogNQ6Ckdi2+/0oZFb7dFL7
6PlIYVemUdcYuYLJwSA64omxIIY/jJjkqjBLNIW5FU29VDQf6tKgQOt5jeIkUbBE
iwqFSQNCB5lec28Dj7MwoohxTWTQmoLXBqQnxy2oIepN2BPFxYj3lXKf7g+6D0Is
TH07zOhbzp3o8Jj59vg/OENWDv4pwOtsu+UBFVnlYmyl6eXPTsvVQugDBprLerpq
HhI1kTNghG++g036gVfY5OXmpoapYTbsv0gUoffJ0vy5VzhVwnXca3OCPvUY3lY5
B4OOiy+Xq6+yz/whsXP0LeiW7ru46ABqYMV9kBGKL3r6NMZYYkwNF+VSQOcl5S1u
T7uP1WW5kTlV+5c/MXEhp4kVgJ+XP/L2HOFjVJmWVgfXiQm5LCtJIgkyKEAga6Fl
6g2ecF7eKqNRQ5o1mm7cKRRkMnbuvfcajjVIG+WNwtI84Hb5VYpj2f1oyGhD+vYe
q7xcDjJ89Rp5Uw4EV6WhGZW0sQwbilAQqfAsug7cxl/r6v/DOi51Wf4Cr57z/GxZ
XamAluWGGZKp7r3s5sBn2u6zlqD3aXdYOixlSO9e2oMZM09Twj/2OVXcjTrZ34BD
IX2qqsZWleE9pq1cuuZ16I29i69z1qegXcAG1CBHY2Pw1c8q42N4VgOpHNM9hgdp
zlKNeJ3Gq7OTvmGw6TWIFI/GgRDHW6o2qsKw+njS/jTiviSyKfJMpVlGDM6QSjjW
Hy+ARF+nbHJlb8TBQkD/OJFiDNYKadYeSD3X3ErD6CB4z+gqTCse8vkSoBi6Azkl
cSVeE7UYFC+hGUNTwz9Dn7r9SuMUXjmnK0TZWBRaY988fsgqKaMVHgbPyFumF0JX
RUbiyckB7eOPNrrKZ3jGBDUmfaRdjEoozUFf7oKrf+4LIqUS3orSxgQpz+EiIXLX
shiKJbLcWXxt8FB/4yKGxaEkAUXf4RN/XsrTzfv3dI8uTCpI8Z6IeCSfv2EEqeQH
bNrVkHrMg+L1RnJFga9GfJUjIZXmQOHxvm/ZWoWPExwto7Qtbl8DwxrIFoF75qJv
SRDSu7iJCi42Tby+pFwC3ou9Wz5xezoW5D21SQfq2SupLNo84lqJJ+3XQuEa/CjB
2tJn2s9O6gdRZbnJjfpn6D2PIp72rg+R5qwwJe4jc46U9hsW2WoM8ybHSX0FjvQP
86ZuLjAW+OBaZXP+HySUvM+mosVeDvfUsabt/OI4VVOdPFCcXiNMng5J48nRRjiw
QTEGmiqDSGpYhstNxuq0NweAvlW8A16YIEq10TU9Jy7nlWJoeAAxJdWWpoXiACvx
1YIh/IBSK1vvlbbCHMMcJudRfyDiqm9OoGW+XFuE5JRIIwZvVva4WE9EyN8545Af
V+W+jgHO67buLA4vhdrxSLapBt8Db0NXLSCy5DaPVpx4/yzdHc5nyS4yrc3oJb0A
3whVfOaAdNTlHfZUb5Me0kj2qQs14ibvDQWH7+A/o1S03Xj0jbh8Z9EvJfHCvKmu
oiAo5fKiamZpMv+MwLUwgxNZFHkRQWxjOuD9qpcxjJICNVU40jz5rx6FAXHlEutq
cJIn0UUTY8F0+m/suY6tEIoCI49efAqIflbhB+yVZ7xFAmgJMOKHobrv6bYlp/Op
7WhehFbQmNX2LCbN50cHPXBhx8Gabr5tV45zDdZSruzj1iumdav1Cwrv3P5IbQ1p
LDxVl36MpfUrrEpuRaQ/vMCYvLF/kZD4ZRscbcKFSwbfdtbe/8F0VwyUpgpjXo/j
azkkwNx1H3H2wAEYrzQZjAbe9Cbcr1TkNjlqIsIgdMkU038GvaGJSyCUtfDmzoxZ
QuzA69d050OGOTRha5MMtKexJHy3kcp8RmvvQhmKvaUCo5AHTItJ+ferehNMPGTs
l73Wjh42JovqYrMaEszr1LoJ4qYVDkKi+jd/SGaxbDZ07uCQNZZAQCOzrHvXE5FP
UH6NX/r/m2Kz/4CxW3ORS1Sz7bIdjRlDtPG28CqZgu/Fh5clBSV7S1lTUY/x9RmS
kyoIUy/V1+60SouKN/lR5nQyLfO72R/KNGC+49lqSkvhxZsW9zfaqzs1lZZRp/Pn
Xlw5/oeGKiU8uSf2hgzuvUzEoLe6MrEqyhIMmshGojEAoMVHBZDR8qsEniiXBOei
vIYkh9Btem7NRTSbq7J/3Rpqk3yJArDdYTPLKeDZtbIExTSHfOiiIXROYP5fi4Ej
JXbPy0PRWOvNBxgsKE6CiQ/ae1tK+3xANsEF6cgKnrYMoyNdcegUUy/BFxra6a1r
A3wA1djPSXjnzCVHsNois4YCTLps7oIi+4ZlfhZ9nrNqyjudwMsfPkY7+vPCqkVF
bUgEcuUe3wp5nm19LfZDXiu/SXnJi/QskDjPTfAI5gvVURa10pbjs7NI+xYkr2Rs
onUX0ndgVXWukzy6knc069Jny+Q64tpgAofddIr9S+nycMSUUALKkq6Vgm3JOcIM
LTqe8mS5gXklMGqWEaxV5xRN4ROr99zGp7oUJToV5PE0sLnKTfOlw6bZTxjuGsO4
um7pLxus6+9OjrH6eJnr3t8AAmBfhkhestGWJmP9dej4W8Npwmrs9FR768+rfYDa
SfOvEJON4NtGk+1BaoxcwxX9K8n5wk38LNTJv3myOeVDf+ESafUuMMltVGh5nBcb
cvu2O8efJy9yXf2qaKXUw3p2tdC4m+NDN+hK+nL6wuA5MoxBBQ+QarcjfwChriiz
eJ6D1O+GVNUOSswbdJO/YqaT9buVVnEVxxpEwVqXg9EMmBiVnTKwisZDynX65ybv
/DfhrpgL5zQQH4UCXlXMYKSgzYBq9wtZXGt154ZY/jv9L68gFIa6/JN/5ccONXR+
5xgEVW+8JSf6NKGH4j0amnfC2cPfb1ZzW2KvwGeL54rFJ2RlfEZTPWN4bhVNcUwH
R9jQDeiveLWXdk/K3Hk1jGdX2bB3U4hfB7rBf6BHpU9oySs7IAzli61rukpsQ87Y
sjmf5jtfEH4dtxOqcg3G6BB/3WC86VZ71L7VDkAj5vuzKA3SQ6+9j60KxDX/zDLn
Q0TtvV2N/7w+DZQZPiNm056Vpog3RVJzGy+SdJzLQlryWPP8Tnnpal9tvTtmR70a
C5d6dpXMg0wtrI2le8bC1nJQTwYrsI0RmcoC9jnNCntjvnPn0OSh5ofY9VqYCjPd
PPyXHSttGZEk7GS0JivmWqri9jT+LTv8a1wj0YCNUMnyz12eUJ1hf9h2pOdpKqKv
1jNPrg4Qob/G7Daw1h/AS4URX3eqw1fmyotidPjvLpuWFOYfhNvD5Jw9a27T1fHI
UXMXhJBrtw11jWw7wc/scgqB9YoP4XtNIIyQ1pBYtYIQc95ONSusyOaSjytX+SIU
MZ/ZhCsu3OkqiBgt/X2SLOViATL2UXwSAm8vU/ZJMRZaj0u7vjTQKJOgp4USeHhg
ezn7deoz5c44ZaQ9dpTt8Y2JLReNIJhe4afUikZjcDmwQH6AMKUK2q7uADVdPXch
RPSpuT6gPM44Qimsd97hg+RtjiGZPxJbJc27EyvQOKaZqlEQXGHo3Tpj2HaVTpMZ
8Ms1GXWg0LkiElyVntJQc6+RvmtA4TjQWhOgJxBJtktyC7FI/4+DsobUx6bV+D6s
/q6LEuxgrEUdBpml8Yb0sD2omgWdXEPJZzhKwFFzf9eY8krp18YdrDSilpElEGL+
T+J/6UzVPN3dQd8mo1DwFJZt7RSWtpBMpeB8NnZLFRaeiPGbkEx2m/ZStMgY/sJX
tVWkdtVUI938PVPbnImkiH6OAtlwqGyULlnkY6rNJR3A8qDUNLbEVNecrTBKGs0r
bbyeJye9Z6VYXPO25sg36K+AjNdRQmOScmzFP/mc/voqX23PyvAVf01oV6tZEZ/t
RWTzo7wXTRb+DMsibxnqBxxpvUo204Djw50EvgHYTvv8m7H0VQpyOTEQf8cG/WDS
DD7dyF5ZvlHkS4uSTjSq66QOAK8zBCvLKO25xB48Ylp8W28rr2ShCsE6r9krpYx7
g27yQIz2UZuBuo9wDS/CVpvvgiEpQn4BOwU/M3nh1DqVU3EZclF4RCPaF4Ez8fSl
W4kogx/BDDQUHee/M/R7t21nDBA78ePzDSY04kjC/j6ofHaixWL9SvOLDG5G5K4S
YHElFawaB6cjaRKAQ00cM7lzjVv+wMO/HIxioRfT3/dVmYEKOETJKQcK2nC42AUF
YThJbQSzeM7nNf8M+uYPyyaDcLmN4GP81pK0IkiPDMLbYVU5rL8IvNixPcH9ETKw
TfF3TMII91pmKvsFSyufc2uQeO5Shc0UEWkJwormF3pKQ+fQpz3NUKaA5QQspffW
HEseonJfCny24Z/d0qz3Ymo456pvj8oj9Q9aPOO0YAokRDdYkuelRFY1bLdLUFOG
XUqXjnS3K6pHmNOndvI97JMHEhMKLt4jMV+d7277LTF/2L/XSthhpjUp2dLACo9/
E3/CtkPA76bcM1gt1OJtCWBo3BqhHkEoJrfrBK7bOFikO1aV1vdT9dusLPUWzgM7
E5eSF2fd/sOQpyBZFpNAbXlxVdI/hR/yvoHZUF9/gJ2kODQSiok+PyEYmNeUKjlK
nqZn0oxTFOWSTZgQPrFB4Ux75ozlz6GHJE2p57/8soqkkts/YDMHQNbUZW0/Lj1r
eqpFsvq7qfzp7320s77vj9BwxaWVo7x4gk+QtjUs2QObE/LrNDGPcohSeDwH8LF3
y1a1QLO1UX7PGct/T4wtGPmLvtgmytNpunuZQeKsgeQE3DiG1wBcfi59l8HkfxSM
x5YaODfc2hpRr5GDuMvJeGEK765lFtBwlA57zgPTR5LXcjQS5DOBnekuCVm+snkL
fvHLm49cMHpd2pZprRS7dilHpO0TzXVrqV+7HXPTYuO/2iQ2nKiBOJdY5+Y/BykV
Luh0D+mLI1R7AkcDzarao2i5hJG3wzKlIa1YxJVWM8xB1mWHHxppuPxjep0ZZkzO
mw4xyz6l77zwxrUtdza9c960lTu6jrFjv6bCRo4BuzpFVaDYoDRZBSft00be1GjX
SDlwtLF9pc+3f/OA+ekY9PnoVDe2nz3nNCQEOTXE5gZrZwGwW6VxHkwuUNBC6LPm
2iYBqpQISuG2riWuSNjmiPmDUGJBxAF0hKd2rH+R597SBGc0WZHuFw9xsgnrozY5
DtkZ9IUg0LSB/AAYyFYh0HFeFhiKXQgrA2lBAZrt3ALoDqxasg0nEpIoRuNOD780
ib00JkiVU8LvNo9cJE4J/PB9JZ64QWjUq0wKDcTBSe5W9gT84TAiW6DDDii077aR
lhEYk6FJZnfOReO3+hYs4vRmcldf9WPRdx/Rr7FrUgv+fN0hAYoYaAC/u+8aNsMY
iB/xd7dYqlT7cfTOWuknoHYDWTqK4WKs7XVvJ//vArv9az6dGc/7u+QKjOtpPhct
sx4m0vLQsf8OK2DHuqITzC07DE+5U2iRx1xcdMlBxLjN/F+NpjfVvw0rOuPcqvoR
qFIE0l2rsecBga/4oAhHm2+mpeSWAsNXtyOV32q6e0o14oHVv7LYLqPcKQZD50ET
59eDEO4OSdVrR84kgMhedhNePlyI4vx+3jYJg224JongUEh7fJKG2ku1gIRCcDFT
vytzOaENK4g2BjDR4cpm/Pd8yOPoks+Pt65DooCieRGqAKWE873TbjkuaZut+VHD
24WN1NetQW/zzLvN5fedk7FieSoEVdf5Yk5gRPeyhvZIoEtXBKKMTJ6d9U19EyoQ
bum67H10d0/H/uybaRPq4R90RxEAcKfvNqY3mNM0Mj2FJ3XKR2KZZN1Db1D07arp
w/TXU48WlxAPRIgqI709k7pZEpmk/4pFn4Cei0D5XeJ1r3E9MJ0tcpvY9czQdx9a
8u4WV2GCjJ9m2kXXX8OrNMCXMiXkQotSHUWjQ76cx6mZtxbUQWYPH2pWYQ3IYSEp
cFqjkFOX+iDSr3b2uMwVjG1a3iw8HslC1SgP8zigzHFRAHhg0CUq2hYajWswKKEW
SBhNXUiILy5AX+Bs4DrUrgeLYJL9sBMBxJld2CcRYKc391e+dzh+dvfUlx5IlWFk
qwl1u1EXdV6WNaFn7ivXGY+gVxX1KBOYcyfkrj+Z5/vVcn0PAkkKPM1s/pGdgJYq
1rEP1K5ri0HCkL9TcVu0ouMIxhZ3T9DHhjyGD/A7q42yXrm1fUGtikDY3MSlLeRs
qozTIzAh5u6Z4Fwo0/A3eGNAwMm2adpw7k00dlwi15RWpT2mz5rG4mJ9lQOmWoSA
05+xjXoYCM2gpcchuhfHok8v/Hj4kOz0/nfkc+9awkY6Y5V0LaoiNpeOgemP17pl
rOP0Goqo+ryeAL1Q+a/MGYYw0ZF+3UKd0pLvl5zitVdj0zo1Md3PlMRgsJ2nLOvU
zTTyze8kZE1IsLfLfItgdd6yinLIHIH+GhEgdq8IU7eWgosfgcIV2OgugIno39GJ
b0y/V4X1wfxiKZ1E2YSqdW4lF1R8P0sF7FPwqbb0NZ/fGqcigvbPyeeHoh3tiM9m
uFN3BhtPahmXhqP0mzzCqcDz+M7k74roJcigUBfrAcvL3X7lmxuBBQVwnakmAh3a
+WQsfHaipd61x9FJ6zoyiLBGtjKnlNKdaOzF8OLdE0JQFbbwxvUMlQCmfKsCb3bT
b/qYRewgLchfv5NKAbCg1GYQDCMhgXbtzEHXeisGWTXRvInm9ui72LzwXx1dDGNB
XmWM6bSw5S6/QuiyQmV2XXtYTyRwV/1SXGu1JuXyCZ7x0B7Y/Jz2pqt2VCvVdIb/
W2WBQI3bKunsmXlHe2USVvjJO2fKvKfsWQuQHL8yYebDaHxWNGZN2TZOeh6wIVxk
hSRfeldrx8QpfiGDEI2Sz7bTNTZTjcLGWh56MELjTCMxzO4zipAkCO9oiZPX/C9q
XF0uPHPvsuWwtqQbZnbn9zOus13FfQ4TizDj4YhpIYkUOscLUK+r02Z0xYUDy3Av
WZXj1ANCJLU+9b9/dpF+s/5XQVH5rc2VwekjM3iiYPwkKkdb+3vuWHz80mbQYyaS
3NivBzCHIcqJh7cw2amoYKUb2xNwmJqAKG/cmf93etGMlL4yavhuMWFEPSEnNQMw
F3lxOOHYzDvAlqqEI5FAvphHRkT6qghrRvrO/V0iiHooITF0GYVkc6PQUHxtVzUB
wIINAgMjRqNstJ+5mei+FGlqWv/tMaODSBEzS9R7/eyQXzcpcqNqZblD97Q0U/b4
yi+OJwL4pCwWfPja1uTVR/i1Rvy0FIasJXMXIu05mNEcGIamAPAuMrOm98VYJW44
Qd7PheSrI/RF7uXNKoDIb9gPgbMWNlYDTW9DSTiF0ZLhT88Ns72QZmXP8i2kdkoS
b7zw712RLjne6rzVkZLOCzuM2WTY6lY66ML6LZIsHM1gZq2BHRGY+z1DKkUQ3DD3
cgl5WdwkE0h73xwTOGPKdgF2WwrWoAJu3a+nqHYNZsJZwbyMgpzXyQ3Cw9mvTFuk
tDQwdq8/IqW2ZCahZ81s1KAvS+abZyvINuL4pqXj63Q0BlDpc4zudvzrekiHY8y4
LgI7iVyjtTN+eOrhgdzo0Q8jyw5FK0s0iq8PTU3rQgIbAlQeESls1mo0ZXVWCtPZ
dBnt8aZ9uxpgp1LA54wZT48hFOSuo5FG/dar+prElds406E5R9cHFM1pBl0bpVlY
vIsSDCaqblgxMd1CZisYjfCbxUOJziduZYFJRW3WQNkQoiKDNAv1twhkfm3X6uVj
VG2HUYtnJ725VICexeh0rD0KR/SQVpqii+2PEVnaudHvTZ1TAYUOrZZg9tWRncrE
6u9a85KslBhmHIdA9pRM30RMGLeCimHlMZBw9kdhjoLg+xMeq5gl25FpMiqZBv4B
FyE/neaL1EwgHwMk/bMa5Ygc0DuwCI2MflvOMTC3r6ZlbIbeBboYIO24ffRvqGyX
UTKYXmlBG1OjSf321vkSxlzcJPqoaLVQ/fi0rqC7XFmyzdrFEhUHXRDFn3xK7SRx
HDQZXIMWBQUBWNyemLZ4fvSWqIJBT347+tSfYT2ba0o1uoY4YHMZwzFTxUSvNJpw
xR5lAQugExVEJktC7X6CsgZbakxU7V5bHG1lDwJsGo8abxrAqlc7c/coOFPBohRr
39Xqw1NzR8B2Iew7Ojc/NsufxrJ2Q5Ot7/IdiTgYtWZv58Lc4H2RsXcEnMlQYHQP
/5zIOnCFZueII4FwPNXMoGy96dW0JdtlXfJpPeIxNCoh3e+JhVYJxzdmYZxR9+Ib
0quzrX1a/+f9/jgqgbC0JOEEOOr2J6tyKdBcpGMoLXs5wnRa4nl/qB/30NqXJTPx
WiMJzcJG9MQ56o0qerixf1BZzSCBrecDDb9oJmROcZLkHVZN0uVIDaZQ1c4jQ2di
QWZPHDlwKfZx296GeFjQrflTa+ySh6DyPU0g0j16pYFbgxc1jMjZXioUlM5Hzm/4
Ax46BuNaB0kMA4vRS4M5kkL3DoamCjn+DQSWOHkI9GIZQnoOYCY+BXePUd2dV5gC
Jc2YmVA4QTra8l5ldiyGNAqpNyezKdPzu1ZIEhPXwWav4RDEQ55vCVKqrlTledhC
FFB7I1KIvyayCyextXdzhq+hp0zh5YHB4/oLNw4AKHZh1J/oLaJ3DEqtrOR8CotX
/zsQx8jzYLAcgfkQknJWZo23qCgYOVy8N6a43iGaJOhWqjToxC8NWY8cB+kkuFKG
ASBiV/t4z1qkoSjgTj+63M3f0mClwpFUXFnyo1ucvGmnoDqihI5Cw6QSM+MpqE+q
4mn4rkJIwp7E7A/jlsDx1h+stdmRcisZzOix9ZssbMMyNYqYp6FO6Zb80ma06/L0
DKpPidrp3xjfavrL2ysqdFdvCRNNRVsfw6/jb1hOHY+xNtvD72z0gKBIYT3nrbAN
YgG8FW4Z4MVM4K+gg7X0qJFSNtX98ub9NEyGR9wt9KLbaWsJEh7TMrr3n9TmcLiK
6wAGA4qV152ujRnKVSbSyGcAWBeC/FFlMWkv9CQ9afEXAWDcYHa3ullfFEIZSZDO
/s1X4VZGeDr93ECmNSre0GERbhg6QVDSqtoXD3CKaiN8d5bKBKOK5J8jCGDMxo6Y
8s6ajchnZSaGiPatY/Nqfsy0DH0h7RpMLdrhK0KLDFl0e1/SAAa75dofytzH/fku
uvnWFiVyr5OP7/f58283u72QLwvqreHaueelc/+6Eun16Qu5lmzyQmn1azC7wLMT
E90z8YMwNykOTYmTcCjycLn4vG3MfPjbncb3AdCmWg5fnTppm72TeR6lN3v6KPZd
v+e/lWLmgoHMBMf/cb0mHZ1qkHOMLKXt1W8WsONAjKsBPuN8YHzWLAZpmTH+PMsV
SWO0L0GNIyxc5BcB57+K6r3Re/Md7BjDiJ29Je0th/E0sIoobWwyq1Z4Q5iHZ3qb
Z8PahLJkICxsMBaNLoSjdIR4cBmGW2zi3fPMJeIMOvjPa7f6xsI/LjwBPTFeZ8/w
JY4gpmKU+2/N7ieikpX851ic2sdm6/SP1oFvLjvqqXUUo71m8B9TAtF/B9VWksqI
4oW3s1y7RUF+NCE+dz8f9Mez4wnRJGzaxhmKhKgoRAjWI4RNzSeColXkz4I0ffau
W6Wh4ViSFeWSsvgpybhJ6QypJLkPUpv4h2HfvboapLOwa269T8OWr26bCzTrlXPr
At+1ublqzOwh0L/89WplUQzlp7a4d7IH9ueqtlH35Ig0yEZ0x9g+w5mTtrbabv8u
zT7FDxH94MVin0Kb8ke7uPd4rLLZ2DORw0DoLvYKXCKIxmuIsSqI+bxfeO0eV0ql
cCbdOUl7+Jq/dLHKoQ1IYFP+lNMb4XMrABiTZ1vtRny6Ci8ROSqcMwh4V2ZVWfGt
2R4XyE52G7I4YqxsnXwRl7WJAlQAnhBcIxTWrDkxynoz4H/FMJ5P+FNhAPD5tP27
Im/lZRO3CcrxFcBN/vcEQ+zpDyeUpcqbZpIVeqIsTQrJJOgyUwRMOzpWlqDppnwv
Nzk7I5tdTVuo8Ha7aUM9/K7ztuoP/QHoOfJiuLMqLh+0K0LRXFMAS88glGQaUOP+
dnaiF9Ob0vLgnZwHB4Y2OlZ3zkYzRvhb8Ebt9EOQEKIkE8uUYzfARHTypRUNdOfz
AtR7xsasMp41WjdhonqCeAWvSxRb4OOiPcm2p8HAqr+wu0EJqCGRz2Vsl+g5X+CK
7I9AO2+/X+k30L1Ekza7wVQTISsOeXbfkqnEQHkNpe2oqmSFARi7sUmw/TXEAIu3
e/oPfQXT3wAAgBzvv5yIzBfWPNTyQAWl7HvNnWRUv2h0edRj/qZbt9bumPYcVWQ8
IHjB2cNcLaStwdQSL1RY+vkwYP+PdM+gbhzudV4JRX66wrt9CkMbPBKhS46Sz/C9
P3lrqSZ4oVOoFw2DC285YiBlfVUSyuLaclDPt5eHRUWd2eyz9DBIWTnUxHqSvcoS
36kIKEnMcjqW/W5J6bInu4MMTPgmDbkj9yJMqW3+07ffUsZWYhNWpUoS7OfpiD76
v5ds+zXpQ1r04tUG+eqR2ax1sQ1x8uz0HsQY+J2D3ArGuhfpWoIz4y5E7xtRpYTL
5xRoB0YB1w+pj3dsvgKA2pVomD35asigiShoaFJ1MhImGbEi93WY5HcxlZKBHXAR
Jjc/yspKe1DicEkE8c8yl/hTaU5rm0sylZHm4MrIkWLl/NvXCHG3kdd4vem6/oCT
TS7o55D0hxysAK+oUz8TZpoLm8aI6tVL/mWGj0qOvEfddMhZW7UUbLFnM9UYmZBr
1gBe111j6CQB2kNxKX/t9YYErtfrr7L5JABqqTT4goO0JITVmG1JKHOPvC0Jnb5U
heBwtrx4AjoryzyAwCMnKQmqIsb8p9aAgLmWvnH52QEsdF9lBcdtVAj+uxXNEisd
iNHGFVOIMdi6CcJWgu3XWBRq9EO/lQ2unwcua2b/qgfifnESwxTmwDpeOnSKASPB
c3he/mTxOqP/CUlZKPPbBRoj9xcHnX7fVvwbZCwqdpkJumfK39KfetdTJrB+I/rC
dndpSaMsrPJ45wLGutJAfeJxyW1AuIlk13rXtdm+8qEVBLk6+FQN3YCNKsuNGIAZ
LzzcjVLt5j8gq3/HT5jbe//nj4n9nLbpMalSckoAJqfUyhn128o9VIFP0CskLm3C
zCpRDrpR5Dcr9U29F2p09rlZsfVWbyZmgFRBzGSM2BJ5urcpUCV1jVBS9HWEyjrJ
+rK1Ngcnu7h4gjt6fyMf9BUhF3mULF+b5mtFFE/Jd+syTJFElIPctuxv7AZW61ja
Zl0r32NrTNFGYNIUO8sazZOaOcgmpHp0tXNQQXWU7dmVHesTSDwbgNHyQAoPAYwA
HSV8q9QBNIQOabHq1TYhMxTiLRK3jhKuAQlu2gZqm/IsMsvL2EDPts4ggDuUctko
8aEVrmdmKzGvN6nZ2P3mCcFqwHnIjoYcVMO/axQys0RscwJG2Dkh0GyYWUCBtDMg
2UVSt2l60zVNHlJceJPfp667IQJNlnkiPlC3nt/GeTr5OEoAY468NpukCVt3WWBy
qjdTLyDc9ZQEE91KaMoUfCEmw+Ym8aa1K9URGzZDTPOTBvzq2OuYQo3yMvV8N/2D
g2EEsw+grA+eF3OUJ3FR6Nyw/ykKg0D8eNOZRAq6eElw3IfKF+ulGS07VZvSD0JZ
AgEZhFCeLjHzwmMKl06heaNTjnbNEOop0XgX+w/J01sQRzE9WleoMxKu6jy/hWJV
QZlyXavxGrL974IbX8YCtMCsiZ6encO+5R44HMPT0IXuxTz1oB8cnOWEC0BTHTmO
n/K8+BtfQd+N9pPBBQcagdjwg+WlwHFlg8f/XylRmMNlfCsal1IWqf7NeG3PlMgw
zyupMRBXiuXI5tEQqAonEK56XELYdllspexh4EBZglmvk/0r0k819bAMgGZWTCQe
IfhXjW14HEIgH4sy7RgtSKflgA1DE05jzW2sOScmaVufujyvG2/cOBt9R08obrXr
4L8qLDGanVExC1wt6e6ib5OfiTppea8HtAySRedzuSrA0l4G+EXJtTm5wsBtxHTm
F1FlSAei4GOS+ZO5iVF9fsIAYuGEPwA7DoL2dVFhejula+u8/sy4BfLlpwTonGxP
KhXpkLu7C9dqW81pb8MI9QqRvsrsuvaddh8AHT39yK5cZx4Rp8z1DgPeXSWKOegJ
f3paPYa4vqoyu1r4zg1OYDF+tirZkTOowoxnE3qYk+62XlWGJyiEZpTtw51xD3hU
xVtAcsdLHR2FFvio9Zg+4YfP3p6AW4ibjhzErWUBVnbjSl2Sda+ZdZJaqWxObbfZ
0DICcarlL6+AC3px9JAndVdAaW4C2LugG4M7EmSaRzPs+2k/fd19/0Ywf4m+cpbg
/eDqJQe2qJ+ZltiCMNoLGGGuF2wIB1wUxeW8BlBjtrqlUuo9whzM7wvG1pi8bZ/w
6TxXnqlnKEXntm5YWfyGGfrtfKcoFd4Kq6W/+drgxdpnaCeKqPqojfgsQ1+ghABh
KIMoSgRzlvlSgePq+rxoJaokrFbiZR3OOibb0Rx4OTi/BL0cAQXStGR0FWbo7LHv
67NLqG7hvrjQkcA3ukvsIpZwY1a+WncOCGKcmSU1KmN737EjSyHe8SsBUqaE8Bi6
uW0vQ9qRU1u/MGnYz95K8QfU3tw6CDlS/vQ3opw9onmMXTeaDwC+yhy6owWAsNtP
AQRDNvqOn51Dmsv4M8EHMhvGgbUSRm6M5TKo6e+7bFXjdsHYwIoJBEj5qOaRahzx
H3MidHjvfhS7rQNTw/ngYYPWmYuGZnMlbproSwGkeXCaxyRYSEJdr7j6CNz66WRh
2DD0TR2OG+FVlgS58Xr2NVAi5JP4t1i8vRHCn8vYuSGRkveumcEGNMQC5UXNUYp1
EcE7rd5Osb2FzmiNHAisMafihLsYrhOveq5InMzVyCLOSaUnhCz1fO+vYEkUL2O4
WWHaSQa6k4mqQ2ZcwOmf68bY9hMurtdR9n94gpbyh7JGbwac/zC/57NiibsBH/ck
9dWJJ0IeFnkRjTjpfu4Dv6aYn+USSxnS4JvfTDZavue6Z4baenX+SB93rPDLzZ67
XQ3y2rDlWFt0wzshWt7MhujAZTWaEq6QMBP2HY5ktD19FgPfp8UUjlK2vAqqOxrd
BsTplEyRenm/LQZpJ1fWp2ODREy+eC1gtUZKdeFSIFdSr+dfp9rm/ySiC0sR7nfW
JJSZqI7CS63wdRnc9YMmXxTkGt1chbSbqKDDJZGksb4zQtJ75eUB20ICB7hOHnhe
IZJSufmHY/QfjsMQXLnHba2PbNVQnLLeuBl8iCTFziNArOA6tx6Sx7Dyk6/58g1Q
W31sEP3A+ot9sL0Krp4CPGEgKKZ8UZxn1riaX4NbCB2ZTuSdR0KW/oYZxR9bI+Kh
GrGOKr+Sds3GY4MpE8xmwx5seHcoMHtPNAIpurmL+TaT2y7wp2XwFjWw8Zdp1clA
JhUeDZ7eDX3SJzOKXbfzSSlOuR7Lp/fh3E5HDJf7N/vX2ZBk1+kfHF9D4bFiw3XN
JhSKbGtA+IyyTXTuKt6e1lovaMprH3nELdjQcsXHfIQnm+BckJ+OEfCkpnP6Uz2m
A/xT4yfrkFwCCqO2KXKSUYEALX2fk9CFhX5r/PDgCvEKgs7bJq0ZZm/Y8N8i8pyE
hSNyncBOJbRSkQ1zCoeQBkTypdHRxrZdk0ucskoZmXoBZKblqV7iCp1yTNnDYcZj
sDJNBt3F8W4UjYp1BQ9T0hH3Abq+udIWd6g2HM+Y2TyAHh/1MDUEyVO0bn/UkIOw
YqcjEKfbDyKuJwlahZiW+E10dr37M+wHFtH0shi+pTRdqXcGyXXxGNyc0dEHpyfm
6CnrBYVCQV1eV2xeUd66P5yb1ftab/4QAfLEce8E38FHyxUWuUdqkQ2RLNFGcZ4n
ysP7J6gPSTpGfdJghPawOlPZ0y4W1EKOsjtqPKK6DJvomXuIzkpOu8fAAEuOHZJ0
5X1U+YzplL13nzLDp5q6+sflFymUIpZXSA1otOTyR1dr8HRiYGojz3J/6qQVY0jO
kvUyF7seDUz+wjpuqwnNW4jMgy86OWliCyfHsSSS7/yAMVNzCVAorqve86l7WOlu
hrlqH+tfAiQKqQN6xTUe5riQEk22rdzANi9lMfHDCnEzcEbI060mIuXABTx1NRVV
gGoS2MXemBxhiHjurR4d/Kfdl+r8xXijHhjLqX378WfcL700MBaY5Cx6zMemsIRn
XSS3NVNnUYLyHubPEMnNMazNl8Hi3uu58SFTgwkafIFV/uIMlfwNnFngwEVYtqWd
xV3CRbPpuha7j58nMCD9JQbaX34MrL4MWGwZksJ9N5b6mABf8nHtuuu1J86qMEvr
lZlFc/nMiNA9PCueRPgaixe52oasjGFMcY8WUhIiCtb6RpFlL4xZjszsKBAvS51f
HCvOhEjFCSrFj97ZNS4IGBROGAEc78UE8GWJjDlfUDevI/MhtXxqxt/q7y4Wfjm8
RhGRzz1l6Na6D8CrKGKklk19ztNOyb5jxDsH5PN25u5cVXt8Aij+NTqCmP6IT3Zs
pvE+MNThXPDSO+itNUV8/q66QjyzRjncOzGs6UIIFsqZQjTQHcY47euW5aOy62MA
iOjI6XS2xVWUHKgjPDAqmacAGZi7AwLWpNYpNBbLwkt5kTdou64loU8Wpq4iUTCW
ovmVZdhO5vQyCpzDCG8balrRtQ9aY7kqjOaNf2SCaQlU2rJ7GPpW6eXa3N/AcKa/
OjfK3Bf87lBmPwAopcJECNwC5aGvp9sCxTJRPpAWbKOLVyujLepoOr2DICfvAwNs
AVlUdCEJrE8H2lwmig9Hf9SR5zruu9mXb6l3BhSgI/dwqxVfgSdAVgv6O5TBDVNd
uBaZF79yOzHd1oiwx6QdH4w2c0tST16avqYIv0g2z50KSsA17GmoMuQosVQAy2zt
bzP6o3UfqYXNQy8DmYZHfKZ57Ej/ctAOPIDXXp3+nxNAwQK95heVyN8BXInrrS7P
QRQxPNoPhE/C6dahAMmbqlzdoOV71Q+grjKQyVKyAcfAo88gf9+hm2JzqHvs3LAL
3gbQKOmDaNTglq02YOECJ5r+ki5D2SdZZefsQDKffUQiNLvCaxo50tcTG6sMOXyN
X8BZeWYv8rjdFHtDKesvkC3lxg/46n6pPadxvK7RuhWWn+7cp4GLoKRJq0zSyC5b
l4GocAqbquQiG3FXkGQcrJTjpOxi8tHhPk9eGXZPGVpD+Pp+d7ZxeRJapW5eHEI7
Yu7cY4+TIJdQFfLjgobcL+wNtkuyd/deh6ZZz0kMRR6u549ACNgwTGak/cTWp9N3
B/N4akE/8IrSdMfJjQ3qmo4TYF1AwO+BPJyj9US5WrlF2o6yzmQdReicWO8U758T
uQg9OQRnUqDWk9Buw2ncyRVM6US5mWdF4DQwQ47KlESqZerwI22CmIy43rU+aEt2
TjiLsIZQ+j+cFDkyPVFwhwab49yWYFRyn6r4xR+uXiBk0abmU0aUTOAntjBLv6cG
Mx2TlN+yydQA1danFEve0CiThoJa9eRYGbkXNqmKrfQFj5wnfWVAPiiFmA/VXVVs
72iykAGDmw11nEm5s0P8XxB6rbR5rF6NgBYBg7eg4wyTtYyUfFYHsd0kq+vE+y4N
25mZMPS+EEBdCUs4ASQkyr1Fev3osuuR4OCY49ZZk2WUQ3gM80tDxJQVcQONCX6+
uRHFId1cP6ELsGWHRadE2+GlYczUO0RsbujutgVfSaHPDLWLESuXRoAL0uHdmCez
hx1Nf+N+RY9qRUDwxRD5khHRoHTQlj8xsJAkMJVeH1IjuMLoMe+peawvBvFFp++1
G5kKpjTbwWFGaZ4guh1IjQcdpy7/O7IRZXWB2Iq3LpuEvR+/pCilyCQyTDXUoheF
XbGmj3hz0G2ue8wUHzlehgmAUIj/SWVVNCgu8PIIQjaf5LdyDgmvylsWn1CWa2N2
VmyivnNphdVE3qbwWOyUmwzmhuWm7hKui77eh5C/kQGcD1m33tDD5xMoqL8ckWwj
4Eayto74I+GL6aA76THfn0v8RMdY6m3sK0tRIZiMOsCzvuDRKWNmCawqE/kMNz6o
3uCXG24VYmdCkKgzSg2nBvlK6i1gGAOvoqLdc3K5sDAU1FwYQJAMtT5odQOqycZD
V2sTC4AsDAShp82hPf57YVcNW3EaS4xS7K3WVqlYliRQ9O6gODArUjJuEACpw8mJ
Jdrs/9SFY1Y7LJNOgOmTtXQm090icGV3B47fFCGHrv0goyZ/6EzuGk5D7kh95IiR
HmOQ7G/DFCiIDJghQOz+DtD6g8OpJMe+H8vt9gh+8Kni16BMtflYRzWUKdGfTx+8
FzNcXg3hAzO12Iht/40tS/J0dMiWBji9cyMZEmxDUHNtOH6zjn/EgThpYSF5wkQP
Zb2GKdLtyrn7TDf5GDLzTwitYMQpjtH7awoE8aTYQONtxPua6A2ILP1RSsCyN6wq
uO0fIawetSV4rSy7AYmzyN6sI4OoZCzQFNZnLscKIgqLh5aaUxrXTkhlfscjkvGs
aByWO8jM4k0cxh9wH8Kuw2rkJidMnVq4Bgs3SlfdNKeuTt3k3pfX90xK45nHpUO8
ARvRHL8Nsf/deQ9M3AuV5Z2k+ZvCYm76pxzqyBffX2CrJ9aP14PLcous6bNACMts
udTEI09xgzB4H7rm+GqSsL0VDz8Y3zDN24ngeT0siDoCC/Ql4N02KNdVT2xQd36u
/IMC7kFvMLxAz6eMF1wgWNqLG/lAgU3sYBwX2FulJKzJaxbnGI5P1XPBf9CFG8NE
8aYKDJ24XbSC93Ce9RPls8IGU1vf6nAXxnmchBRjEwZn3X19fgZUy3PpLWJ38NX/
MUYFZn/Hl/srkP/TlI4YnOJQqyA/JW6CVueId4bJJ0hv3HGm6TQmtDPk3HXpaoT5
U/FwEDl42EUDy4R/hHekB0oSqw5wlDXZDx8D3TfAx5VUSr4b8/7r0euUpC+lBPaN
dFL4Lftd+bxY2dDnQO0N6VP9bKdjvFcaWbG4f4ZS4/wYVcEnD2ZEWyWWN5v4zkzA
UpluZqry4cnfewux3xI7/m0bJXG2YbrH5BlOb0kCjrYyqTrmpTSOAcxGXBrYrsUx
pRrsI8XMHLTtAyZ4jQa6yyA5UGqIvQiMgwH25lvhpTbrKcXXBTIRj+UAXNQe1zhr
OUUrG/t7LsmIlLPZq3e9q8eOmJVoJSS5bE8ukL+xaAoRc1VVuUFkm0SLLtNhuEF/
eQV6XZTqMppbSAfRVF+0e8IvR7TTJ7P2nDHtCvWDEOXnxnDfG+dvcSYPYzR/Ok51
Q+pZiuQ7fKaCim7XEvV+eJ0KchEioCkbdQzS6nXS9MXEizTc/JOEINIW7ogS4iv3
41AsYTbAcpeTygeToA94Fli5NIDEmkFwcZ09VEuXJs+dMUib9ynaIp+nARVq98xk
m4XVVLgWGXat6MhM2OtYANWYUhh1vWh/WQCYOI7fvjsNMc0a+hubVtDIM5FGD15Y
EjtdDywoI2OMUUiXhskQNvezFILnjZ4aMjVchVD+NPCuy0XCPm0u9PoZ3maIsNtV
hT0g4hybA/hfpo6LESyJv9efvLtfkZOQXGKVIWYF7OAIznTp4EixPIdxfiwhYgkb
+3AkZbes111nXG0B7nHlw1F14J9zVGHdc9PhdEFBteg3RO84pEXOwtpjdjBu5bw+
d3Lt2gHT3sreaFfB0d1nr4H82N11irumNjMjNafYQ45sAWxXHguTFshAdvQFoHzk
3xyfydooHcDYy0643SzcbcEFe4FHl7iNpaIIsBArqsvxWduwNcRuWTkDRDRq1S+D
h0odfu7mwbcM67ASXT1kgED62L0RotX/Xx5NxlXjkQmrDyLxXLIrgIVMqc59dDN0
ZawvFXuRezDVtbReR3aJWoWL/dVte4qrXlL5n3vCd3X8o4xDrbz6M31mhluZmxJF
pcm/XKUKseUVMqV6iyL5/2BS30sq5HZosXGKPT+AqnnD/LI7uTT6QOqrsfG96KJe
QuNL6o5z3ZwAJvYViCxUNyzZNL81l60cnA/SkduMy0gm95BT6d0ryGL8HQGYh+Mg
ZeX3dfGoH3819hcqbFw0HYv9myy9mBdCWT4lvAZZV3toYKFsrdMrpRQZg0rNYU/b
RniRd2rJ0eFfjouaiTOZSbuCABu7RcwILUa6leD1hW2GCYVbXiVJPYVRRA3quuXE
g2kopG3FdZydQzcNTVM86uTZga+vWoD1zoF/Cz8iqJWcCuzt9ZWMCM3C0Yg3MTLF
EnuXuwfg/rPhf5DMq46RRySuMRZbscWagkkKuNPfvbYdgkp4THQSSrP5be36X4+B
8b1AUhR3CTXpKeMSyMSaVAP4Kxp1kicd7Xpm7MHz8ROf0P7THI6p8sgTayr0Tvsr
HcA2eIEICHPW/0XMZL0Bi1sKSkw51BCmVoIgGcZSFBc5vRsulb4Ixd9/KVlP3eGL
6xaVsfCg5mX1XikhNcjkwGdY4szuNjRUdpELcH2+s6vp5eku2gq+pmmvugfqqINF
SVkf5SKCpYO5LMPpsuXhs9xmzALY0ue/J+7HTq9yuWs0H9zi1MOp4qZZe1J1FXFu
aS20zvUVW3IkLrxTBCwrmzW1v4OPNGXZzun+d7qZ3oTKjeE48weNsfpvU6XJEl7m
/Q+01yIGHS1sUBXVqRKLEM/t7UlscEMPM+f0NgVg4t4C5Uz+eZInxJJj2vJRWXQj
swsfg6Wb32M9jG/N1k1kMKSnkLxqxXMU3soACcE01/rmJ3AzqFVTLc3xwchwOsLC
mTQ6irK6sf9/fDGJxtmjLlCgrjSeO5BOWfEYNZ454t6EROJZUhIQJBUIm0SdKIV3
d/w5X3bFpEEAW/+jU/w3w4sm+MmdsWer8tb1AuBjBCwPG5UGq5o72e9yJrcrCCdd
Ju0VLobWvgClhTxwYnGPsgNZYExsr6x7Qqj3W0ClLbGf8/dYcNAD3eQMgMhYOcXc
ZXkWsP9PAnLXI+7Y5I2y1G2UBLmPkSc0+dSLwF/IV5hsRjkdQhO2e4UAWeR38ld2
A8nbipphtBP+VU6w36XzJeZ6Z/h3T42gDtY1W2J/g/v92cXHVmn0GHD7w+EnRBIm
keosg14AK2qu3XGSWV64imL1FBwiZNnrt3ug+WRuDEwn9jxwT4rGl5vvzCtIaAxS
Y0ozpwYv27gCW5HopG08Xei9GUOuH3rJTJ++yRfOUEZkK5+AfxWfYkqF+jeOpktb
6MurWUdzDZPTEiDsv3E6WAps0mQrFt2Q22sbtR0X9uGJ+/ST52cf0Mn8oLj4ldvv
WKlBp1yEY1kfqSUFIJUVcwKR6wZZoeBM0jNcY1VnMQ1yanFwxXvqIDIGXUnOxw72
Q2yTRuwrVrkmEQLRy8RaSHHrmfQ1oIlVba6mx7/Xwqp6RHMwtqQ9iKs0yt3ByUUD
WdHl4Qtf++ueWBemv39HVbwP+IYPMWVkIGvUCeDR9eWBF/AZxTQxhoC5kHB8Kiqk
oRZizeZVdfrGMiJoXSCVy4Rz5Vydgn/2fvIeDpaKLFDFkqhyWrRZN4KlHzufe2YG
/xzNW4Tyoxl4zwJrhFK9Fz+dIQaRust8l3M/Y8q9TRIn4hvYiTh4G65M1h61FTxl
XoIv+YIUWG4q9Z6tm4DPBNAtQ9S8+DdCVvZ05aezDNLyRNVjx0GSUMae7xbRfaVU
X2FtVfuIIona+UWPeTMJ8Yhj6pimnQLmTgts+mr8AFb9C5cLwGp8BCn5wNlPURtN
QkgSQl21EppOCzkTMkyN2m7jR6cQFsWHj5+UjRDn1Jkh0UaECQC6pSSfcUAExjEI
WiSl1o09gvsBwUuDtmf2r7i3IDhFySA8STlqilSYRZ0dz2usQaPQF6VcskMD00qj
vzOGxjfNn4sSDwWCfuXyoHKmECOueFIaHry+SqC6Vxq6MjBqJSdV9iSM459SozZM
tqQjlm9YYK+K1EQFhg6G4d5SepU9moJrjAFzzRIv9pKV+LZUVq6I4b2+mj3OuqDA
80nOc4HG5FrUjYV87DT5qF5r60mu6ODCzCCZVDg1n/XvZI9isfoKmM2b4QAberBF
MP6B+npzw/Kg3+x3PiXAAhcePLKptCuF9kfOJPSavMYkezRK1diYwMvEGpOnAtaM
aa6mAb1aE4UYmPmky9pm+Ex1t4HoIALMdpB5RFXIN3/shk2ZrI4pmH4IBGVap/vc
ZVO2zli8QE9E6A86yM+9joNkbEB+RqeqNjyeKmYPO3awxfdRdg33VxAu0f4BQyWj
M8eIZmh43RVRR8Hg6D2+swLdBlYlroON2YtmyGolPIS5VQYc11t3D/KEqZ4QZ1Xi
yuiMTuyXPfxlEJY1ZQlfNiKXcg5naqvXe09+cmbcQKVg/b73TSbZVndrpSKUMkXb
GKQDk8LMkjym9iMhgfwYnI21Eqi1tiTLTgcqHn8av+3sxXRTM5zwTRil1XKMisQ5
5XmCXYh4P2Z+Ll1hWR2vb6J8l9Dwfrp/Ej2jPqTXGwjitih/DAGwCWjf6LemKNTZ
/V5jB39cbGJoPvRYaEmf9FXWo2/uiTY9YfAkPJ1Hdh6Zj0n45H6zZlioMCKhoplw
gQUorD+fxv6vZl3tKWFy7iCo+RFbamBuVhpmwVYmzv5uzEXsq2f7q2PzFOSHbgwM
dQ1D8dx/FvW6PY/zf3cE6ZDRf5VqJi24sQCmekra1d2UWcQzKo+D6rWeXruEQ+7g
hUmgMVUHBpOmoALsgOoqXT+eRKVjY1j2weG6k2yXZFb7nIAYreBEsnxi2YsrJd0k
6YU3/TXDfAytUNaaxTp68rEGeOGl+5DEPilX5jGPlAZJcN3B0m0Wjs/PZ5CEv1rL
QTB1xZnEphD8mJXbw6KVNpuUHTxPy3VeLpKIgDQDdxvIDkmO3JdaBr6Uvk6loM/6
8n3Kz9K/facjKaVlD3KVkdDUeqHodWAXyASi/AsKjZtZ5r52+x5Z5ZqQfATiHumQ
RJBZ//V5wE7d4gl4cob2seCyiQfdqgcd94Uww0Kr5u2yCR+2shwCTfPkHVE9TuXj
sj+GC3pmzsQ7iPI4XtnbogYGMN+I9i8Q2FC21cM0RXafBUQW6P5xYNMXPjlNj2SG
K7t1f/oLLSPVFUJkh3D9jZqeJoSAd+iS1my9NbmCRn/35A6gjHcUltXYmA8RwnvC
FVWwiF2MFeIS8W3P0ki0J1bZ2St02bv58hScwyyu2I+eqH+0fj89VPxVk4VnZ+GV
Yes4He8XC684w90a781XDURZwKexd2vH4ef8sU38Sx8XfM0gKz5jbZ+Hy6PoOung
EHguJNzqXv9asFwTYdGHfoXwZbeebpY2pHmJZTNW4H1BvFdOkg4p6ExMFmFLlRie
FEpC5LeVTJyNDD2fJ2SGX7p61Cf9rIxYzSBVp7GfzVsjQLzGdX+CLotYhmEIL9ph
Pe52rZSfYOb+UVIafAzVbfv6SddBKnIJWH8BBftsodAggmVHegBuM42OHFfxuk3Q
fHQSzcXltX3Srtb4ZVikiqmK2Nc9EMsMrZek8CHqk77brSj4zXB+14oyiFXnM21K
730tK8pcaXwJFZV2k3G2NXjvuBmOh7gU/9WXXw2ibNL4TPHRxtSxzOuAmJb9kdsM
CEejJHDP1O8BV8GEi1vHHBnLPgrcHB+y25RqRS/B/T693k6q4neSlZML13c/NZYb
vnywv4VgtEuLX9HptpG0Xd0JuFjBFocVWiUgixq9UHifFuN84lcR2w75AF7wpEiJ
DfGQ9eFY50oEGm2XzdJu3FR45AP/OER10XO0ckxc6T2liLiv1iwTctO1MAmOkpAh
MgNWZVyesgUNGy5v3+Y49jdYMyiMugAa4obAMbmULUB1tHrUT7ULVOW38sAcHJ3l
w+q2xCm3lhOFupojuHBtviMSKo9OvxE05bWpTrybRu6cnJBSfbOZWlllfbfiL53T
x3xZmL4lSSyatYRzO/3iFcPyWuMjmUJa62Ec63gH5WkV+/OWUoKD1Rc7z5i43fJF
pAtKGju7jI5m5sOJW6KgQ98zYlNS/eu6+eeNOdLPal5C7WtWeyjDR7wQaBtDnuDF
CnuQp1CT3iD7N1qLvnhVYaRGthx846pHeBcY/AT6SUaRQJ4ljkJQpi+FpkcZU8mw
koOWiyi6/9NL3kXecgsZ3t9SXvBnvmQWUfWkQqc00oZAZwUQXwYc1bGhDbfgBkMu
X3uizUIUSpnciWtZOJsb+1SOc+6Y7g+8ZS+BmhkxqAk7cv4PTIgXpMuGVlj7phQ2
hA1w9d8oCJyJ00OhCm49FKivOeHi3dflMoHr+i5L775yZBnwImUVqrFRApeVjI0h
n8H9id7jW0izQF7CymqKbbwTevMtThLj7xVZNlkw/LrhQ21uHSR0ie/UjPN4jAb+
7lgL/JvSSxZAg+euabowXlg67IIT4LZZIEHxvvFTri3wvQaoKs+E/BUI3dy1dcM+
IM2s0vF92qU/IEkdK3BM8IIkA/WwD/9MHxs1PZCEKEup2G+03is5mt+uIhxujGo5
yag88JV8Qg9CIPq39HHSvK7Gx2lNRZWEsTCjUO6ocbtA/gIwptTxVQdN49XknphR
cXPyDbKIREPzSJ9ykT0iAnU7wsuHDqUgbVe7TfwTgXmjhwoVFd85+RlU69lt8X1o
YxD7f+MQ3hVzZaw25Vs3I2A+EmhdRZ3lqlRjxuSRYIa6i4catJg6mLzEXrFapBnu
4ihVdwBAlv5+cMV0Mkjo5enmC/zm1efUEoJd6NaRlqxU9jZubDLPSb5Qd1Jsvf2e
/YF2RCaRcUdcosYuZ2EOV/br0Zk+JUv+12EBm7cYGkCniYbSNSggqFvr6VyaKCG0
iSkP/n88wQFBo4FvTwgSOpXpe/+gFHyt1lTdaHiqlqr1w5SyWYVOMJaAJGkw1ceD
+jD2S8Gj6bgQQcZOCApjLsGKCdykAoL+OGturK1dbK9bBpBIOzk8HQAbqf5fguxV
OYR0GTAltdM6UCj/78ccMUaGYONjaugjBOOLD4cIh8fk5GAOcbdvWSlD2Vnk+O/E
FZI824PfZeZ6Mf0ylN0RbLrsfycP+kMUSb/vlcEliKuAvveAk+43gkp8fzOc7Dby
0Vifd9QcvPAoiafVzBZJXcD3RCdwnANFom6i9RYzx8g=
`pragma protect end_protected
