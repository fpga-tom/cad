// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:22 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
U/Cz/QBYVI/Rppl3o50OQga8Ap/TMXBdKsl1a2LRG8RMXr6TV2M3bGsbxkzCUd0O
n1vJw2J/sGK1r1ykQdBv2Z0OX+zoI/hC9uM9lZuSdhSMKAtSdx1mn+ZB+c5kTcgs
kQWFtL21BhEWkswGQnovZ5vGPOwVdY/yDBpXJ4WFOX4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 49328)
juopbp9YXPinEcDILqhjMnF0rZOG61EQZW1hYe9KbHh0/zBWxAq6hcJNb1N2s1fV
dpknToxqOad73vLi7EhmdKsbQPBhNyb8Ft82r6EvC8bWpMGqpkhqFov7g66i/uHi
kv6kjZoS/aDmzPkneMjJYtlPY9YdfZIzB4fU4sBMPt/CRiob7i1Eel7UoWBIPCUA
5IV9SapJQ8SD06ch0qUNhM5SkAvQ2/aEGQ1PKpQNGS83gVTcsx7mt1WTq3l+JCWr
cBNqdWk8gUhJA4NxtlcCNnnpnTx/ZELSNx2qQKPVGCA+83KnQiiOhYvFDurzr7Bz
0xNQvZAXJuJn0jRxIfd5Y8ak30J3jGHbi2lTftQKJ7ab2d3e6gL68iKSiKgNJxUR
NIV1/qFzuUDXEuZZojmuaSP5bzoB7bNesxxXnzL79P5xIEwL5JhSmNweDmCplpJU
i9G+7lo/IOkh7wq7dqXGyqdX4qblH8cdRz2kTeZy+EXYuuV9FMs36oi8vGLq4Q2F
fVdrHMNe+2luv5h6uXhtvgKqGRuKdvk8+a8byzYOzd0jtSqRp/JvTb9cYXiuJRNT
gmCUcaQyXqdhC2iu/fJgpq5RewfviqoiIzDHHeMomRtebaOp4rYbEWLa9UpXkyhZ
vQ19pxaSoK1ZDOzhbqNWVPBxiYqiex/BBXJy0QSaZhG6VAds7ii3OZq0xn3h8lky
GCOfRjPm70kwzT+mDZqM80oOjdBjsu3Py0wBtkgzv3F4xAhXtp8/Z8WOGr8HqHfD
SgPC69UeLWFHgqhM+YTnGcNH2mf9LZWNxqfZbekGTPZr2K+MmHv8uWBNVyQSmzQI
hfCF/jVwJI5Vz/FtzBZgRXDWdHYki86o+qYRjvoaB/RXu2YdK1t35PLH+f/UvXZL
JDuU+xG9X3dYyQifiyfvvszQOd2ZHd6Kak9QtjAekO76tQarSMpU0wmBL/teQmHz
KMCbz/seGRy0n0x4fAL4/iVj8K5P9ex7rghmRzsverGOccXNJi5Zmiq2LlH9eSQN
VEyNwtMXoEkmh+OIWbJE67l3dXM92D+gcF7Nm5BLfObNba/TPs5D6p6ttBVdzzJK
SWBE+ymsbV3rF5ib0x567okmaeokOisbv/RtgvVro6mDgcSsAJMVzeHJnoDVL5N6
A/YUQsF7/jEwrbZGqSDX4hwTsIqJjrlYy3mo3UMVyMnWK3greCgZ7iOlN5HoQ/y+
nGABFsdG9ZGAOrPOrxJFd8mkutH4n0vgy6MFWyptKC7k4iddK0xl7PiPDPsBBOYl
gWDKrRqw7XuvrOl5Pxa3qF12G0pEc8+j3f4hCbrCY8v62vk9VLd0KIkPArX7ToXZ
1pm5eGFtq0JCpgZCxVvu1ysMoXzJodJvl+H5nGYRMIWCs6FKzVSDEGsWBLuNYzTg
24A8yOhU1TK6iikThnmYB/BCko5aB+HMfyx8AFFIUIN8sNpJ8OUr26lZxUCMB7Mf
GUpwcd7Rd6EDBDvQ8q6kz8j9ozHs4YRW0rCtH8DzWyoJ9RAN1sphKIU7YUUpwynv
gnlnou/uNE/KlO6IPFdoPs/sMfxl88vXyVmHCslBuRnoPky4MVRqCikMpIy0Nh6e
5QQr72u4Chn8Ik9t1sVQ2uSqPmkv8Rsbc35losipVloDul7U9Ifw6PO6XnWEQyD9
cIRejYVA9zUhNZcG9bNjyof+sZ4Nvda6aH94luOOFvCrVOted2sUCQev6/xnIZn8
1kERxcSGaU5DHYS96H6XrHf5470IbU3L7I/ujNE7d4s51PXyvP0kyfnTQgS/5l4y
PgpiEA+Z5dEaBnwqitHGhvkl5/OidTU8k2QwdMYdQ6eHoCleqlIcZbusB2Do67QL
WuTntmlv+ZXwY5UQnphfJ/gNGPjlR9RkxQY+blCeE1k+Edac977auc3DAPD7M7rK
aodybXNQ1NPIRdbycu3ljgNXVI4O4bsC7gpwzkMeJ4jP3pC2DfySfHmZB7FCSauD
+s+buBiwr7AZFT89KVOiYA2ZjYjzLcM4W8oF774OSKHqgl/MBhI8XfE9AuiPlKCq
x9y/GFW+YZkE5lRJDOUxqrGO9C4jetvPzDa/7Ax2F8Zv7rE6GbpmnflxWeTfe0gF
IdKkZcFatlL9ZQKYjb10f7pFQoTMbEzE71qEF8DELg9gkvJL+/4pOKWqjLYQACRA
lUl4g59R53cRAhuNZrEYHM9LgOkFU6Hkrc7WznxAcKaCofUzpHgWWVC8QwP3ofoy
ybZMH38Gu+hhhj0t83vbiNwyGtU5HCg/VI3uDJeW77p2+CYJNWZhgwJ8Nt/okz8D
5JS0s/lGrhDRKiraMrcALNL7Lg5Z7IYAMbDb1Hl/iiSGj0X3Jn61u0DnwONXHeA7
suXbdsDtA4cfn4hA0+NSnXssbHtuvjIq9bP4PfjJhCUcRuNch8KYYwbOKM3Ovd1Y
UDwguYjfEihtdVv2bDu6ggn/gqudh0fG0bB8A8txteVy4yFaFWbh+l7q6tvu222Y
hPqLjSEjxCEkozlxTYfAg4hqvcNIXPBtRMwjMUrcbA0eK77uSzu1VIVZchKyiTeH
SAsTV4AvS9itVN41JKNFn35hyeUvqwWlRRrlKjzTGEJxnJgG6bjFMrnUI+XaBp/t
jXuyWloyLchFhwrmXVM77kuxkhuxVjhduaJAFqKRRGDKyMwt3nTllVoiYemMbxqD
6Nwhi3HU6I0xuC6z2jsBr4qHNhqNX/aRvvS2Jku4qPLjkKSrgfedtBrtKkl90Sda
EHYRyIMV41gKij751kc1JRrfpZKkNeQaKNBd8Wb2B5Vl1ayFaQAFSc1X/+m0uEay
JhIYXHU7caIv+AREz0rSnktK713/+00w6P38szTMkx3OqMqvXyuIqWbIMJc3747/
6/y4q2pk59sEmVciRHJ4YmO7XY7EnRk4sKi2Ha/hyUw1yRU2wiF8oyZTmfnN3+pQ
Nm2I1zA/GvcAdL/tRPiNTkWZ0KW5f32qFNYXWs00+rnqxmAYsPjPcqthtdu20bcN
9YTVLRqkWCsK8xzJWCrYaqzrew3rJOeFriS8MmxDMCVI98lI9taL3E//xYN2cXmV
sMWelZ8ZdON1lpTg0310wMM2qTWql2qcG4nVthhMaVgIitcfbypLyhcoMx5kdiBo
0n9vjx/PH4/TG1cZIAPLi7Gi8FYrx8Drp1N2Ej14rLsIHKjcFqpSELl9ZyVCAElK
rjrksEDdX1NhCk1TR55pWBgMdbaidS9cM2bbUzonjDreaMoMjFQ2rCrHp6/a3osL
9pPDoHQlTdFUnALN03hOk8H8RPnQXe4pUOo4N0SbaVHhDIfjHVAiqRf4VGt1EkZx
4ua3W1FRS023swjD0Jf33gzBhCxVP2L7gDESW0qNYL+veZl7pQHdHt8tL1sx2xaV
S+wAfP74MjZxgBMCMpyQFYRADp5w/XbfH2Lk44UKw4NgPOdj3xMtVTpx5CKt1foj
t82QA1qr/iAU1NQbSTn4vYv6EShmcUVpRfAmhaxCs9opxqMxqC1AL6EkVNRxcsN9
lqAUzmzFnWkd7iGt8gN69Vy1fGXaFiTLtkVcHPrL7ER/ujY3ooUBvpf3SCEGulsS
UFy2ppTwtR1n4Pcf8H/V2UovYILTVA5H2/9PPLFOBo0xUiTyvtuRKR1BGOoYDj/w
lQdr0XqMOIlev+qx6V0lA3p0ko41l92B0CPhmMIrZGUzPPCjx3GSgn6CHr0Q2/gB
T1e5EAQ0bSJXE1xUDOp71vzIPSDa4N+XsQyH2f+e5tIG8KE+DnyPr54IEV2OE6gk
lv0a/cn8Qw9MwopoTQBLsDFxov+J+aKFY3zDHP+9J9pARO5CPqv9cHaO2QzEnqXn
Jrm9V6LeaIlBC0filZ+A/9PmQj700PEwEOg88WZlUUaTrhxhQB3aXAHIc/fTeF/s
RVrlWnDB57QHtyEv7ngoDSkbbfHfDd0JIcapreFuUqFulgtJqacjZhc3G/ZVred6
Aj2MTCJkIcLc4Y1ajYoq7BfdLMWh4iGQygiTFNiPaGngvFZYEp0hlUzuMUaSnTYs
9n5FWlcdvfAtZisw2lu0lJnPnMZjAE/teHK7wyNBNojp9r3QvTjOAuvDZ1WphHnQ
grCThr3x0tv1zpmFQ5Pbxuj+PnA2Gaodvq5oUOT8nNy3jUw8xGwerEGZzNV95t22
cphD+/QPJTmu4FZhOpr/npJMMBvJrtnlkiCRyi5++Kv8VUhWxBq2W0kVtvVEm6F2
2pQsW3dvbOfGIRYCOLd7SrEQ04FjpYGkatgx3v2uHphcZsvIm6JYl7tNv26CF7UP
rvVIcLlaYtX/FUGbN7fEswyUiCIG5hNeWOWAEbz3mI+p/oVZglDCkYcEikVWwrMu
JYG0QHX3bAnR61WsDrTG3FFZJryAlgp2mCcdNoZ/01L22BNtp+/KyNdAhupGBsNu
a1V9kxJ0S3gfYlAmmVY4YzHDsCwyQS//hSLaw/cJchcTpuM9Hujzsfri3ke6AEcY
wfnR0jyc69q5X+n8P++y3AZDXQFrhMY/54+fEV3hTgLqwnMTiYe1+PbcJyJju6NK
5aqgw95kPAmUF8dULbPcHDkei+Utf+KjDCB8tyFBt9BV1p0MQo4iPjaNkkjHPIpR
W9Ce+RtpcZ9vIK9DappM/TA5MMegL6kw/wUh+Tw9jiMPV+OWYf6cwCiDTE4nh3aB
eoEY2SPwGylYdOca4XArZw+lb3MfhbEQf2n/j0xKOsg7PJr7G3jwRV1eI9YzRO4M
m/aVDMUe86260mgyHaMR6vX+qtoAnsK7riUqPpqMS0FOvbsbYIw72TiVT5qrd749
/HCeXDxFIHzZWNM+VSTKm5vi26eNSM4H4IbnbXvn9vMSznW7O6bteHXEIVpK9/3M
Tyej85W/9aOnE/Dd4V2HZfv+kNcFd4VVjijvNpYL2tDevS//GmGqKYFRQ4VIbUAK
mlWlfsUtBODgFL/Kwlzm2UKf++iGiaV+pPb/As/gCztbnuDh1Tphk7V7kx8dyMwq
QMrIpL2nObvNjhqL02A8EirxDtpkRpLUD9olN2rZQSoDSkaFc3kz+3kneyXACHkX
5c2crF+RkKPqUyNY0T4Kaeb0IVDr6aGuGCDfALkZbq1OTkLmechSA8hHx9sVWYZP
V0PUfGAotBLfeL9i96SG90VHK2uncjgAHD/t5q59Kqvj3gjJoX1nYKz2vplHa3y2
3Ufy93DR6WkfA3oWtyPDtu1d9nlBCUTVFMt53x+2cDx0sNRMjoeHxxsOqS67mS2w
J3+1VVskfCDbIbCz3EGSUEKQaVKc/MzOVQwaV9mcQ25Mj2rf4gMNyLDoYYbXKaL5
Img9y7vRztwjx07paqin7Qe/rvOTGtyF4M+8zZ5fBXpyvOwn9rXgRkM95Yo8O9Z+
TNAr3EOipZKlpWit9tgXV16dyp6H9YzGriYWofOh26KEWOnTySV7oN6LukrCTVOd
Sj2NKnB0hMZ/MDSOuHyNMbmTqcPghDFrwJdYQlhg4Nud2f3VAAwbXkHMmqr/4Y6v
Pe5DxTTZ0Wh4OJ1Z0mIEvEF2uwbDokEj9VjGVD+PLV9PkRBX21LbY0mW83acq1Hj
XrkTS4M1rejTJpt9uP/+cFVC0SLXFqZap7R5SfVrdAwPDJj2voM8tqbTqxi3hGdU
+X7e+JogqPuBHhsfzFCSMKLZe7qvh+NCCfZtACK2uO7Kl4YdAseyduA7YPBvBMyW
eM9sVHrV82N69/m5zxWD6mZuQRC6UE4LW6/naCVcA1WcglISLGzscZMuoopns1a0
HYIIMw7jPWwiTnvPQW2lMUxFrqY8MKcxYQVd+wpfMNaGJVE6cN8/xAj/secshdTW
qQm7HAV2pTzTcs7YmGsFsB9+0eF6ybzaYK2ZgCPY4ZGJakwydkvv4OdszSc26BT0
Kj9fSSzmgdJ3vKhMjMp48haC9wdCo39bzr9J62bcVV4+Q9qkBKtKYhBkP2nG0eSa
va9zwYSwI+y8A2TJFTvNDFnush4OabmexmVwIwXCj/zkcJqJ7sVeyMr7cIsc/NNY
p4Qb/3GoV2cZMQcHiojq1jfZZkYk0RLYcIwcNzvAt2o7KeORfq5rL7XDHt1ZKyih
8ozyL0Q2cscW8FH2ACXcoIcG6SFMgFSDrF9uYo+D3FzCeGOnWrU+81+MKEH7+Ja/
LuQiuuO9zLClnqar3wGRysV31D0a8RspRPuPD1Q68+6z5hI/Tf0nFxmabhTHgALr
C+/IyMFy5YdnhFfxXF/YrCGhUgmI1x6uDqdpI1mv9wmunS9JkzWdRnvNeK2WBskX
msNbubMDnnZRYxWfU6a2H45DV71h82J25WQQ1fqlRJzCevzuAGbDb56vglV1y++y
Wfc/NPQBPoHWuORfiktLFigHIDFs2DxxkZIC7zIr7IBtJ+A3vJsY2p02D5pdODB1
iZriRv531dVQcnNVfXnmg3DPGDs7kUAcY8m7SWwjMsfpN/Z+/htCfqzs9KNK2YVw
kMjfyZfChIjdytmJUInPacqGEV1BxsNbYLSFyMwf+25zTQuYfYDwZOG6RvYBvXeu
7d1jveaGcB2bcAMTqT0isAhHpEj949uwbg5uCt4ZHncMbmB07f7DJJh8W0UARo+p
rW+jMWSvAMuMUuUlrVbAtQUHwSad9g5q4CqfQxsrORFPOcIhqPL4oPTBRrwrk/Bq
7rasp9sy9qfmmDBY5K+HbqdwQLAjxWg9oGKnn9fYNJvLzaMlcXI2Nl3xIe2vYSXW
HRPX7B70Jwz3gkQNNn/PVzBNRi4hCvBhwajis5O1e0NkBSwVmuGhMJSIAxQK732R
4ZjxK5mZ57XcmkcoxXRU0iH10W6FYYT+fAtGV/BjUF04rzNkTG7gFQLAAT+1G6jo
MlsI55RYPFuVAnQeDdCtw/4mGXNyrSHS+JQF9tJonI5NwAnBz+yWEx/wEloDZwPv
O7v+jmLR6CI5CoIBoxvF/BUbJy0Fl2isL+i3wfJie4OXpG4EboF7itdtgiKukXHe
oy9XwcVnuPgyRWallUmdz38pz6Qfj9DNmeGePezieldJztON1u+dhtDUyjCtpa37
AnQAlxOBwTlCtxSfPAKD1da8jvGpEtWiCAvfmJEhASlA4S3kl3FwyyfBrmXXRtpg
zEjHztrPrvnc0W5j9Aj2OGHrA0Tv+N4D9fhNW5/MS9LaPKHp4kFVi6s7usVguIJm
qF5pFfa6Js5QnRkcfwUBj+dPK+fIb6icptvgMwCazx1X56mMqmyt3T6t/f57qrau
icu5cUB9NKg662/HxVJ981HhcYefsm0yInmPb34t4afluXzAzVK2QKiuBgCnPPsa
jWjZtMLVPokYuE0ra+6KlZ35oT1y4QPJvaaGuciPf3GQI0AC3LT5DTEB443qDXuh
tCGQCS5r5pBgUHPbBNnvu5ecypXFWBHb8Q8nat2gVguYAcqnGWhjuTOvhEQ/KbD+
31KsrqCYv4SE6mxg/uRu/1Xt9Jo5chJboQsh65SNcvoYAYvOHjn2fe7wkr4FYLnP
TkAeZ7EUFSIyoKuq15uotwQirwI2keQoIzVyAv5Eyw3ArLgIVQvnKu7isacqbdi+
tSVd4ZT9RGgobn6g+XfDESlzFV/eiO05K7DZHuzTa2D86JKl1pYQ8re4AhlhQUAE
k1oYx5Y83gh4v4MFWEgEk8LMBgmtMwVdyY3R4Ze9PTyRtmD90iic5zqD9GTIsckT
ZBixp0c6d+SKzCEqYDZg+Wd3xKq20hxQ9Pzj4kveoRts32/+6nlS5e5pqCClSJa6
oCF0SDCPFPSq3MPSrZSm/diQeO/5usG2/FACEZGBjm+ah2B8pzAfiDkZCV1HPw2c
vlD/Sbghcad3PVLt7/PqOfwZD1vScIXVZeKExFXQnxNEIvG0OjTy2L47sym/Sde1
CaJNpKAb8oqMmIPBSSIAEwJz1UF7RlbmUEgXp6P52t/2bdo/6ft4SUjgS8AbdJZV
iLfV6NH6YowFXlrKjlavsyciyAIiL6sqbEymDuZhfYeO/M20PD2MGel0IGqQ7WQm
FwShC6boj89R7Oh9ULjkJWhNVHdus9H/MXS1/SgHcNWK6cYKLX+PH+3aeCGYJf8c
zEx370KBqYwrqZPWYQWMBNGisXgs8KBmylXvBCnzo+dihv2KnUD7i2eTmwUC5hOr
UDwQQiCVtP1tSKrEPlRtn6TxJV31wRQ2CNkDCCVgFfY8SAziDoUqtOPsDbGDaD97
Nva716rLzVAhJx+/O8FdiEVc3SHLJZcA4hivJpm1tLMjgP9GA8IwGCSz6dPZr4Ll
WTUNERvX3u9gTBPkDae2LeqwL2WCbr8q07hobXqtsYMouU7pT/ngr8H2TLGyKCoW
Nkamv+K8hsZzbZen0gDRWqFlITmXzqv1oUSNLMigW//aJY95IffJNwXl7Mv35XAJ
MZP5HBz8C8CVmhu3BmMWJABVjEIEwC9MD44+ya+wg7qZNB/CyR91SQ3c7qrWaVgX
GmMGsyalgQVN6XbiRsWFo0r14HuMdQjro6cruMYdWSzwcz4rECpYA3DjzlzMrm8W
ODOZm39KGjtZlllRw45s9/w/siZbZ/GKcSnKG8RPLk/Acw3sEL+7DakCdGBY45Oj
XrcfrGCl05JW6rjWq7SffXBRVNwmJN/3cCe+5fi+VVKjHgqrL5UjaXJTCg+ND1ei
/GSoA6x7HyWraG155IK+ySg2R9LCpRCzaYlc45OFJPdM0elGBvRrH1yrqeqDa0/h
Op+RYA0skKRfIrOAB5/MOK7R1pi3H0zx/ZFS+U6ElPABOFBroMajS+3OJqi0b6QP
mFqAELWa4i5svJoQ22rIxPYJj7djcudO4PZQmjrDyzFZGWq0livZAb+h7XJjIMQW
dUX+9VdFkqIXrOpr36ugGUHTMQYWsSuQxzS2eyY8VH/UsUI4wqLWPBzkpaa7TsoP
6GxJzVQPnYR+V3fkwFz770qsoJoZ1Ejkh253y0QNniEfv6Te/anlx5vKqRV5sZ0C
y6NSmy5en2ZzMds7DDnXoTQ+Q0LmvhOyB3hqA1iOFVO51kQCEvL0kZH25EnAxijK
IEnTAdpOqdJgikqWoLAMPYgaWg96TuurUb7IIzi9hOvd2IEX25GDKxPH2cOQD265
naNT8vCjNaqFJma8sDpWw/akv1cICIHv21Wh0VKkLBXIoOkGU+76rYD0dV8aGC/L
R9AEF7EnYL+8GDeBPk0ufSGNUV0b6tFPYQIKMQg/VVq/pZzJZ+cE7optjNjeH7WJ
PyjP7t2w9aa1mg7ryUt8ikFajDWVZ6yAYqcnsgaLXYWHu4cXmdLZDc0Xm+qa77yQ
AOASVJMTyJ4CbY57PSnSkYokZc6sENi5sdHTSfl90HPMjZ2ow0ATmsWwJAZbTg2M
Jqp8Qki8WH5VbYJ5fI7Z0rhCy4WvUWuTnuuBD0tqLCX990VDOg5/skfsuuc2cBA+
CJM3dLi7v1osgqXHmk3pMNLeA05icu3rjvxtpmPC7tqkb19VlTRsTzljVHDINAHq
75M21O7WKAphz/5hOjwTik9+vX0HJMqOrJlLj/Kb1m6TDN8VOlSqE97CM8Dyh6QF
iytDmelEuuMC3XZz0CvwS5ZvESkautqOjRCzFQtIS6yUS7zHqmqpMXvryAVESpwJ
MVu+5CWwnlo/unWbZjJKaKLWhqk8p8/xj2IOF4E9oMVG7PLnTFRkMawoU+1PSyMU
QPz9mxcmle4BNz/N1ba5hBGC/OfoJ10y7KGTVRUrs67OKd2w3EzdBYm6n9uZpktY
uUXnR8vxWevl4GwRXDM1zbE107sLtcqZ9wapFlYMRaSLszeGvNStg9Z1UxHsyLB3
2u7Bj6q74HXFwXdElhxn3SEUX767wcpBrPNAA51Sv0DCrHiaw+rs3BLhIgcy1NuU
SpIwkC90KuM/Q5sTXuXp7fr6eSvJx/rqdkpsdpQbZ5mm//mDfo7Pvjkqjke+I6Jx
xc1LmuiE/VzV6rBiyE8p+8bDV4R/yo7OFh2JyAJJuYpuevw8fy1Dj3ihuS654cuv
f0rWnghpVW+o7r/qBB1DECfsuU0L1jQPT5JKLgkfTlSi/uiCwWA5u3Qs2l2p94j9
XlhDRdv7toTvhSAEe9xXJOH7qFXyj6/l0DmyoCPo4YYm0U+cRGQNBcCH3+twpW/B
Hjbcf7HZU8a2yR8cCSfb9GLHd4tsOGHDh/LmntTQuc/ebQbKI0KYUaZvgfsV/GPX
a4hVHrNVSJ2dqp4Su33O0EYxc0QouVePeytmDq6srxlew7+PNzPDfM3Ly3tv2c0Q
oW2L0aYbkecLHPrrEKqTFNnhICrKFBIoF/En+O+WgSotyXX/YT0riD8DnOit+Xd8
E8TsDuO0SfIqXE5+eBfE+yJca/IT6QtqPpQkApzUadG0pKglotcDTD98qatC0DVz
BrkzLHjPiR+Sub18p6EQR2QHdbeJ+YMV9FIa2izO2YKhvHoIXQ8BtCfZKhmQw4P/
/yWFnOk435TvADP+2FUPiIV5lD02dfAM1Bxk5FIGWcOaQ8bgwvnx8B8E4+yEvCzn
SZnt5MzucoH2qrGdKZic46InXAX6CErFCDUVKAimK+k6buL6xHWuc1+YNYrHj/3+
C58DrXtSMiQxHNTP8GdIC7S7oUcyNc8rwW7Tt8rBOcjoFgG2XkE0A+vHMTwQ2iVT
J5c+dTZKr/ekdPneHHFvtB9YBw8pGabn9UurrS10tCIV5CBSZNPT2B0MpP0drVgI
JMI7rZPtlLD6/6uUaJu7twBANjPwtYXs03knJ4N4hElZkE+XmlAHpwQDXvBkjAh9
6T3Fa+JvSBYQBfWSVj/ntCgy+wjvZZfMzcZjQ0H2wVYyavPyobtcnAWGnzeouXpV
Bn63HR4YTt1dI8CpxDiv+hob0HBZA21CZuyHDqsGDFabZ/FSscKvOQiTZ4yVHXj3
6sKslRjwpiAX7ebPodeFppnb7YfBUpw0ANPEu9x9KUttC9dfX5w+/bm5ivpB5vOj
l7jI1Z0QqMI1d9+CtcZ3msyoJF5/v/YIJDdWf/YKxuM8DDkmSA+WKJJyCwNJcqxa
LS5EEKzktbBi/hhCRpDk5dWRHRvElCjUw4ps9SZO5kP0+PHkn8UwOeUNy8eRAARS
/CFsmyz7GI57k9NnTNkqhyhCbxd5aOU764rR57y1EwSBo7NrIB4Iaw9ncKSXjsDy
1inirnEYxTaR9XfspAlJAHUmenEPfEiJLBtR5r2hDsiqHWALbjDPi4cYWRFk9UMw
iw513Jhr0tTbjAaU4jKEBgdUbeplKXbWE0D+kECHq7OuYnMZLJo/4DpK2ABp3sEI
cjGELpoAxrskBWip1J1f3avhrdwbWHhL2Tvk6CvY2lH3FjNWnhGAStF9Y1rCUbWJ
7FHrD7w8e1xg0tUscKaawyHRyacRnlHKRhNBVsqWzUweqFTRGogMvpP5H6SxyWEM
0cdmDOldXpSui/+X8CICxSqunfp+vx0ryqbJJVh6OrQV0rXkr3mLJLnxb/mXYavW
ptIemFvliGu7ahAN+canzg3XDXm7jZ38MQHKWdu3OSc+dIUJf9/7RA0qwuna3G//
PRkDPCCLTohicWKme4WwPduUThvbDqrI/csoF20adLH3cB0hTSBL3MUpUF3J7WmP
nAhav8RmgTA/fPw1xgHW9CJNztIkPKYxsq/Wj+TLXr7BeRa6SHmmkJ9Q01u1TzjS
RNb9ebiz5EJqnS47xy3Q3YVoJWJaHuD3vHOgC33L0u5LWlqjiSiGBWUD7D6ycvQb
VS8j0t8ShDGkqtSwYI23CSYsXFLOnvQGtAy3YXVfMOQcB6JmvcGxLW7aykiW3aQi
w2oWQc7WziEuISosx63aqVvb7JvQFjQqJ07KgiunGw/xO5WzIUVERQXMEJDMBfmC
qjf9qju6zwTfRS7sOVf1fBVJ7KymZBe/Dljo5ktQq7lFVj7EkSGMp3oEkRaBkXZz
FTGJyHDpvfXYKVOaLntWSzA1S0akif5JpYJXKUpTgPKSGtwAaRqQPEz0lRY2qzpx
imrewUdqPyLb9tm+x8VieloBnkOPZcTlqcBtTrq2e3nAmCBlFWMgnH+3HG2S9lh+
HzLcHTWq2LlrS+AOYGEOSoYVXTZVGJFHOqhZ5JTpwvRSmyfj/3EovhL3l5KttTrK
wwaeBjzAWBS6vOQVx0osgfjVCmqd+a0w0KdNZ3vWrgIQUGtvHHd1+venGleXfJWQ
0srVtq70mgu2kWjedkFcEPdaLBZS7vk59WM00j6XpMqDjh47JFUStvqaXZNDrXDS
ISpBOZzZgRSXGzc/cPgifFHQbj78fmho5eYcqJXioTqbOlIcV5ePqv+xK4xAdjj8
OeHqRo+6YWD5LbPa8B5OyuWWCZv6Jbhe2Ny7ea0m/JEbn7VmM6Ol1kALy2qUouo1
vwAFWFAe8fphoBu4kZuYiS7RxVJlfSQIrdh6dkFU/Ww3dq27Se9uaGiGZnzCwzBI
Z6GINF1ou+I/cG5mTSOeNrTSdQ9FJyeBgWH0855oohS2r790tn1owMWuk9ydmxzm
QkU/NhRN9ZSqYAmg2kd+NwSI6Gp/JsP8rLmuItt8dQiOlNqBsXhZfMnuqTfyJPdJ
SK4hGi/cPKaI7FH3ZXLj8UT6vPap7cYdIcZDMva9avbOckgyapDlWGKM7EqqzB2x
M5e0htOpilnJBF0WIYnDA4Kf4trT1uZTsXmysF+SY83swz98bMkr+7ux0Lh48V0A
Zru0Hzcsvg2gSjQ3VAtxeCHj3UvPgUI5xz4pJjMjySYa6PflyePym0go5TkjtV9/
2gw+1fFMOJskIa/y0sOGnjBHq6Y3nXW0F92CcYjV6JVY4EigMcfooaqwNdkCSYsO
gyqBGXoRE7Sgqzk4TUdG73WsqNbpbJX+s0bi4EPfD35kNAqmyKdxBdBPf0ITPpbH
ORGjq0RAQaMcpzHYnQAimnTM1vRZ6wnsrLkTFFWwwbsvC3AIdnqPKaLwBhKPDnZI
lpnAFaZGcbcsqZrMQglkvhtZYLCxGpLE0l+Ywwhrxcl4U1vrCtMP8Qn8QmA71jTr
4nXymOusR479MXfrx4DcXOp5YdcQqHrmn2Qd/Xmww6Pmeoyi9H4NHvvkfMHw4CgB
ax+LvhcyY1fawkUydcQPQhYY56FbrbNq91gtke96dqZSy0QiN1mWgdqR8WwPVoom
pZB0Io5TuUWg0nM/i+soRSMgLX73rrUI70+Qex3UmI62C4HLLOYNOLOr4p1iDh40
6IYKNgqiJ8YB+ANbOeTjgBRVlYnwfg5M42uJl5dt7MaObVRtZspH2EeZPJ5vVNTF
c/sqKl88zC+41OG3aLGLbwpjAhyuyiAs8EnWbLm9DRk+98wrc9xtRSd72eFjwBtf
jyie5HMH2g+F6SW0II2A9RFUmnw1sKrIZ7q5HpY9BqEbn3U7b4wKu62J5leeveeu
pq/h2rad1SnyhrAP2anoeGl9+gJ305sfPbqLLuyYdjKfkmqJSS4g7Q7NF0GMmVpf
lJCjC51FqWZck24Og3MIodKpiYTliDJdN6Go/QYF4doURraHA8Il8JKDFi72S/QP
hBPUp/e5jdTvvHEZQY81iqVCtstZgL7BzjHr4xqReRqvimm/Z1eJljDD2RFONXS4
xQMZSGn+SrKQjzePvPNHdnG359luR//zhiNnChNfFazqG3fqsQZKsM/YRyzHmRtY
SnmSDfZNb16dGTRmi44NbuBD9jRGugBxhRMchg0FiZQdmzgRc/e7T24PrMyFZ9xn
VLvbebFWc+fIhyhfvce6ys83qU4cMxiUglDGaFlbAf03eWbk88SOdLwECOElZ6A6
yizMX7yflAnGDapkR/XGRom2GBiOkNlwEEnvJpg+PIJ/IKnktL/YWBz00ub21xgP
NLFIUwkUqXbh/HQ6WofomPLXjBE72MPWcekdfQFo96/Hqrlk69diEu0ER67XZMWk
cVVlbIFkqmMGy7kWlxq5AY62anwj1xtaw7VeApwE0zF+LTsnhutueizRcXCmodUy
Vb4xSSNP6I5qqG0GYmAEqhXH8KNN60zjYpT9zdnRqt3Kchi7B2ZHguEoZJESWFq9
j1AVQcUdgyqAC/ie9bsv4jpybNh10qlx/SPMRQf6NjvxmEJkuD2zJLfPqQ4YqESH
kH1gUx5uVFNLDqfJFWsq1yvoAiwY1UGjnIrIpCfLknrGDTd5erzT4lIyXDK6OiwA
7XK5iuPNEcFjPQuI71RqjYxQv1HzGkVyi+PCn6oP/+AcHa2VfsQmdePN5bjZKjHu
KC4XVNbjZur/HfImd/9olsij1N0rTz8w1pNvRhoJaTerGpyUqVyApYD17E7T5wM/
Tr1eQuR2N/BI56qsgspacEvFB6VRTfnS51dmQ0eDY18AUylbqUqiNXtyWJrQFKE2
+EobY1TQlwQDvadKwHix2pth2HbQD6PEBPQxQoamzb4l85spmPEN2QZg6CeTp59N
fG2DizBx3yqfPMBiV3hCEXdUd6Zp8C6xXR9cOn0a2PgfvfLdZnn4BRbdycZRq5j6
PblriWc7kKEU50/5ANZWmlJLD9ZKVd7ZjMunCGmDqNcEvvdMXkG26VhKeyzPa+BJ
ESmL/QBL4or4X/4xMPJmsYeGMfZ7r058AaKgVJrN1bd2TN4ERObVKYuYIj4octJg
v8R3ss6AVzSaIxhy1AChZzlC4UrGcWq1Ogm2jswYtl5ykXgpB2ewkIDmpPQDzcIx
e/5USHAdK1IH53/TOzw4/HIQrLrEOxOa/Un6J/UuIyPNgBp5L4PaPsSYMmveYHXN
krJcGt0sBfcDK+gPbXWu0YoYlQjn31Sr7rPc1rJ8+6SYoxeYFdvOmUHL5Z8sh6qn
8k7O7sRnkAp8Dmzdr5jCmxUgBVbrvOUtR1tYlkkt3Hd6VixTqtaeJNSzFarWyszL
0UePTvoB6GZpzUBwHmNF8b48kS1dqP5Cdi8pIg3WcFuolDJOGb4ze3XxryE7KCjw
ZNkywyo0KzmoF4tvxwO84mK/rgjEClNGlV2QrMLuO9P+y7PXSpyCupWOZg3d8GIX
LVJA6RwjL1tvqHN8zYVjjsqj2mCGgdV42azto9xcGiBdZZQg/kTsnCsFZvB0njUB
/GyVGbPI5yUdCtSdPRa/YYnDyQXci4xdSVcNICF/SjMoPDigi3x75gYaGGcQnthH
pmjGcykUl7nk9wLdMdmnZ4kkhbaq7A6H2eY7mN6Aw95RbIW4UupQDLQ0lwsdz0W4
GHfh+ne2vr9UXvZTqelgoa9IB+jA7PsCa1TrA70vK+mIM8Lfcan+IemMlVizEFMm
sy+znj4d0FNwY+8sK1yAQCI8EhXQ2lMv2cLF5J5NEOmem9umC2aQnT6Gm/XokKol
q56+1G/02XcUke/8NE+m1gHLJJAPQe/YtVgpInECu8aXer7VVQmLfZ3vIY27neg1
Rn54KACMCyV8Fv6SYoQHHgeNHIDrV8l7bZbRHZGwe2S6NEaevPW9RZ9lxHe/iVsG
bLcUH2DreIBU5JAmqhhLAPLJjzxOJZk7MI0YYdJJah8v6uVnf6FfbRQoj+X2FPLR
7kax93rciLCEwWE92rWaquN7lnDus6NOPqrHJGKUhfIa120YFU2Emi0cwAvw5Das
Nxpa9z0gvQaFA3Y2caMKWlu5PPuTfYecT/fbwUBVIv1MAPKUQxHtmWrjKY1V7XHB
mNehqOE/1dSVfLHB3QuFPgwmuEC9OqH2HagaMz0A2f4K3zhDtq/aZKcmUpNYpZ9k
cXTG/idy/SuHgKkcZlFOg0oEb2PmL25enOHL0NuW9A16nxtxjiU5kqCmDOfmTuFS
WLzNlMpDpgTMsMd0TilL9SrlAotuihuzBazP/0ib73XB5cNY496eYyD3lMP5+tiZ
dZroHNoM+AixoHLCMu9cl6G7JSLB9OE1zpSgdQtpU/W64vslVFIRMhrVYnhF+e+/
oESZDvSeMLEGQNdLECdhxeTR9AjGpxb/4Dmha4cDEDTcP6xGFZMOM89XajWyPb4b
7RnB9xTqKDJITiSZKAkKWwinVNxptx/r61KY/HWOyBl34f0l/1fd8+ivXu1vGCB4
0YTNfKJr1g3tm4NKA9LH18k2Dia6+5eXh15iohA4kn9KiyDASlMW5QTqb6lPEhaw
EzZqsYy4MYhIE73D59n/3H82tgc+FuOqTIEaAZmzUaM9XnFrqz+T5v8h5Q/fCc5g
7ptBy0Uz6r8IhLgaPmczR5ouWpyen9Cel+gpgHkvNIZ3Y4Wcr4x3QFO/Vzjm0gv5
nOiqXo8vFBhsETR2042n4LCz1GJA/jhlKpN/ryB4VCcs9L62+rGQLRs1RIWMQh8k
C5rIYH9mZL0MpbpKwof6cJrIKrmSE8QGIYXYVv5uNwtaMEkeZLdZjwRhwhuiXZZs
SPSkwqT5myW90J0DoNRoja7l2m1T0a0qr7045xP7sc9GWaDTKgVtNSNJItUmwaPB
DuoKjSSX0UYt6ZDO6nKZBOwf1B5XBhG+JQDgz0XjOii+f5uV/rP0R4wAHaoF55/g
6ntOSfG4CnpNFkj77qWNIAP8VPKx634tzf4/NCrsuO6k77MmShcVYqCIedrvigFP
zQY1Bx2pUmfQ5gjyFEfQEB1DG981GH1GArbLy6Ark3px7AfXqHBqUbfFU8q1af61
MrnPXe8DRppsoxHIYYfcuP00r128p/88U0zPtcM+4Y9Pa973C8xPmHCMbpceSzW1
w27nRBHGT+byP9NuptE49fwuVLOCNX2cFFwLDuSUjrTxgG1MNLRuSCRpXXZx4WHc
sse8dY/+QwcZlfnOMeL+rKMQ16DXHbkBihIsvNgzPI6RnhWGXpsbBC7wdCaZnbt9
7BmPMZiuGA5xKdUC+UP4KvznKuISSjEssxhCCt8F2+k82iHLYG1ekdi7ITP5wHqM
U1ztauQ6gl5Y4675Ee5hVYNBEbldFxmrjadECyO8E0MXExd406+ij6szat/c0xVv
5F2FzDm1glj6MzK3QoSGhUn63eJeWFCj5BsQcd9apAzkr2x+4e1vJjhaQ+k2TZ86
Fx5IIGf7y0qWdyawdt/HaNYOhU0Pi1Wz3ylB/kdf4BijpHem+hhF1HmDsUhBXSko
CJsIV7MjsUZD3je16m3xXT7HJcxGaGalWDMLem4LnI/eRfVKqQyCPGwIIoGEdmrR
Umb9byt1Qto4MAHwpNvMdrg5LpZpmwjkinZ10OxD6RSdgknABLYQtWQFXFbmiR9x
BQhPJx9qXUA7bj8AcFCHQI1T4Nm4wvaC5qz/TkfZa7xX3gMRhQS4PAMCMD51sDbf
A6PZtfm7cJlbRWyWW/12VCO8TGAVJhWd1x8+YQ+9dLv/8Om0QbtBrGIP+VI7gqsd
afmbXwPfGee7SrvoVHa5jNpBVuI07Ek/tBgeTJPHsJ/ywFmtQZXcPgy3rlOLlIZ+
3/vWQtJRvJ0dAMYY0J3YPpIJ+a00BaZGSQHezHSDQLFs6MMlm2i6rGKVr6YPcjm1
DS4OXJOtIHT3x9SwXjrcLJ/NoJhYluSNKQW8jM6//wFuZq5SVze8vJhzdeB9XEJT
TexG1wn66yntZcVlSpZozqH2sQyizznIAusGcr5vee+TRt61VvqUPC9sMouOUlsv
wMnbynej8zOmFP81U545iXAufDtjSKKgAyEm08eV/zi1FZVfIJG4fP0+EYbCDwZ4
Ja+rLcIvRb9cF4S5kkDbbgRUczKGSUzvEBqNACBDe+YVcbboFmRz1kB0gNIiU0rn
Gnisqoim0vE5fr8wiH3d6TmXVH9NUgW9Xav28nn07JW8hrIxRXQKubLi6sdzngWU
B97afnUixEpdPz8WMVUG8cgy54Qh/ePuIxsDleCieNU7rqHusE3xLFeElJj5o87P
OAkl9fO30uAGbQ4GxN/fJaimwMqAvfX8owCrfqQCzX/dQFR6znpHaH3EUXrZh0T2
hbe8h94jhJBO8+BUomisGyGaTSzHMfFszeSDLxztPK118u6KX4w4/lxWKDYQlXix
jzPf1KqiQKq0gez2fCvlF1ebSA+heUsdUBghAXKAN8cbim8EZo5XZKaiR/W8hulh
2LtZp6IKKoMXcnminNHqZjDTeDn/l4PTepievtlpxW28wtOTlb0muZrJDH6sPvAi
if637NZs4h4a1xtqL4sJ3/8ZCMyISrn7oc8IoFT1CihT069e5q1QiwmVxKwHZxgB
3+LQe1IsBthAN47hJ0nS4xTgVi2CbhyR+iI/o7/Y9kCyUvhhaO4nw8L1rfkezDkt
Su7U9D6Hd9AIspWb3AXU0YAQJMZyoZVq3VPvFwWMaYE8hrMzTZUIfPwj+/S2x4Pi
QuMs0vffI4sHiPdCSrGFOHAWKc4MfJ13HSAFqFxhyBHRS28JMTPvpzYV+0ozeqlv
ak2tEqtE5yj8qE72QR7cmeht4y788oX0P01S+y1Ke+nSbudFgS2uxkQ1QEg/h+qi
x9S6ZLk4R5yhCI2UKZLmuXBbTuxq0jpIZPRK5hyUIxIk9VkPHqD+UciXEBIyq4Jg
EpvuGMlNZE1qLj4wngRROxFidKtRNpyJKGxl5xEK6BYnWzSBTM34eLDV7lzncyIs
Yo7bGPvqcKo3zv9q5E2Q3RTY427BjV2FgDQzdlYHBU8Es5EgHSZWezr/WIdgzk3R
Bp2DJinfvjPpjrscFKeRXbVI/1j5Qd3nQ/2bgMD1KmuWi8XAcDI9MxUvDetDUXuU
SXr7cSyNKIweD8J8hTYzJBeJ5UUrqfCJLmKL30NvWMtiSHIbAJ7Zh7AHN2sKP23Q
Fae7TxlrHbOx8AzCOI6ZrYnYiLLDR6dvRDGRgrFY49klyYzikbVZQxpvs+ybldyx
+sTEkvGQXn2izvNovqSQULR/YeqGv7cGHEqKoAcQjOBt/1R+4Od6yIMiLcIm/aMs
FUaoZt7gOOeIp+Uudsn5zh5QjaCtAur/oJo6K8lAewLJLec08F5QHBzqQqlI7Cio
NnESJMv717C1N8OjyeM8ZmX/5Feg2g+OHfbj60QhU8v5ud4HMKnbKjLXjI3HP6H8
3vF4V3xcnRUm9YbuLp9KfdUuS2bwkYHitAjb4Og8mV/tN58n05tAyhupEF2eIXUQ
Usu7Qr45TkZSaGqvOF1pbhVaITS6f6GhbGKvKuxc/YJLrot4sr4A/tiqVle6JUwn
GVBt+JdDdt70wHq5ggP89wKDDfL6OJxBjG5kMkrJJCDMlVV7Va8X82Pa5PYopF+O
tRKn8jAZU8CsMSsWxUjJe/rBTKzhQYF5Fq393IRwlpinG1zAh2YCqmrkZwCH8799
amf6mVaZJUGlxwvEmwijB8yOZdOpsrapSQfB/A3TZtffJ0nr7JQ8mXlcTPfypCF6
TiCmorcej19IdiZZy2rM+tzH5je5g18wmw90RsGxzvJ0XXD++EBuulLnimwxKmzr
qMvFw9Ee1jqF7uz2xeAPWiM/+m+P/KUKYtewhNjLm3o5fKMT6H9huyO7E2f843Ce
CTbTe0LmN/B3odhSMBRx+NsqjrVj9rXJvBhJECGfPcSIPnTu/Lbt4MG2ZIZLcLou
YOhkJzjEanoXYHB4JUT9x+EHDMM8TnGjqCW9yhYXXtjeyaMSnHgJhU5wiiSILeFc
MhAmQ/OpgZFFIqXDquKk8UQDx3BJkVwR2zbsjezCfWE7LEynkS3+tpWpFt3pHHXv
NKWNnLwK2wPLbO+6yboeQRdBiM1O0da232pMTwQcvs8TkYkOtUwOb/sMYyrpFLnX
BTbQfXqO/4s/XyfIPcyZj88gZObFRHu6eOjahVkjLQN0RJAg3HKsRQk8vTOZUHfk
NY9fdc3UQFfOZgqFguxYA8uroGggowTiUc2A14OUj95f17fK+JbVHzzeqky63ilI
FKQomxDFWdk4T8TWowOBGn40sIb7r6tPMAWWkiNi5L030TQBNLmuf1A+wgzE8b1P
IzT2bpgN5XV6crYt1YXEkXd7TXX/Ts9LC1Dhc6E+dDDd7vXvkDA1DyO9+W30dZZh
ZLCSLxDsGNxivpxks/YE47bIyXTFdVEVvf+gPl+sO2154ZVkT6nQc/KA9YrXTssq
HlLmg65wyQAuQvScn93ee7SyQAn0mrRaM3KkLR2gdI7s0bqYPB+1fq0qFEg9d7/+
uyFkoxkCLRb0AIGkbnERBp70UrAmaqFcAu3k9XmoGpBVNYeXWIRpQ1ybgJdReAJM
tX5DKAT3IzzCC4lb5pfOGkZgn6K3//hJJiaH2UA7MClTx9XGjDfJQpRSNjLWQshr
PClcViHeXjcMdkoJuas8cY6GRB6XAN3+DBWI9Pw/AEep1N4haUOWv7IAjNLv23O/
F9YCwjox9TZPsJ9W2ORimDcTQiT2zEwvCUCd4jwPxClE6BpOE7Hqz7cCh+URK7c7
ErDVNhnWSOYOTDvqeUFkbXmKV8gXtRnxLB/JuR30bS47xexHKtBBJl7x+UpWlBrM
tKaGVkTUFmwPtyp4zmLs2mAM992KqtFYGhZOCRXt0SAbcUcNqeHOLg5NSTQ9PUIg
V/bQUyT8lFNWLCFsBUFDRjihcCADTROq5iyx8EUoHpS++6CGS+r+WVgyud2S66i6
x3RJu0Mb2o+Xpl/JO4VlODExo2yJv6OC5GtHMG4NxF27J1iUsw6GYmwC1KrKUJEV
hNP+RbpfrlCxNGhrixukOBDtD9xcRuuBLlgfgC/mJwkThYvK8RWARhHr9jBJhGRZ
2WE0VRq7tUP3pHmdVmdeDCX0UmFPIQCuuomiv5yRr9JRtcEBp53RtH1qsRlaSyX2
FFr+2DCsVOWBLc0sLltHp4llgeD2odxbMPCu3rY3/fVS22V20TypiUfodIsfOhdx
joodYv3Y6FgkQIRk0eg7OjNm4OucusylMV+ewvmqNS2s5+PMylrUJnP/ZG75fIxt
ONf+Ry3iWn8oVR9qT/6r+mer5j4C/kqgGqnc3mYEmbvFN2WFxd0Y0/yf/ZB3f6Uw
hez868yIZpv22/zqfCxaZLxjaBLL7NtDdVqnPqJmKbyKLahUjY1yoOqKgQANe58T
wUs5A8NC7SWou+XhpD1+CjuEi9JaBUmP9YkwXtI8AqsUGAmG/9TjSPMb4pbXBg51
bZm/10JFlXPTD1BiSGIC/6eSe06HtXjZvrdClQA1u5LRZwpJzLBMV0bwkwj7uENb
L0UViAEmwcXmB2kZTBlLxIUXGWy6jfIFwULpjXaI5wTHxkDzymeR85qsRCG1VUzF
EVmZ7Xr+taP5IIMfg8HIvM1a0XXuOlA6jvR5bL/e+m9AMQY758et9d2V+0sJz92N
dV5BH7Qs8CxeykzpZNUeDAOBsOgEvFApuKuUHmXRtJYisw6ltkiWUe9iy+exExHb
qdRe2ZHKzXDS/N4mzSrnhjlFysXdXWxrjvuHpPND06PrpJtMkWZE+jlAbYSzL6ej
UfYGKky6vzjzWdHb8gXJC/dYmrAH4TCiF+QHKMhvMtMJyGhJZxK277e2f5mQO5lD
H0g2P327NQluM2LNgDspjq0NlR2iGPM1W2veUZq22jtwYw/rprf3SmUhUyzHjNHM
yV9z4sx2t4ljS/QFxFi6MzyRDySs61nB1W+aGWOkp8hqEpZ6qAn8CEDePcBCnVux
P19FiuZQG21JsQc2RB43MdcyPzZekoM1UkrhS1bdcGFScUdvpideCbEn1zgeSI/0
mzdMKHbZr2DsdxI2ArYZJIxiQeOcY8rmzbi0EQWv29Pe9M/5/Q98vEgc5abXpvHE
GooPo2tslL7fZcUnRpSCJEkYYHOrL74ArvHs4RFxeyjjWRluiThZiN5NsAaNP5xW
vD8RKeVPm/h++AvE4SuI26R6axdA+uoIi9pfXbPLLLQouVizwu1TpaCn0Y0tUcYi
o7jZQ3ghDuhcgtgJlbu/QWoeEcwgOYK+zcK4FrprglZEFulVqS/NDQ+aN5mcSSgt
EgLJtB4KWoGwWl73+pzW6db5lzi6xTms9BzxhBKuuwd5oeH55l/Mt9SD7AQHl7EU
NG82+Da1f2cRvr2C+Rs0s8Mn9stSW81UzeUtyBC7ASiJGwlUR/LQhi15kZdwiXkB
kEULfVu5+ZVBppo9rTrcbkU47eiRBzOROwB/Pgu32dloJjtOn9JHNHeneVSbezdp
vpb0HBX/o59e+Mc4r8wsABCwjVhzemOlikm+yRIrGsWZimL4tVG2THSFJdCbt14z
bVuzz82zzZCzluWSIc9DxrzITJtBzqn+RoUZpOD9Lnz9BGjlMaTr67PMnYjo8ex6
RTi5JTOzVG+Hak3tCm8GMe29o4/0EY+LCgCvMyqGIiVTcyRNQG14bIUg8GZC2r2a
uCCXThPA8+sNC68Zg48ySKdu9T2GdNcRbr0uqLNdmK2UMpO0oZ20203g44S0ehRB
uOcICvukjFnbK+Ni+NWQuuNyiY58jEFVERmJ+rxBNcsmDwG1+WUyr4GCEUlTEqPq
Yyjz5J6Q4ryp4g64EmI95qhFzVe8i6vxjbU4QElP2X6jc3Mydo09YqKWRupIFrdB
XD5z5z5htdrOC0GgEEEcbyvdS378aAc9vpuITtgv+hpjs9bJgm+nmtCkAK+ZmaY5
PqljQ8a3Gte11RVpud0lyWuw3JRjddRPIOIRAtAp9AoGhjlafp0Op4r20L0Sd5vh
vuOa4ApSoZQSCZWDYiy/9WQyOLU7hHGLfaNsOaVllY6pBjP8xqL+nE2FD+l+bdEC
JWGzstKt3O371jcOa7X13DpIrbB1GAYjiFByIbUi1zWJJU/KQ4ko4fJnX2evvx9I
ELKcKcR+GuPzxul1PhoE4ZI2lkzDYlU9knSRZYOw76EeQ+AKz77BMzuYJJewaunI
RBtrsywzgMBkQnWceUfqXrZk+/kwyNrMUU0KfwEKMPl7B1ZpGea8ITb5vpT9sVsZ
Y9eYTHctFP/bTCuk0PeeKsOojMfNrHAxtwOUxaICjZn+O5il1oOaZ+yJFKnBMI9y
bTnLBb+bFtkdtTY2QYV3EGr80b9f10z7tP0fX2vNEtQ8t9M0cVM7qCBf7Jt188UC
/qu0QNJGmkPmup/0s/1ZV8rezq+egVUrLt29KZvsNuj0jWLQrl0Ib18Hr8R1ooho
CQCcrxHlSHrWhuxzvPRPmBFiYyTono19A+kgKJgi/XubFTrVWKbfZaZ9Z3p18eLp
8stYs/cUXXn4fsk9EtPcIhZJrSH6IEOFQlrtvEhBZpZficc5Ak8eO7T1+57Kc3mN
QCknBT2SyNqAClcByoYpCqwtDbIwRPnf+MhMjKvfhuS05KOJ5ck6OIJXPMnZDT2w
7AucyGlPsJsPa4cD7FtkHvXX/0ZAxzPY8n0sb0Cp9Adk3G6vzzZrHtiW762f+MUK
AlTwP/oxZxfQxxuF5/jm2W68iNx+aitD5Mlwd0vfc1Zs4CLFoXUBhRObThj3Y5S0
fjxJLJ2uNPoZmyVO0joezRYx2h+0c5M8gv7xWr15/J+0yVqbv5WwkAHdtkCIokDd
RaPS19YrQdysCXegUaKaTjaD4Bg49h0kOFKvl+eg5KXOTAgIjythFsUj6+4HoF+L
rWkrafh4mIrV7NUsEnSW14Q+Hsntpaq3z+a891RueChB00SBGajxePqnAOjOI5G5
RU2zBLBII3uVWo+8gd9aPZeR+Ojjj+6icEFr64thhuBJuo1Ee+Ymh8K/gzhcWi2l
f5ICv13Ab8uTaUxcbDXHXFvb+JfYq3WvlDZP69sruJdX5g9TqVKvwyvMsQRzhB3+
DnuPh/jxHXYNLZkqOZI88cjcrTUZMefA9+tsKs15jA+/hUUuosDMCdatU8xOKJtq
bz88CUlNr7kJOJC8tSgQx6IQBKd7Ico34X0PKmyVeyHMG6u32r8U9T2rsuTVQthL
Afe2sSLPZpYOffPdwhVMEoj5nbtPRgYPJ+nJe/OjPB/Qeve2CSNWQHFHQXJCi8M7
qBe+qa05hVZoz67hliqILJCckG797M689gZ2kDBZKYUAfZcwsJ3pHPGobWBpG4Cq
Vh/GDmgxI9zY0fyGp2VJmtDatA6YsWxhYLGZDt+6IiqQhbyKfwXnnSnlyTI6rzEK
qKac/gVPVSw9HTQKahMlLdh/KDZ7/0DZmxVA6cookFg5/diz6NqPzYplDF89PinQ
DnVmKaVt1Ome/1xF9Tva07zDOD5Ltb4pPdOxV0COCjM50atc8yPTvnTszbPPevao
ClifEEAf7/v5oChLvhsm11AreNd4RWqMpxxg4UN+kXbhpTMl7dINGO5CgxfUavId
9YQpv4RBZUg3mZWbGcRalbWSS1bgiaFpZTwGgNqHMZmhT5uiub0NsureWE4NyxnI
6MNbswZP5SjGLoBjFLNc1QtDQVSt7YWiWWQ1oVgpLmAo0bUSn93+poZaWspn/emG
/paVn8+EhMvgnj7TPvpeNZ/ajmeQSqqkQGjP37wP06/2FHNEv+P4I04wkBYJyoWZ
uyrQc0Ya+xnLlPUAgx+RAZMGJunG6Q5Y37eLV4kEMVyAaEsMYkq4TMNsA5vwgBYQ
QdVNro03it6IBInS2cxqk6NCsIPHeo0b7wsK0C1YXL3cStCnGNaBvCI5N1fF+wD4
1R5nUAHgwuo64T51vmgGFW7dDLSNTg5OyIf+BGzSfxNJKKxdBBOAk0oORtkmmpWj
O1fFyvPRzaHFzQ3bc5cgEbqKxfewmjqLIIZFnUO/3+8J9zkmi2wZf4JUaxiFxJKa
tnO06GZpE6GUhZakVGvcuuI45aP8Z6Y94E8Ti/vNEt0XeKNsN2SuS3uKkRNAx/jt
mu8IPeiB+0y1urybVnmH6BuiqfWNA9RaIyIwHkgyZyjBXULu3Zi9G59JJUN3hsn/
F7YtnSgr3uiQDw9iTKTRImPXqLLlzWpT0eVQ2VzLyOW+lgpRTvPyscHcpB7Ljf1k
HHtiYh4CHSWUiTff+/lOdZSKTOSHj4eKiqeHuOC0aH5bZxT171PY7wAt2+x4PXDR
X0EUVoS+wrEQYvaQXfPJj8NJ8Re7WBvZHLn4ge9+rzrO1MNYhGde3KQzQ9PSKrLs
PVpohpvOheD91OsCwS4cTgikOsafhlOMP7olb199L5vGTC1wiu/GLjLcMhV8JqDU
QDW72kt8ZAAY4gJa9wC+s0ozMTKIo7FlCmTKfgqwjo41ZVVQFnrEcHBhEG4wNNoY
zaufKw/gewolP8j4ieJ7m0UqH3phnrfVk7OBo8tnN6xejQyiZGMqZNc9bWQGac+U
bIU14fCHZ3526jE9LyJsQHV7Nhdtm6hu9OdoDB03k/qBuguJSzpZO0jcHHB3z45t
b1KOsP7KAgPgDZYwFVzQtzL8aOXnMB1BnCu5KxalB22NewJeqFklTidK56VUmQ80
/hpEEVL4BwbYPxc33H2uqsLVxSch4lP3Mh8V90OMdQdSffg6IPDmD/hImZbc79rc
B+D4nnGLGykyOMx8fULVe6ig1Fo+HXKYFk7FflVpqGPWCHz3JMREpMksRGgk5sHo
+Vgr90tZ9PslWbSQ9TFw31HQKTKO5VCwopNjxtng1QYQKi+0kYBrLeqgvP9ySgMc
cBqXx7klZWAHjJ5Xn6aj7Q9DHBAAAyVb5Tud3b6qDvfoRSrOzOknd1bZZDVvK+3i
Kcbc4wTgLI/1TaaKUD2kweBearebZplN5YQRyXC70gX1ETfnsRMBMJuicQuhm4lx
vDrbjpV3ktNYz24LxOyLQqauZBSYOBrhdFdmViSji/AMV0uycHTAzTGvtOjdXIJQ
BnmKwhGYa1RlwdX5Iuc9+K7QWOYJ5HYS7NlANUeQ9ZieRRDU39yATMpHTsKupLny
wGsZNV1p8oj20P/yF3XCcOYpLz0zf4/TgPcxs+zaxtMCksedwGWjWUKgIhaD4UaX
hdOz7HjUxN79obt4ppqTYbZuKqPucxuaKxCF6MyviahrG6jJOt7NwRwJoKtOR7QR
WOqyOf+/QasTNaCBQeoISb+Wj+DHz5143C+e22U6FwLIce0UT+7JwFYnhbhqjgZB
Bh+UfEFR+vCVGnQPh+8p4CEe0JzAVHfJmo+H1eV61T4yMVEE+9fYICS+QkYlW4pY
gPSC53n/38VWrxm3wbUyv+EjkQwZ4+GQ7k2Bzu5MWtOwlcqmNM9YMaJWRFyqH96z
owSLjwfLsdOdnOsHoCwLaZcxWXip5u0oli8om/9HovalQePUFR2+aDSrWP0QgT52
xFi7DYW/7uHgvyf2DRQeFSka6jpAJ5sNV/198HTjrKf9V2Am7H8oYJWmAoGMpmJT
DnMJmoY33vcnjU43QmNZ9IOgVm8zUnuKSRjxzI1Qps3urqAkIl7rUoa16ZwT1raD
LpcajY3GvHsg0kyr3cz/GEpI1qJZs9caaxaKbgeq6j6zrK8I7h2w2Pil2qSFBNfx
R3tZoS8V4YqR4sB6ReamGoLCyvlKXhsKr4oR9/u5aPW53aF3BdYrP9r7eENPswQP
8DW+YN68zU+DZvpTx4mpy1anFDyKad2xeZaiIB/f7JlkKCXzOZSz0B1T7nzRuzsj
+8Zgj0svp54UL7t2PSVGa72c0Wpz8lWZpi4Brf4WcevHfjalnjHsFu/jPH/815j/
rOhyo4dzxwDPxU3964IkIDfqtrO9ZOu/t3IH5FErKIda8cPlJSqcUjKJ7QG6aFJ2
ArRmWCwhIzM0q893XMc3wr5Hv45zTdWjahDxhUzVziN28UjRh9Y1Mr7RPAdqKnBv
TVnlYjX7zVmY74bM87p1RIQqeT8PAjJBOQOwIX+BcM7T6zEpDmzZHO2I/f95rCk6
AOrSFp7+kZZTFHnH4slvDrwDmygRWkV8g3pw1Nj0bh/noKJB0cQRV5OmyQ9DPajA
55BvhWbPKn4NQBOZnTBCmvMU+K8oaFn9OS+Rojc0rzGgnW8ROq7Ap+d54JxSn7/M
lq77tqd0FVLl/lk8XUDwRrbdfhTSlDVUy9qveUzylbeJhMsaFkRIwnB+/cmHZXNs
1J456XwNtPzU9eLSPctM6pCZw5Uq7ZemOqHuzTMpM62N4VEYtTtcJADEnsLcHYff
3LVHFNSC6K/2Gk3vvoMCu4WambXRyp+0JnMkNxP9Ft9/1LmLJCkXg9+wlTI050h3
rIpxgZWYDhIEIJiopbmBTov5fSAEtXOvl/5PuKwpxP9Pp/zXOAIgKGsHlUsWpVql
iftDE0Nl/wfJhuCydXTMIO6poYSHV9J1oMpkI3qzQF/c7tZa+nkJDKP3JzpfLX36
ojXRyjMhNIbyM80p6dqzta32yTFVjPqLEgdDn6WYErj3u4szAt3o1y0C96vs4WDu
PqDSnFDZivvT82XIpq/MGdmrpaHirVn6kDtWT/EZWKzulmHc9ZgF5DM1sXzqIjqU
RZeEbsaHy74hInfufnHVkChaht/sk6rsmra1a3ozmunJW+dyXwsm5p3Zt6n0bHHr
i/DOlKKn3WLOEoIu5YAvKDgeS9CZ8lZH4sCy5JAGTFckthVkZtMFxinHo8zPWccA
CsQmUWvGk6sFMBTbRYWXrijfqu7MCW6s/moTR+rFoSQuzI1zyQlSkkTSxXF8rq0E
cTJjlgbweusuK3Tkz6ESKG1HTLnZrTDHVAkjC+x9uHYsjjERUeHy8K8IaUOPof9i
SflQcLNSGViN05e2xemH6WqMoM0dLnhw6kaaOQxnQQLZQV767ZEffjIpjX/ztGAM
zOe4AcJmaktQG/vaXWUOa1sNTq0kcHqSRloCexMbslROyjrdkO6q/fC9eJJ/LOnJ
0pPEVOtD7tY6/Jl/4gu9Z9IJI9TRKv2qHXJ9V0goO3HgmA8491n67RMygmyqJ+9L
amG/wqMVa03mTQeqBzK/x1Fq/YYLuPqJxfJrK4EOjDrhK4pXLJCAi+ugwiwFAw5w
0czJjzgMzCUh80Utf6jjcj6OntShYjkDEF/dGyVauhdRzLdIsGyuwmw2HxApF/Qn
DKDsXjm2QyWYxxY40cFy2Gwrld8Ces46j4weFfiC1kBjVaY8DuNZXUupHDrU+EnF
i01YbP7hMiTn59IJVZ2kBiOJ4kou/1DtN8EgC2hfFgQcTl1ksFQOSkaR7P2/Xtv0
7tKk2VJ0qLFoNazjNawXSYN7qYgb9f6fqpKvhIbXeFhvFz9PK+19glxyNPdqohXu
YKTtbXMe3aroApmTMSzPaQkDk/7JVjjwCsZftKnAP44PGemSL45iL0mRNfyb5fOU
ek8y974yudFAyoQ3ALxQYSohMcewQXVHE/BvyMyDn8b88dJYaPPku8Hm6IPqHrX5
mPxVpYbENIp8pNO9wlzPpxCZJuzLT/ZoKWj/6eMvp0vbe3lGD3GnUgEhjnpkhSWm
O9XLAf9Qx886PjHLhYrc17n23bk7ZvtnlgEfHsl3tK14ZJ0YEdiH25vzuzFaNf/p
8u5RC7w0mzXWwFbs8x4qVUCovpIlPhP6gTkxGm56LYNaBcFlossAD8ipIe0x1Wyg
CRoUjMBKuBKVVdvsRazpNZIwgazF81HPnc7AaGbCtkJHeQTP9m0d3QjU9nqV4mLs
GOQ6Ro7VTgtak5vaOzKeoqaoNLVofQ5JJFBDmAKcJmpNNfohRkysFO5U1lbCl8z1
FOmBT7DpaBIq+GkI/AJk40xMnJXmkMy/j0fNnoWuU4677JwFactfhvmLvBNLVLpf
XGE7tjnS9LUvE/Pj1K0jjHIUJrMHh3OJsIqapUoFKTyZ8fTxQGCfhyIPAxoH80Np
jCq6Cqw8zNtEE1GO7jOOLFNrvXNx/IJhnyF0XUulrZB7dSpDCBMiUEMtWwWDLTyj
KVM+nVl1U+cRJPG4GSI5Gw/MHqELoDCIPqKUdqAfOHwd0Q66+eiv/RCpMa+SiIjS
sf6f2gcIdoQ9SfXthuB7Mj/fzRY31C1t2yNPmtQvvlVO/SSR5KEq8c8hV2AkijU3
o1cEuk+j/oHuRrpu00eISbz1iReZq/LhHvlf1P9s5LVEOrjXQphHBe59t8wjWG8z
VoJ5D3TyxkmVtZIfJPe2tBFqooJLON2fq27gAdHTiCDz7I9NRhTP3L4+W9svxPah
AqYLqk1C+NNepsKT5wRwmZVRuxo+DIjP3RLWarElC7xdwSYxDqVjMbo9Sxtm6LKq
ERVRPnpCRkVjhk86WDCpP0JoQvtLOdpBlNX9m6u+LjqD0d/hHoYrhBSlRI/3Bhjo
4FaCU8X1ZnOeKKgzZ5QS9SX+4tPWSj0rUKrqHttfKe1zwnc9Szo2qNMhpo1Uarug
cx+J75WcK5n4BmOgJq0wHCb27GhHP+zuCy5VYORE3qbiyEyimqMBhHhaeg1ZGiy3
Jxojb5YFM/5DVGMM6wlq1DhQbIJ8KanNN1if3EMtj4AgJZQrQESdyQZh05/s2Q97
GgqSHsamE87+m7cVnmXdv0WxtHOc4JyHKVKwlkSuXbPdEObQue+nPLrJLwYfCZgF
t/+Osyb/FI+nIYdgh4Kx6XumeTp1vi+MmzBzg3W4aYZKo3tAL7NOy/+vEpV00VVP
v5Mq68H4wwtNaRtfGAyB5mISJ8vz8mZz4/gDEmOxoII/8Y+UHJgBKOuJr0WZ951t
tWiJY9jpz5VvcxfKV3+Gr9Bg2lQ+Y0vRPiMdBuVNBdFoyw4vVT51mSzcsI/nFPPN
3E2LyX3IvgEiFskKks+XPdER6IjQccoyxPGrN3dSmgwPo/igOEaWE694jftaq53L
MAu4blwrRqX87eesH5aev3l1Ofzy5zsURbf/fKbqIBfD7FwIxCEl9JDBHYkxIWUo
9SI+RYdYMwII45aHbv17Rvz4iQFhHa5NE3GhR1y2/dBDlSp4srRxdhX9Qlm0g9oI
tUiEtTCr2x6f3NJ+Dy8bh/PvqpX3fRqkHc4XIfapD8VoDrJduIjBPYGSEIlxnkeV
EjFtQXRG817XpMiT6oD8p3lJAESR8tcyhoHyCEpJZaFxawSllFaY+GlRR9A2HcdO
PIpf+Vhm0xkr4fvKHMlOkVCIGIY/C5bq2XFZ+IF74npKsObj1KDrcG1VZePjlFci
xYFzw2q4ExOzihOUPKcawMiPwu5tzbG7GokoiyfGKVu2W4kaYcT8jJkR4pw9A3Xb
XDFzgEeNQSONxr0q7ttHh5N/VFsaxmxdmSlV6xZ1BbzfWrkjn7//k3R7LFES+R7R
t85DNh9soJhDhzqwIw8/excorGuug9S7Q4p8jKBUAAF2JGBPA0BXX4JCt+6lyb8w
NMYumg24QdVyQsWgIG5xFEjL5HsgdxFBuomb+XUFEWR84mbj1cEL76x0oVvOzev0
E9ttcrZbV/Im4WrXOlAwzFPrKdDFNU3YzSxbqa4Yh12bfk4VeNaBqwP6r7Z4AZ9a
uYNukQbRxBDF2FRY2MDrV5kpDO/yGg+fdySZ7RKn8UXyvg4fqJYL8tJbVFjlcrP/
n5i815N72BQ0Xa+cQE355jX9xk2cRDKl46RfQJHi8B5GU4aRHFymVMBr0VK+n7Z4
tmdbZ81LblhUoXoCO66HhoDglhTvqX25Bxv38dNyCeEYB2zaR4FARUj57l7yEGhu
Bp/pdqYQLCneKxfZE+Z5zUne9l6YyFcUG+Hsi3xtKfRr4aSmLSR6m1RAVwhtQw1r
7w4Vp7Nap1lqDpDliMSCJz65yw5WZ3p71J7oJHrQ10LJv7adRX6kfBY8HRAamhKo
DlHJDF+rfUuNE7ksvN0o5gwQp2z1HlhejalbAhRSUC17g/ZeuNYjAkKiipqH+zwC
dXo2PRYejDWBfK6Ty16NoBmuHaKYCXsj+G4YpkKBaRJDbQHvFVVpmL0zLUhP0lea
AfelHO9QI9YyuJbUZdfJ6wBNwaPJRYMvjOloHD9JtvxSq2u2X5UwO2f202CfXCn5
5DxWcdph0uRE56j1uswy80ogrWthiKjwUNGO/SVXBaajw8KZ06JN4BRLso9eBppm
9Hp8EJ+A3TInoi+bFqmY/SYEZSXeAZzS54y6ZvqfvxkDBkU1Y5o3SjFPeKhqbB5u
jDuPBqJbSIHqkutBpK9bg93XUFPJ0f0QC+4J+yQayjA9jEeZwAco+oT9pUaBAN8A
hIhfnUVP4CT7peiMGy9N5FkOamk8izDPHzQuDZDYpECih8E7AbHLcf+zUPeG2mcv
PwwSUfnE7T3uP830/7/+jk31TBLbQlF+2wZns14tPRaTmj/Nqtc2dAouBOe7riFO
gaU7yop5nU00CUluGVgQ4ImC/+JYyOz/1hIuCQ8vExr7hoMqNA2H29xQvykbRMjj
wTv9Q+9cG+UTxb0H5KWJ7FTkpBDQYEczs4f30tgxNBFzxnOMr8fLAXlO3SODrV0h
ehxUVZPba5m+MoaZ9TvFOKNKBQ+fheWNJ35hjM/xJ1xVFOFsS/b/OZQr2Ql+lmUN
CmOPGRLC76zfgEjKU+21CzXHaEutB8klnHlO2rANOvp62DE4GOAbqioOR5ErEQvx
RrRH9DIS4cIu9Qa0nVGjsUZpwMCRhyxNJeUMDMH+w6GHBzKbN/zVFNPhSJkCFAzx
+1hfq+aDGLM1boAc4uqZK+PdZhB074XSlxOrCLfAjMpiAIpMwqBc5FLCH8efDwVV
nVxMV0DTqYi2UFSjbbB9WR+4+Bcg0znXwb0HyJeIrDLMoeYOUOk9PF9xRprBe+Fm
A/XerjRLrCFyMJFeW6ksWzFKMeukw5eYVYO8nThIxdZgAVyeKuuDIQlcRYvr7+/C
a/ryT7XTiAjwe//ZcQyUa4JZF1lb38kn3GJTfTVSq+zq4xi5Ybc1uUSmRQC1oxaV
NyRzLLVVqlgc4V1ExPHwoizHXrCegSUoAJ7CEiKTyHMt7BYcQZRYLGYtfvmg7RKP
M+yFRVGdjwEnJXvdj4B/BK7n7pMVNSDzD5ROahq9ecvWD5jDUNXbxkLiAxy1SoVI
3OwT1uaXWLlibDaKpkfeGfKFaEyfMXeiv9lkFyKChYIGeHj62l9sMz2cSQI3wDjV
JzkoHH1TbX+Xhusp58GndC3MTpa3qcP4jpKzXpTLkJtlJcocT8CiHBMV+4ks7w+Z
iJZ3rXRlB3WJJtvBczL8DLv+XQFGgO3nPB7zm75uRkG4Hic3LWj4HYyI/CSyDUAK
/pw4/+a+ANjbTuISO2dqlhiu7oLo1LTvO1DHL4yZecDLU3CuKDcB/r4nhh8XoCeQ
vOknYywGoMQAifhug1vNrB9z2LANHQqqWf+8DvnSDirs7vhx1RFk+MfAX0kmekYb
xgLS2+rpTcf7+JY1SDhYH8kxCWDuZQAluIouduKqFnbGI0fBqkvN4tC16TqXDioK
aqMLUEAT4YClsCLzecl6vtrbbHMiYTqLzY6P8P9qWZc+OB8vRU0V4I4yPKBTdFET
3g/xi2lSaHgKC3Ql4pDPqkp8KoIZL+1o3tyrP+5SPuVu7nqUFpy8h/OuheMnSkX9
ohkOUnGWK05E9nhNP3BTvJ68I+P/9+ND7EnN7u+nMgln0Nt8zND+gqnldb8MWf1T
BcNGtbdbTh+7QoujsFW3RI7A3Ej/H600uV0RcRD1qK8F6/aRZKqQLkGwEHpasYEK
wGxm48SLuvxw0GdxMnYPGqUp0CukyqVm/EbcTWdmu27dO1tOPlIotqd2i2mospcu
lBKyIz35os5rDFXrIcNn2KFUzcE/jn7XMh+9mkyroMz8wkm2RAgim8qX5bc7T6yE
HXToHGc1VlTh5KuvtMlNx8hDkeN5f8FCUEfpryWYltn9jaUllA2FKo7VPK4x19x5
tEcSAIOq3y6q91RgKJ54CkavgLDTbY4BcSJ3ImJWP3mYvmF30tSC0ApAShrt74NW
kjHyLQG1VTus1x9jdDIKPh/0I6dqIDimQwpOLfG6tpVu4/9KB1mSkQkAtkSF7Xra
qy0ILtk1pkEsrpWgL4tuMQ1dfe5C0dPYxTqZaSKi8mXs5EVFcrwltRAFYP4g3DJ8
/dBcAY56JIGlUkkuMEwg17gzZHjDXPSO1so5GPxEnmG/ii2PkDFzyvR3oVG+Tbt9
H60hJz825gVXLiJiU+fe61F5t0XiLmTdroQEg4xLBfxeJl72cRb3nWtZIiYlkgHd
7o5sgqZfsQNQhrTM9ph5JYOwc0Uvq5QvFjBR4R4RJX2WwGwfIIDuzi3frqk4f67x
SraENF1eYCSSLQ4MAhgWQ4uhhHOn3ivB3DkIGwrPQRM+uc91qUr0eK5M+dbN0Hm3
X0axM2ZGwxD9rv2qrN4lpqpFjAxTKZQWxqdl2SVnNe4ckQ6V9omvpca/iMmW/7bI
m3r0kJT0SKr8Ls6mRjltq9d8PgC3Hej8sGi22swXsGBNkviLWDEMXs6yQn5cBFM0
HoEiPWGwXB1xDuVmsJxbR6bPFLK8+o5fVfdP5PkWogAg9bVbfxW7rzJZLqLFBpYg
FIMpt9B0mVrido6KnYQR1CxgTBVMhkHlhxNtBeix7mhT2gJ6xbt/UX4rqzDkxCjT
i2NvjHz3p+fOKMtOHFnERGHwEcRTrY//wG2xLgNruLHdibyNvQzZOx8CnNRUsG+E
kWbuEqomKyYbSoD1HfBoWr1G8BdkF+oMJFTo62FC+m9tT4y/9aI5i2EjvWMRttVV
JigathFN2+XUvEaGOJwMg9cjdsU5wjhvdUbtkXV+YiJhCL3U97O+I4rss5o7wH6A
kSfMmWCMrIwdVotF1HViBfA5raXUvyvO3J8AhWYQWW8tgUTtlQ+PJ9G32gOMcSFz
d5ZqmNnMsxzFZ1Yj5I+EzAzeGDZCQSayK/5w9PvqhLJYgtRl/PnE2AqOcfLKxXV8
b6galh6OWaiYaYoPGNoZ+pe3dica24tcSypQuOvsiWoTeaCP7HUf4w51rM06MqUO
OG8JcADqA1+IZ4m8wGfUQygCK/RBnYwVQ4ZI7QFBQfhECiPFIJgaCr0aJ/v0nAb/
VtcE7AL7TJ1/OOn7awAncYSBHA41j0ETmQY5K4vG1VmjHjoSPctUQf0xwzBLaBMJ
/xNB8Q74Dz8TyzP/WwnunwOKUGqyuaYqMvP6FD3NnTl9oTeBUJ4fWUYNbss7L0c+
U6VFuvx8LlUhIaXMogby6XH7OkQrEE1VYmgOtRIx4OMxTOiCAA8il9DaMufraNeF
3pG6HT3S80m9uhi+POqOz+ScPn7H4TCwozr8Zuqm9wC83hQtwML02HTjhaCyUiQs
rwxMhubqkzWKnGM3bMY+zbP//fK3K46SCvnYRD9/lS7KwSnGDJsr/EgXEN1551JD
rIpiSjpzXDhQnrgMWnIFSWo03InB9lbLkhIAw7YDN8CB0YPQymg7noO2J8xkrCUm
MHBzhcUTwYR/phRb8Ox/XwKBn+c6VMcK9ZJnbb/mfIH5ojvwm0UZdsi6nZz86EPJ
Yi2p05/4xknfWcrVbCLnP1fWRhLJ7HOxnVpjrhTzHU8hRbt+zmNCKW61rNqaoDFB
610oH33PgYa1Iog+7iom5LZ5VQeTcorBI9JoxcgL5SNxDIUS9n17G52pkqz3R5Wg
EZmkqxTqLgSFX0Ch2lVEwrnYgDFCE/cGak937Y9h/Xd79aDysFprQQAD2LStPHKa
e6dZIa2a3zEhnXqiB5EYYaPLuH5roRlhOSyM3oOq4mIAqPmUf3zRoz/vjmL2UfuO
QfCqLEHj3qXM+x3+l2OwFz7txZMMNqoc5l46nPKy4tlkgyGAowM9aBJ1m05gIdOn
IB57ITBj0vdXEerY6mvBTEM9JKebFxCuNnAOkkSNteZ7t+2lx2UhFwW8ATah4BUT
j3v6RTVWSIADoHjB6edNekMBPwtg2Syxa9sNclLjN5RxfUqjTrSfQPlwMjJ1ulbv
qL7Az5sElA/qvCt9q3tZs2Bv0Wg83yak2YzqOQGLx5gU62KqP1w8yCuYLrY22YOj
Di50QdQaR5k0fTu1RIcVm/Mo9dNGp4diqLw+qoikHEPj7Nl6Gzklqi8VndGj8mfL
AIa/654lUXez2kSlJ8g45lqrWnALZXouWY41QfRujxNJ8tIqZcuq4tRM2JXZK2ka
216dLsSfpl/XvY1C9EM3hJWpawjDQ1QGsEKpv7Oic5A8GuwgA/cub7kUD3ZcU2Qn
Cqqs47pMYagz5chsjptLT+GC5QkbZpQRXk32xtfkr+iSPmFuRy+dMNuBeHwchEJK
STiOoQFEwTuCQ+rfQ+btE/t0jjj6sDvKRXrQMM/KDf2KvV5lefOY30Av9AiIdxAE
5Agy8lvpRDwbMhc8N2L3G/Q5sC7W7oYEQyHfxobFrkL9Pj84NUBcKS6HMZXb5Gv4
+2e0Os4BEwyD9dJ8o8fT7vMZcmIZFxTj0QDS8PxEzD7LMnOYBrgBDuhVtDsGbORv
Faqgk58WDwihFbyq1K5jEHi2097tND8fF3TuO13kRPc8DnwFHflO3uqxOAf12P+S
xuh3H1P9Zi7SH6b25X5r6IxUIjeUbaMw95k3kH7Oy5kCURTM2Ybj9Pl7hCeZVxuB
AFZ+JZA3RctVY+jgI7KD8Qqa/4Xb7TvfUX94cERDC9RSp6p/0tK/+Qp2QgqCL9Ho
We7/z20sgWLl8p+OyYQG7oWLhvJDYtCJXR7aRZ9MnlCvIhKa/3nkbrm/v6CmovXC
HuyKxzIUpGIEzS09RvdJpUf5qy4JB2l2gQ0DutqAPOlAC8aseZfnxvRhG1FDxoBk
X0isSNp4VF0gNMYddeZxYpuWUJN+w8xy+B6tr6JHmzJflQwYGX4IhmlKpSg3VW3T
k9kN4Q+xzkDqzMbF2xXIYnY1Ijmx3pRTPiOFeyD2QUNcsVC/YNAzK94KS1oZNJZO
+lrBzHpDMRnzEdjB0Oexj5unQY5PuStgm5sT4Z4j9W8p/NLOiycK0JVuak+4NJ2f
2gDS/XbFgOgLqxFsK/F2eS1sdiuVy/9aId6+JRJnbEW8ImExwMgx8XfKFuq/800B
NmjeV3788fvE+/rc1xvI41GFzWRITADvfBiuzHtaN1uvQzXW9h3ZuS2KzS3/4nz8
CUSIqo6B6syFYC4qY9cKKMkQgc4j7htsY13Yn5Uq5kO7d9neeKyE+6MAchwKIBTN
3g2pWHDc3Ma+Zk9eWPsQ8u8CdKV1JJ2fJkr7ez1pKpatQUoleaI6fK3ZXu+v6Vf2
Q/ZjrBH05YikyTrRfhkoY81EBcP+28zM+6bDa4n/qQKma2Tf9/TMiB+Zds9Zligs
GlOxRCECIR7kP2+N9ZbvAlc9rMiQvaEOnBtUYZXB3uZDc2Ge/B+1LEgq3LdCToER
/jyXEUNr/ypSow1hm7uPRRICEO9CwkgmVv/NYV5AUZlv26jvgXlLGp4l9DnwlAtC
8HIMtPbzMPHEoGccudFsdIT3zgUBsWsM50iigHenX5VODscPvyr2c7Q9b+8WLgci
IS0B/zxZWtPUOcL+av14BVuxZ5tPqiw3i1bfJ22q/i9CV/mKZNDsTPyBvMImzPP6
Lg1RNoVR8vko2ksGujJTtwa3r1dbrMAyPn+6xmRXxOTzsTPqCVXGmtgvqz2qWAn0
2in1V74+dRud8qbLJTCjcTo3mTsf5DANBI+C36N30vExWVakhyLorNii4SEFTItZ
LOPAPzHvUK+yTH2IgAbvg6Rm87h+PgicXbHXCnDABmuLAOxlnkL3RIWKpIzkpeDC
9pU04Y/XugtRsfKkSWFxCZPJDS9nZzQ5g70K0WOBBP4V3eojMGb45bAAVSeUWwBU
4HrpbRL7uAJF7nF2glnAfHQ0uojCfaZRE7ZbsQH9HTfg3eRr8nhEX4hQlHQPWNk0
5gVjkaLAoxoaEizhNooFcPg+HRsXhdHH60HsbcYJQzfmBnwqhP3Zd+EwPJ99viXL
8wYdIHxbqWXzg8MDjyOZRNgSkJF6rTKWVYtP4Ih4ZXqmrb4RFGJhwC6hPeWclZMB
5BwjmYUdOevRieWr2eQa2Kb1cP6zp//2+tcd/t3V2I/LqnHOZKSGTkPnDMa0xgn5
ZB+zbwsnQv8gU3/v2Y8jzcYu/c3wmx3AVWqjh5lhjBtHvZPDbfxSChOAlCpdEwLj
ptr4MQB1YKDoj8trgiBQxsJO75lrG2LTs9hYOk7Hd0booangNaVuFJGJqKPz5ajH
KY1dBNcjV/S+kHslP0Q7yfmDEjpdoJpxqBlkr3n0gqTB5wvGIraOPGqQGyK0oDeM
R3DRzKcfY1RNhLldNS8tNm0E6oOMv8bhdhE9TLia/MMsBAhhk/gTu68dP/iUPcup
iqo921hVtz2vJrUyeL/A8TPJ4F2pvpFK3Z/zCDGg9EYpI/ny3ODsuiN664aDE7jL
k2pW+fa8yalZb5F4DX/8KbZUlzoXlrC2156vDcqODBZnozpzHEJPLIXXUlla8Zl7
wPBiUEGDJphvYN/IBSWJvgOKdOSrogdlf9OpVHei5OaEUDXsW5g0W+8rGTCQeA6p
1J1WLlqqowuDc+uLwMIZgJaAGFb/EzLJ714aAp8Pg2ot5BMPLeWYbUROesaIRiJw
bHx5/QLJ/O1VeZHtyjhLzHupyAiNE7O1wGlVErd8lg0N/wA378fpRRxH6pkhhvWK
ZBGzWsMiKplc3cCE06dBYLzXPH6VSz/IEIO0cS3VtYSZithMGGYj1bmBA7DnnCcR
9EGyQBtQByWyW0PDzun04xf3mvLiTYf4FD7dhQrjL7xmh/K7KlN4CGba+T4y7clT
GG9YHYYHSUI7h1D7wLncxuzDY98XbbR6UhlXh+IPZ+rJoo8xdO9Et/3bUGG4WbYI
zeeLXVwxwpK6b00KDTylecGZWo2fhp6pZPQ2he8hopyiE83fe+EFqOGMG5gv0yvt
vgne5k/ZWpMfEii7TaJLjS34wlPkhGDMymXgUoJYFdpoGqU9LEhuWCYCW7C36/mL
JdEHluPoCRbB6M8Ogm9BkYST3td9ksF9ZR1bbrexqmXtTKqLqSzp/z8F6QbG/vqD
TQKa/+KG6JuHCtfplF+6yIUQWQNQbiY2UckEf3FnKwbUNyGAQjWxdfdgvsc89YL0
9nwNXX6Xy8iCeZAiUKFbzxGzxZVQ9uEm8NikvySeymsKYBYwmbOhgMKrt5iHKjsN
3f/hUlsdx3aDr8SQHwFVbX2M+sjhSlP+mSGFmzbOkcMLp2SpHig64mWxHM3SoUL+
8AcgtEPJQBQIEf3qr9YZeUCVbCQATDhASqTu6cD36b63LD00OqAt8So0Ahk/32Fo
oR5VyolckQnSlQTMd3z/0T+LHv0XLCbaQzI6uIeGbF4sOGIDs9kD3z7e3pMr1EDJ
ZOYyyuiGKPwrXEvdRorlZZudDqhg5Fv73GRcd6dVhrluvXDPeLecmq5wm4A4opdt
yoJq1DLeRCd1C3lr4iUi43eYRID+AJuAvI/zFQ2hhwgWIlz++hCMajVkB/5LkNIm
mmJPDqeLF0TIPpEgsmfg/PIMxe5+WkHD5MOwBJGCuGNqRBLU/dAoUu9D3tgIX5+e
u3iWtJZrZe8WrNiSwsjZBicP3uNz0dytnBiHjdksZqRM5YLgcCeXTJFD8gF95/vu
zpyHAmDSF+fSb4kv+/JXCBXhqRi9EhkxL0E4Obmy8Kiaw4kxjGjwu1+XCnDecEBM
XhLRiyK4H3Hln5ZWGUyQ/xAe8Vm43EfDPezufKBOYz9nAvx9OTPSgM01I3EDTUbt
+pb1yghbCsw2MWYqY1n55iLf5tyvFPqV0Cd8nPLx4WDfcp/1IEztLEziRAtqV7wH
bcKG9SbmCd3Gc73MbV81y5wBcuSW4Fs3FXMib3QLB4KKV3d0kPbQUyDJF4IvhA6U
0txM14Nhycx6BKCsk9xCVRVpuA7HVtZIk3Zh8iRt2m+lSA7986iaZwV4BgPxPNE4
soXxSTd4wfJhNcT1KeZ/+m8fZzQ0WHdC5c5wRGI/KIKFhoYenimVcdczNgsNs/9v
gTXCZZY+LMdBW7x7VPkHlxV596HsZm58rcfknGoZZGEFzg3H5ZZt21O8tTj52dHl
noB3rhQEr3EO5J9wuhuE7fu6lPE5WMz0DUlCD6R9HmMMjxM02kow0G026QKG/q51
Uw41vIr/qFVitKdMSCe25HfyaJ4eQEmtL8xND8d5q3xK8FGpA9ti+M6Thh1HS42h
bsk8ApuJ71K/V01coDRzpVQKtSqG3pCVhGkTijJVOM4vnHLJwPqp9qARwEoKzT9u
NsCupKl7DBRdGRSJnlJlXonR5Lv0QDRibty644niqZUF84TIanrc/ZHjQ4t+fDmd
9FaZXsVB8lKWH4d/yIXlN1Mkb/qj6mN56JE+9DOtihynXiyuPiCSKkQJUL3SiDA8
SkYubPz5I3S3gfvpaRRNvnd1o0LfycmZFfWzdprhGMk2Iz1Wlh5KScE058bvjXff
k403Ijwjj1APzhC1A/J72iNRZ3RZ0IK3H4gNgsbloaGG+e0yEm95Ffmh+NMOtj0n
hTmPvwJMx/qXV0f+daZk/gRZgpfVlnkscOQiRyFhgiogH1pbUwgy5f4loSqQVvyT
gmaNVwsXivbi4u/b01DNYcewhAyYy8H6jeqSENz4VJ6HFH8KHrT0PO0yLRZz0utW
AfkiATFjMvtg3drAhq22qFQZQxXFbqm0uGGiyNapA7l1VAZLodHkYrLTisTFig1N
IC/Ca+P0+JzhP+Ni11cuF7bm1Isa89GNLKcJWe5xqYbuR6JeF89as4xLOnd9YEND
H5RS56WD3wlBBU9luwK2Bs/gBZpCVfFUGv0d58uNyzJxFwAAVieWavPWbtSHMu7v
P316UMM7hrkDj7+hhKuGehU7ayzeF/9j5KINnC4WkomcC5II1WU85XYmJJaCyaBC
dtq+qB1kdSKEkpfws3yP2HUHbfL6NA7FtgRsVjnRXYVfkalmgjrOevC3moLgLTDU
flRErHRtBMqyzWrV3z7gjaEOSutDTyhNiDs8t0I4a0UAXsPJmIE4EEJEhfl85luG
XIaOM834oHqRA2SGgqdZ0zKzNHQdOv13RRWc4xPoB8bZ2IGDlSHHrTKe2wF587ZQ
r5J1Pf351b1TzerCAUSwQ6V1487GWnLYcYKWCmmtuQ51bG7ihKwkRharTSp9J9Cg
BJwy5Z9uk2DBSGvet9oxKH01Valat2IjyIlK6VFNBj8iv1+MeYeXv7djV+g4liSO
pjW1OQi/Vj1v+HVrqYLgiJvcLVM6Gk6sIWBm3k7g9ahAXCyh2UBFlo0Nzyd5WvPL
GKBGbvaY9IYSEAfTXygVrgJDDn8jff11zct/Q8zE8LWzzxjHMNH52GKbyzUz5/fb
JxKSf3qsr6Kc5BWhIyM1JMg0sSlx4xhC0FQp0F2QDmI6miPf3cpTXnI0XC4EgZTm
ko5w5GW1aIsI13Jw+NsMbH143NlPMvhP4KKxlllwBLx+ti9+FRmtXlSKZoe3DEXt
yqabc6dncdwNAWoNBvpxeyRc77KH/+1/njKiRQNJSmIqDDdbXavkUKekHD5tRoT1
wM4SEKrrQMhr4qOlJckIBHNztf8GDCMJP+LNbjr0IUbn1HW6pRo37VuX+7Ibd/8d
ckjuyb+RvOQgpjJz2MNb5xm8Q7wqUs8mgf8J8qrwMbjA4uPF4UBThe9S3+NobAlc
/c67zbO0h6J8ssLf9ay808GZzwc2qvmodWOSDaMmxmoOpSlWHtg9MLlrvugjMQKS
HYy+d6LvE4TLcvqOf7syuG/auUB3hTRzJRhyzidTbV8c/Sb/gGF0KYoI+0KqQ1Uk
TJpoWJ/9+0xHEvh7ZqKJlkp8f9WLI6cdMQ9IO1POURU0xyEDmUTB8E7LlK4iVEby
2f3/nnmdOz1HVixy+kQG4tfelvM8H/6kk40F86R6DVJa2ns0BqUQ5YEltLIycR4o
KzL/V3WezPOzqX0EKhWib60/eSPIJo1zFORNFMf6vg3NPzf/J0acH1d0FJBciqUA
DjH/ZCc/z+QjX89JUrWr6JiwjL87T+vYfdmyB0TwZU4pqfV385ziMq9IyNkM9XOL
hEf9azIxiqsWVW8IMjGBmuuVmIL0T5h7KJUM5Mm2PsPdA+Vau74B8qnDB02EoKga
eZbqd+2Wp3S22waW2KbZVb/LXqjNeHN5ARodExCs2a/TbBf3MLURm0xblcIOmgHE
oP8+fpSGOUabRC3XOYNxno53AzPbG1PJHyEqpskenOJuaejqvBZIYolWTi0Nn6Mw
cjSh1REZitpju4XXu80c3Is66dQcQbQA82JSmEspnRYLMO71ARf3QcERFp8+TR1p
kw6XbImYbdwxrRVzHPo0mU8Y4nBgSIeDjqSXBgUlc7qgvBncdWlrhgOhrlSvtktS
ZuYCgzP/F5qzRe5sqGJRsE1v0HI1JSWHxnjkmVLLjjKuOSpeFhWtDOxsMeknyiGl
O2UKIFeFPFky4bkGBYDjU0zdhgP7jRL5AlzMkKLjPXRm3FU3I0iDP1efLffKcwiw
26wjt/Nzeov4DBBlFYsa0pLXwiyAqFqtGYiqkn4VJpxnLBChwkgfqdHXTrbXPFsn
AwVpqnJh77ecQq6fl5zS8prymQuwFcX6aAR2ETb5K6WMFH/08iAJkYW9DpjTyOPX
TJ6p9jrlxq9+B76cUWpklYaUZle3eNLAuGbS/yxwd7tMW7LbldLEiTftcAkLCvY6
eBNkOfiSIlEE+0j5yxeGC+LhNQ/DwUDFIjb++MS/9ux7Zzs2ldyh39dfNltaiy3F
EtP3PMORCUTzrKX5UJRy3/ZZhwj4/wEtmy0b6ooav1H+CqG9ZTjMHGMb9J5fTUlI
aRfptKUHrgL9j7CJggVMdccULoDQ6B8FtK3C/q/I8p2j+hsCE0QL79MPXvjopK9K
YDOQkOJ28O2XSQMMRX9O4OAQ8lrqBdL0/rtKeLjwyy4TItKXhL/gGHnRNb9HuxnH
3cWO7T8SCqEnAPoObuXRzldw9xE4nakw6WHgGRoMfqZd2nZ02UsQEtdXAMD1PAVR
Lp8JH36Pr/8bhwC+2VB/5rea5hl3l9EfOmec4opeECp5NMCIHq27xNqpV0suyVDX
NJqHOMfbbvQRMtiH154HJtaj5erYzU9V/junk/I2+tCY+Bv2aV6mY2/HZs0nu5nV
1wkSzA64BQ0IjXZuds6dP5jrqUin1e/hRBehG8H3agmumjUYp8oTMr91JSITW2Jo
cTj/uAs6xi1dNKaW7EjPlNmr6JcEivaUepnNaQr1oY+UFuDjz1Mrrj4S2BCQgN/j
zFsHSQcB7Ip2s0au+GoQLX5JxOv3Y6bQMe0IYLX9cVkuR7YXTID3OKgcP4uTW9Yn
eAvYTP7oMdEMJeGuIFLQgoffSX4QpgITLapHcvYBavQhMDbeEGyT9+wkQgRP5qcs
jEL4KXO8i3wW+BiA9pMfF6/2IAZa59ErOOPYZW7keirUAAw2Ikmo9pyFeZmSe8j7
VxqZhoXeb1JcvxGViPArIBEydpFnEuVWUFPSOsYhVZTWZL5cP/8TuME1LpMqgwhu
GxCpYzNIbDhLDg0nNGL5UQWztMDAd5iIyLUdM7of4NHoiYZfn26U4ucjlNsJEnK3
p8sJco/McqYEmrPBrKKNszzctMP+rvoFUs4GThvboKe7WQGnjlll4ynhEd2rHS80
ni9DkfOtVGABQ3ylxlXSQTPyDPTzUTPayAKH1D1aYywbASmUac/RvVnlqFTmy7Kh
LxFFiucmFdpCOfEzk/6jRNSehzQtEam6I3fmqAnZ+UqNPlu5Q/yOLNFmqmwe/z+G
9s5SA9gbsliEF/5/daXMGFgqq9g0bZbbHuL6gPIyOTPPHKKQ1njD10EO/rt1Hutw
T1b9lOsWMzGZt5T35ISE1lnEj5izFMGavs6L4QNiCuPFvQ32c5PXjFNvuQfyyCn9
RNWKEBoWQgAC49qSTPf6Zqu81Ne7rohXGZMWwcAiLO2db0XB3M6hExn43GjvgPtm
K2E94d5cyURC1gXtH0P0NCXVuPGvzkStMf7j28kTZSP5Cxdtu2Ni1ZNByXThihr7
DRAO8jQ/R95s4AgUD+lm2fS/xnX5rpAeCRtsC3mECA2UKBO4CsG4FiBr5quTalSL
+xhLnFpmDWimcOnPi1vId4aIPpkwwtE1h+gSW8w4WNe5Rl3wCgB5wcmcI3KKg2UD
y118i8sZUOQwdRzA2C0Oc1L0Gg1B4NHQ/yZ+FXgeK3eVnLv4yC3h29YVou4gtuPD
N0guR4e9uGI8z1FOJ6rFaL7HOKvrFrwb5HLliiMINnk58c2x41bhmfszorgrHPvb
Iv3wOJipk5Lxq8DlPvIBVzBQkczuKRAuUPVtZI7jFseNfJWnrnkVJ6A6WFLvwqCN
/aS6BamM0MnHzf2cmYGFcx0FzTNlmvxAGPpQmLxBddKkI4LfaUJD9DK5Pz1PO+/j
svk6SrJ081nlzkm4bC5xkFrR3mJksBER+3BObtVsjcdJs3AiFC30WcUa9gZX0KP4
xQw/toONtAflrhvg8DFl6XegensZmlTgUeCbeJUzZ/faWTh0NBwAdzr5d7NdofjS
K7x3HyMGN8coQHK14YZSgHyTlZRE5s8FrEPU25QcHpEIkf2eRHffA5s+GpQEsvsJ
/49od+cHF6cCElO/PwO50jpWUfog6vaFP8wxpZfyDS6/H2hgJKpxRgmcEZs95DR0
1gjdg4HC+PU5uN0RNgyRp76LzxFnHFQrAdR1DzITnP5Oze/DzYC1xLY57S+DmgQA
VZ0qgc1oGcrhLTZFPtKoKzIQmttsyxQ6c9YV2NiTT0jTLA7bvtP+LjJmlc0l6uh9
Nq6THqsM8r8MmduF2N8Yz4h2dMGo4+U3lyiEU+1lKCjiTRfsB0xlbpi0R4IRbvXy
VXotMWCRy8Tp8+VNKHp5GG2LtG3T6N+utKSCF0FahEkAecccjdVzDv+/j7Z+Rq0l
eL/cvWGuXi41lTrbBcxVxRVFXRVDnGHCyYNxW/TUkrMhaZY9GqI/hEFerkBa8EQY
9kF944ojChiH4+723Gy4wGPe0yH4bnXl0lzwAm7yMuf5TPbkvyuIZL3F9jkTfZof
+OOLI+cmTl/NBImsJyS2QRQv6Xn0v9gmfhYhvSWeTTkI7+wzu62Rie5b0upX8OoE
TsBauhzgEb47k/17inIG/lS41lr55itc+//sQFzKKbSmqz1PJ9xvWbC8yiMTMq29
yM6jvi/DybUOD0DfQ8yqIQyTQPpvtR/zQdXxgSbRkTpjRWV1LI2QkU5+wCTpnVrg
44iTvaWo/3icqHIETOjrH5Q5y4C1MA1PmBLIDMF69ZlH0U7ry3bCG9//DOdE3kEb
C2LVFSE/PTXjRxjvXIpGrpxJ1DegOvLuP5njzqiu74JiikXMTXIiZZAFV9uw+RLn
bnJxVOVnUn4R2UD5uwdRULrE3apSbcqS2KwP98A/zpebRNBF8KRfSXmbnZPcNB6c
JyuaVzZSifLel/hp5dDuFNsQWSpF/aB5jrOMYFE1GiRahVltOUhzTiIoBKPPiIAw
r17+f9mrh5237Bh49tJvRV0w1FGR2Ac5UFHfAW8hVJXUHODRzFKCZtxnjJEtBdKw
kJyzMLA+pwg7j02yDy0f9x1xSMCpIpKI/mLnKkYbruyEn7498b67+DGqBL4ZqS4U
X0DUX5tvRhQz0iukNZyRtKs+DxPCOOuo2nfQ3rRyYyrwZ1KVYlAreGkdJ+DIXebo
Ow76HG714oqfbxDdFo8Psu1dW+ySTlm4psonnNzxms+fDu9cV0Fda2NfLv+h7vVw
7J3GHXRm8eP8qARwq5eko6th4yZnD3KuinKOXbnL/X25x45RvVBDCUmapPxNQoiF
njb7hjitDRKAX4JA2HZeBj2b1r+6VbHx4smK+sTb0r0oR+ngONBrOExzGYjvZsdB
V/X3JAuyxa9FCmOoxLn6g25Xgs1Nnr+Ccw6K5vJF9kWOfJC2Og9WkDcHOb2940rN
wxhhVS7RGGS5yagxNvxwA4P2DpGiJJTd6zkpFfllSkFKWeBp3aFsyaR0AG+XP/An
YNoZM6D5GViS8yedJS7Qu4wLCyKQxS52CARdoEw53/E0/MSNLVjUZAwTOZeGn2t5
1HdC8QPNw8+ysNKibwguXbX3X2lY9VD1oeH1Mz+oD+f8jNnODS0CNx6dTcokQtK0
F9WELAZgcc9gvbEoHGcYaEWpyUtYnVm0x2fkGz9usRMW/3wOSTmVszC91Ef4bfMi
RI2HGgzeqFTg4Z0u350NB1wEZb/Kt+adZPYJEckZi5/AmqOegvtmM2QE6kC0JXIq
kmfV4weH+xdZ2f+Xq7qiAaS8Xl0IGUpbwZ0XelWF4zNgh2qgWQUNSe6XccAUTR0h
cF9xUGjyFWKJTQvWimVuftLFg58JbFexZiH3X3/tfCKuMJsO7r4FsK0xXmeFjjNV
AQiYjT56mLi8zG7ihkUuHB1kCqKSwuU4Smrwr31wvvCVAw4uzU8sbeMpwndWFiy3
3mmcP5zavFI8+NpvbemzlHEwrk7sLD51d+BR9Q8BAKuMiVgvJDPE4M73z2yne0uA
CxNRjsR2hvtf5unZcJGHWXvdUbqTQjlbkMDW49j5Yxx+pe76M3fwqiQB2QHmMjnW
KLarHS33QeM4Bhvo/EmA4y0SmYAsyyHj6QSAzLQa6KOk/dnWZGyoxUbPag6TAUaj
XO5OXEQWZGPceyM5WFLfP1aelY7E4qEKlQiTURMhJ2/s/4CNAO1G/El8qr8Zbbox
qYK2tBzXKqrE7bcqiXFO6igYu+II43aojsGHXS9WI2IUt944EQSMHGcasjgkoPBR
+UX8uixEoJMNT+kYWSbm/5M0qGICODJFUNMhNPNa2GzX+bDwBce/JHMZxAUpAFGo
eRCtb3aplbQxcK5bAFFyJOOD+dmqcx/b6mJsfbwm1BDXSeBGslJkmqpHZvh7l7aB
D9A6jnZZ8KWJT74Xt87BniCcKFLPMa+vruNgt7wqCr/8PbO/9CulrNFAzVIs1yPy
Dhq9yGhGcSsPVuxQU6U7GTJ9Vbj8Xww+ca1mhCH9SpRtcEDYER0yFzWiXARuG50y
JX0EgsQtI83PhKMpJmjbExFFODusyyy3QUOvzcYALko2L76H3ZeZmObY7GrHlh13
LzjoOo+W9NEIwLcY2s5Pc3R3I+5AwUvVLg1imiuMLvXl7E3pitPKHJaEVwWxDdJX
JFRCdsdehczqq9b/kbLwvIjPlaS3g8mc7JxSTdOOb7TsMwIUMJDY4IqxW/t7OVCj
B+8ZI8dveXH03UdKx/pDeN3kWj4EM4lAABbxRWxFaOwNwbFlzoG6ZGx0J/1/peDV
wJhN2icMs6acmEW9fk1rPXkNOCOAh4ut+SrRJ/TZDeatetF4yM0DLtZ/HVT4Q33G
8LAPw5RUZiCCmiCt3WyjdszE9Ptd07IVsTR7g8c4G+nw8KHsZcaub1iksdhmS9hj
EJTTM8LOpfTNJyhwf3WLF5dyVTjqFaOjEidt8RMeWFBzyRkC7Uw7CNeQXN5kPPie
OwU1rpp1EHt5qMqJyRaf5L0wWgoYGji2SLyMWYlU4VTs7Et4e+ybE08oHIa8Fdx8
+UtoMfAoA2XX1fgcQxZ1Ei9PDK1g+aVjWgC5S/W2Uvz/dF/fmDdQW2zBj3pxt+KN
ZC6nFKTD78vU50C691hfkTBVYpQ2+dR6Mct+5vaNNz2cbH5Srm0/I3xuD2E/aDoK
Zedb3KJ421H5XyfK4Jds3pZTlGeIxv5bWGXZTjTNaXVO3mrxOenO2ke4ZDbsgSbH
j2lgTc2TmzjoepMBb1LQjf/NK1nOWu5/mxj0TCTkQPMfgFm7fEH4vNe42CYsXDKt
ob/6yop8ugebSK4Sva/ONS87zB5VBfXBJYYXYoqDozAnFZWU8Zzj1AWPKOOXy4T5
dHG6LcH1LkYy6eoPs42Cpcnw1mgN4rTjadapsdOBN6573y1GPzA9Kpj66vDEKGeu
+Ar360JCWjFyG7fWv1nNGuPWrAS67Kg8qQz2dcmWZY2UYT/y+fANQHteid84pb1J
i7r8QT3fa5qOPj6WphPt19h4z28PerDMKhX/khDVKf68dP4+LC6U9+KovmPO4z9o
O6f3KD7a3P2fd4RgvK1SQ+AajQRob6vvvhxCJaWj5YcRpVNuAqXbV4Apy/XLTxLt
6OiegQdzJ4vg2a/h8+n0+GV0h8EzgOJRw6FP6/PU5d0vlV68h0+LxS1tDANEu1en
QuYVL3HksWdsn9GC89MOlFLAUqowa77Jb2aIDj6P50dSiYtgC/2xPooidb5iG46w
PeDc3KA96OC76pnE1u3qZ479fIpjBdRT1FDr624op2Loyd8ibbS26GzOPEAyGbhn
RmFPSpG5ChlH9tHk8hRFbr1aWpvDBw8AS9R0V8ud92bCGgIZx4s0OKwWuKf6/vbS
XxMPE0sBtJgWQtkSfs95hUUX6ZOUUAU3vKuiLJr+r9HAkRITvAfHB/tW+HGGryU2
yhE4soGdQR4cGRfn7coygCwxjRwPPKacZdf2gSsnLRrB9taf17z0XaBU2JAi4MCu
u78rVzPmIJwFNrzCiNgL0mi45UIBS+Jmw3vQVOUu5gV4PJqmKaLnlDtJQpxyEeAF
83081JhVK2MTpcrli5NGmLb/1bAz5m/Qy8VXViT49iaf6P4JfQbndgd/tv3/FIg+
n7ps9sfIBkleXtLNfUyUTcyB6nQB8EoiRd1UDDGWB9YGCovpJOofnjC+dxTlZvvL
JOVUGhHm0/YxI70uHtzaYxWy1B9fPPydqD3gCXYBaZDIoAN/4iq9/uJRoOrJbKgu
Doohsg15ceNe35nekF0dKARdPly7Y8k4JBm02PnKk//32Q0vHf37/yb8jcxy7s8o
jybtreCecVjpp2n5EGylapIgFKxoTvgTzJgi+JXoqAS3z//HQToLH5SOE4jqkAzy
DUK1TpOg9k7R/CqPZY07AfvLQYJQcNx68PDvT8/3PEbs42htF40oxib4eYD+UhkD
zLATuV22TYM53CI73ltWUNLs6KSsA/Z129CLXuiOKuZbKmjnUeIknUZpiUsh8MqQ
NhD5bjZVEKfs72MEoWIxBckH4n2QQ1fepMVHprtE0z2Hd11gBn5L7HC426hMahxQ
89QQhAXTP4/oJKvBxppn6KBZ/DMfd2Rv9D6ZFf++7meUjhEg9BRtD46nL4CqpfM3
mq941TQ+I6tzjLs2JKLdU/OtPAhfwxVYlLZ91pUw+nypJ2m0Pqa1vB3we/Rj9ZAd
Rnfto42NHwAk7R+mh4pNHK1ddATGrliRTYXXkRwMXUA8rY7YEB9/nYv5TH5VWxRI
vw9yeO6olGkAB1s8PkTPszREV+4J1UD939Q00yLKCG6l2SVj5DJ8ZgPeRqGK9rUF
UeKROI+raJh21iC32QolQXPt4J3BovAX7xvT2Nlu4X5IPa3ytivK6Y95KrqWwdwF
H3noGajx7uu4z9cDMcYt8oioxBSuZ7UwOx+QMI5ZFhSliD8cEYCPYZELJ/MZEpIs
AC5uO8t8ZjQ73fs868iMXSKjW1tzddudMJdOgXvduiLC80keWyE3qPVPKOcXM2Ap
gE48PywPgKCg8IpSxcx1nTmVEQ/HCxBB5B2eju55yV6nIaWP4cDU7zkXiOent1nC
y38KXGrvUC07ZAE9RFgRX2t3Om+783/4YwbjvUrdbMv4TH4WG+3CWO0FbMnYVLRX
1P3mvq9GLB8d/s9r6rYjlhP2RHQRLOMiD2Pnx5MHUrEWseCXlCAfbiQgJOpbZ6U7
zlobYhSKFeO7lqUtiYyP1xzDyvgKdF/hvaVYgsBt+a1OuFNFdP2DrQFy2xaxg4hV
+KdUFJXCWPaP4xfyH3jnNYX//pAyHdhMBKl2Xo9TrvSzqKnAwQdK0TvWkOtmiJTs
WuMjzsKx07dsiQNgb5LQU+Al5SDqIMT89x+85Yz3M7eB0HYmBfdbXKpLZo2Mbz9f
irkvtaJL/0BGUGz0BK/tRc5cs4xsIdBzZswpPPvgxvkGieDyAbg1iJQpW10gUQ4t
oxwlJYFKp2sJOwRqctLTO01S/e23Z2buoyTqVp4CfyT11PX4vcmQ20ut6vSob6s8
VUEN5gDEfkQMhp22lm5V8xDsbVyoJexaxMdTXIquDB9JeeI+QPLCRo4TJdowYrjq
x2mTZo66/P+KvGJY5KEMhO0PQ+4ZLzTmadCzlmL4NGpEPyY5a0DdRdqRLobj74Ii
zNqrkrEkGsPkY6yB43hsW8HmKJ3pQGtFy3OTYgpmCixDnozDtMJOxSKCvZ+Iy/wR
PJbEKsHKoGxkirMAPeE7I5WuGF9JVmz/QuRUyDIlJrHupCBCrDPKfk5aNIGf2nJh
DxiaTGRE48tKRNScmzEd6h5+nN2+7yybGOmXadj6ZiTjgNnBvzadz27LjhKICEiC
sZfgdgmqpViDB2Fe/cvBLViLSOdaWxcDL1Ex2uzufMU+PlyYfkPQxeX3vPDSqtgC
k33XfkG6Kbqp+gN2ren6Qq/lPzk2zVFPTLtr0kj/QfrGP2LclrTl9Zir2gm/uCf7
7IXUtzHqNyrxnh/JzBokBCHIDWk5rQ9Xw5cphZVTpw79oEAh+hdNPEE3n2yDs7y7
ymHBzzUorpL69CrNVF77BtBcXmwEBuPw+wZwq/dVRFcXfrrI0Dby5go4ID45xe79
aLqfJAca4URkgi4HJVAkJ/m0JsTZc0ijIG1QI8bEPiNxnfsFWxEtEkjJAZJp+kSP
TPlr+5dCFNX72G/Szgfq/xkojdYzEwJuOTPEtPf8pZrwGL6MijN5YMQ6MYshBRJU
uXCyc4nPJLYhc1RHakH9+xuI5UHC2K1MEqxYSxZpp1ZjceETst5l5/hF9xXCyXQw
Mm0B5ZLDS7ENlfMX/DLJREWySq8yTBAaZhBlbgdX8JayEcQKsgIkMCmrFswzYkWB
ZOSKAlPFoOn9eLSzvDLHkXsCNRDxpwJn8f0WoBiytuhqFKcGVPzzS0FBLciD7khK
+nMKJ+du/9YlbVVn9zBgid9pB0HdArImBIHyEJMMS07+JXo8XfyNe3XcrqNbwLQJ
BPg1HuZKVIZnFMs5ieTzXxzzgRAtnCipdHZKNxtOLThvg3DRj7K+GKflQXb7KZYh
J8K6HMH+UofROmkSvPhFxRv97JOoUG1vB/nQMQ3gPtUEAzuhzResj+XpLb3fQoq2
T4gndPbkgZuArB7BF1oyuggsWv2DUB33cTcEDH8doALeWGn1DJR+UUnUJKudPz7v
207qfPpvjSDq2oxcY+LmFQjrehBLNlGzYewU4wW3w4c2SbKKkYhjeYqKBaSvnkAR
GFoJJT37Xj1Mr+TkZjPbU+QXB1AcAFQctOH2oH04KupHBDEj2XmuAOzEupy5Yb0q
va/ZopQNs/W1JKPRwjOQHCdI0GpqZHJLvFSMSgBEuI9AQXHcALSSpu+f7a8WsuaJ
5sK+HY4OiQrfIwTAfyh1f/OO8ul2W1VXz8z3lPnA5Q8sz7zg0whme78MjbaaH6bR
+5kYfWAJUd+l8w52BaiYI72z9U0R2pAFLUpdefcJCpML8he9LGb3W75VwSv7pdYm
RAJxhlaBQNo9hunKcj8VBNJdn0hwKBcrPUoNWkk6duLBjTuR9+7JfFC0yOpACtAl
gRc3CLR1FmxYC1Z1VxrYRdONR2n3QZ32hNH1wwuxdym+fgctDQH5Yj+S+xzXCDPA
653JYgg3zlL5vzZF/yKrzxbgNXMBcChXbfMcJzESM1ADFFJez/RMflSZ0lu9XGKo
pYDmhIZEH5WD9/QnBJL3Fz0CDGkxW/EbVDg6TlrbfYyHTn1DQlyJrGjCwLQUb3zz
FIZLmlOr2/A7+7jMfesAyAcLZdXKgN9HCxHoNDe3BAUE333h8KaSI9D5Sj3SYGDG
Cc3GXKqZCky/LK7QbErnxbQ1c00J4a7cdbXP/la00O5ZCMNB4uJo1v3WUlnIrn0g
TbmgLukHzFched+o9W05RE1LPDF4GFw2MAG1qRtUBJssaCYNqg7X5OKgjlUmHB/p
SK6eqFZ+XAZzVEzSG22tY+NCO1bX0reVmVIx8FMuxxhGf8RKKF1MVTeGMY16TsjT
Kyh5NGk9FVv3UseZ6rRtjDc+ictMN7o0NeUV/ZxnY+i55xUuiHzBU8mETFSso8wl
331ZYEKxledWEuxov/9KHrL7IJU6HAfIjI+FK0xoOgRJHhm27p4wRo7qmdXE5nXx
PAaWv4q3gWUrmiGcYrgjETgBxGRtmd64b7dLQ+ryi/zTGXDYL77dbbV3f3e3IEIG
zWJYzyubqFLKTzLzu37978TwB/KTBhT5LiKAhT0mc2KcJJI7UYQeCbOiy47ZV5DT
Z/1V5eegzE7j86y4vR+gUYLRYm3ajL/RlaVGsn+ywPqjpr+VWvWD2+sJJ62YuklG
mKxPXREeOfMw6rO9qCuRX6yGZsrQGcK58WNwx9Fl4jUCVTCAumyjHfWQlE80Bhhf
nDPauczFHhRMtmtFTamxYTuE/DykBGdoV3+lSD2Nyp8xrTEU4uX2TweBEDH/4VAj
xMPoDvsNbOoqR2MmJxncnN0jMelN88cfuM6EN4dp2VkF+3fVhhy5il1kU9zOHFOe
fCb0uXhCeXLM25aVq0XRFw5hfvv0V+R/5PtmppsorLkfbSoNKS/5bcji7k/5+GLw
uqUA8NyE3872Q8FTSTA1QEI+qWHoU9tPY1Jyf/9fPl1P9roQxZBrKn9+uMwcepca
D/QrJMStjABzzL0RJlnGh91k0lRsvdBmkIv47At0Ujq+gtpUY+Hk+P6iep3x5ReJ
nQ6EXyAr5C5W/ERRi2Pbu9BdDhCH0LNK76znPcrQWWC0+PLwpfYR87RZrlKE9GGN
bIAh0z7oSZZghZ3PUdH0HNR62Fk9JqJrhKVAoYTZtWG6DZjl12JPAz+YRVxGr5lj
jyiPwEvhS+iuCIvmgM0NJcZ8UUD5BPsneQpR8HGuhGXuYV81e3bIWSNYFOD/0oai
wI3hF1bFfXIcCVfdTRl4lqojBPfbvWwpA28zBRuVZTmTlLFB7VKZh177+UiZgWn1
aMiF8rYEcVlbUDjP0W7oU5FnkmEUIB7rKrdBj9XEzrUjgtf3pgMJlhjh8VsleQl2
ttokVvaKZWOPJRZ4UFGb2g9b/NzheZ/piuTbzyA4ktyGf+Lk0y6ynmDWDpC4oR8+
bL4IEavV7D3emKtgOik6okR2KZ8mPyr5RktX/xGpRXklnhMO0kE2JzdGapBgTQCk
mqcLMiffpeRGXDH1X+pSfHskdzGuUy8dV2BQoSGD21iS5rxNHIsGfwFVhoOZyK2f
59x9n18+o7Hz3kVHY+hYNIguJjVBsQ3vmDqrO65TcwIHSPWJdMPGgXdCETM+wLsk
JfaIhWh8dV9zle33+J/jW94pWwpXZeaQR3xONj7N15bWx7PzNzjgEUsAfj/TuAWt
mCuZxcObMEg2MK6LgNuQGOGPM1owwznPL84YXhamfyJ9uKf0nAzI+kYSdby8ervW
wlL7Cgpf5w/OgSLlmudxSgqh+f8ARJfwj3y9FgSsw3Ha7CryWHB2Ub4jbZ1WZSfG
FtAfok74cdlncjv+LVowFn3QXDBbb1UQTjpUjuMRKYWFpgMxCa0bz5h6pTETvmDN
+RNb7SZd2Dz/pIo1G6SdJYOLYaf8U99ChBkGMwdi2vm51fJ2PAUBNohcyqpFOyeo
STVpWHs4wTcjLB6xdgqXF8ASJ7TaCWHhXeD96XOnobfDo6EA5UIRgb+mwIiNBU5h
BZ964dQnNszE8SfkWQaPxFYU3rROBS3UjoXrJBl8wN8O2m+IKD7etz1muZDuxPQV
oECDH1XOvZVoBZ2Aioq0IgQZcdy78mIgYkzFAK+72uBeFraQklNof/mGnwqzytkq
RXW70ULr+lIFB6W5G1qvoMHYlbMJ4gKuDMkCcPn8e7TaEEQkHKoLxTI+YlpjqXd5
joR5ESCW28oI6ePYeY6eKIx8C5RH/OZ2+Pu3iyzXabxnIW0YDCSUU6Y8j7dGM8+8
vpCURygycYeuGiZyoZaefoLSDnlSgTUIeV/Hpm0A/fVpflITmoxon+YHFgYAhBPY
mZp4Bc5vYoQJDJ5lKg/hTRH98Wlo5M+WJuyM83hYwVTOyZqcrM1PsalGI4QSwN4T
t1k1yRQqedyIuTyt+KsR4MUHTnC0dplNSHHfayzOjrAP0JLX9eA/I6HvNwRf04ty
Uhmmk0F2eSgThCs8V8YsXaguFfawOQ/siuKXPleXPNOLd0C2aCw2vb5Ej8o62UJ6
O323UeoxHeEDsQ3l7fOOC2UgCQ+ZgLJ86qZS1VPkGagtTKCH8s8hBq2Z2VRWR6ge
ilqYGpas+Or4fadttDTfjYWj0vtQPLCZh+V4UkmkLgwi9TMQe27ZKaXy0pxydw1P
pedt9itnMlcMvTXiLp+eydk64obxp+gUndDpvGDlnSXUhC6XXiKMrk8vCNbfT+Lr
HQJIXjkFjcU82Hn3D+8KZuj8WcTtXQ5nXBS9kkRCSWpihyEcOcVZVYf8r0EQuCeR
0q5pRQ0b3S4G2bo22I8ligJmSFVNdn0ogPAPXoDzOwx9QpPpR15h78x7F4XvR/Aw
9jNgrYQJxicTxYbLytGcRea+em3skFvjPp0btqZNSwzZHLoaESDlxkXZsgE/odSH
9+wwbD6Sudtx/sKubOiiTerf4S2vIJaK9Kfi2cBnzhC7p5M9RuiT1RCr993NUbnV
inlORZwrTRq7jNO3eitJHmdMfgsnwcXgCkNYSaDjCTqP9RncxSmrWBTwWx+igrJ8
ERvaQb5kAZKwJdm/n7hVkOTdc9BWOpcJaxqNazQk2BG0kHllu8mG9ASrG5eMy/6R
brZKlwE+1lnyEjbH/pwJeidbIytmE4uIgqQnaP90iTQpNR9raDB/EG3X+2Kr8dOH
FjnuyFPL5A7HFE9OPbQ8RQyxeaoDikutfsW2q9s84rzVq8t9TWW/oTk5t2dK3mve
W4yi5GG3DCx9MMehafmh6VbGNcQ7A5nQjEi5VX4pc4wzWua5gM1ngFICLgq63TDG
TWFrf4GxJhmt2EIIYpFkDq638yAnKB3jZvGfWCaeMORcgAahRTE5kREPTJDVtGnH
0eIWWWG57kAusTcojIMkJcS2TcfVQkKNaRUM5r6OJ9PYqr5sl1sXMdM5cB5/KdYR
76rh3qxv31CiofUOziNOwwhG/6snt2m4qZmCatDVt//mcgZB41/lzn+z20s0ARzo
AwKp335N9c6JY9uAhRJGQQzYDIZiEc1qSUx+sn6dkWRbEcrKZouIKjnBDkYBDAcZ
B91xQQj56l1aRQ7xmYZvsmqtIvWufw3RbKGUGzSi5vsc98nCSl0HZdhY9dDtVRWp
DaGtXkXmck6WlFOg7OFbNGiSUuuTDbJB2fOLObrcvyP2gka9B8Ls6AtuNA6ZsNup
/lZgXtZGmWoGCpR7lJHXYNsrx3ApjI4g9LPkgtLdA/2+qiVEz2tP0O8bCfU0k75U
jtNETfAFjcXLt5ATAR3O6HixYLVyFqMuzoyEBZqDB/a1LfFencSx8oRM3POxa7vG
+pLFaltwroHG+eGdR9bpwNIiGtcBBiiIkfc9froZk1ACB1uGSSg1u+PGv1bZuMtm
OLDOdfQ2NA0v2hEmp9X8IjY1lMx4eSjlbxDI2wWGlBueS2fdGgAvzAqEVZiURbX/
4YaCA8IUL8KFM6hNBIRdEqhx5AnRDlJBV7nnGKtbKDndvA7cmh6SxSp1aoY9RTTQ
hczLAK/jGbMBMTs7btTOOdC+LasUJVNU5Dq2b147/yQV2LeF+1kllTua3NTAJBS2
pJihGYKhYRP+7rA5Ea++++djV/oOoMPB9VM36D6uIdb9WQ2xFGIgugOU6HTtMmhC
oC4CTt9O3RHm5mqPQdaK1XiZk6xMrZLAv0KO4h+amtq9fypF7q+lKItf4UcA3GUV
zR4G86I2KABsvlKFQ9OgrTP06GdWfGYIfldnIfOxRIh8o3sBRtbhhB+dYoxqblc3
L4PM96w6s4jx43EF5eJvyLBnWFAaxnFLgbo687G82Zke8/+eoMMB5pYgOrf7V7Dx
yEInnBzZAU7WVnTAItO+Mf2iMNzhej3Xy4+a75kpt/3/EVNz14p+UnmNFDnsWiSk
EgI+msDWHfN7w27k0WnyPORvGdxQdLxZQAUU8/Jrk9kaPulxhXhPTtI0Fp+ngmgw
8DXUhmp97gZlP4a132FL2+7kdkwv4wLzQqYmSHxuFQo1MRrLCFZChOJfR3ZzgUPX
W6VeumXNv5gOS+tDNN5gwC7EKIskkQquHcipIcZzF6k4vixmlTMJOB6D/Ty5m5Hz
k3PsVsVE8nD38MRENmM4whJ55I4cKV7kofKphE0NsRFCOOQh4GcGkvm4LYSYyVF7
sbjTSKHrP+xSO1fQMLa0rzmZcKCj7O4Kztwp7q0TkwpWcG9ni9kjp2nC9KeQLUAd
1P+Xto6B4/mLX3vR00mdHKe2ga37QhkMbB/NGUqwYCXRiY6tKbP9abDhrrI2GcBS
vHXFG5zDc+WrUMKIuOtFKj+5ky20xSwA+Bd7I+1O2IwVFjSw73LHqBvqQelJPR49
KBqlEL2qkmd54cmSmAbIoQSfWrOsbte9zy4RC1v3aNV4UW1gbCtGfC4tsfxyCJ25
rizAaF7oxMXFfFP0acfQkj6GAHNKkCHbs7mh3g6HqWTabA/p0jHQ/N6QnkWafIzO
xzkw+WopyKNlxgyJM9oukZF6eAEztntyTFICw9f6yi+muF/aUks6K1CXPNU8uCCX
mJyDt94fJ6wqijGtX/yRKYN4esbxWafC+E2lf9CWpubNoLyf7GeP3cYZRtJSp5PV
DPHLGQqEr90e1hVMvCSfHhgJxGx0lnytpOKrtw9SV6knSKD7tcis664s87Y3Y22a
UQ3i/hxszd5EYeEROgEtcwm0DVsjN8XLvJkBOzfA7/RqUGTiHRFXRJKxhOcHyZwo
nLftdD6LXjx/bip3Wrpxr0qBx4Y2/tGoXj053O1fWTcVPU9IctvHan08whtdH0po
hWIFeiuScxENCwC9bdfymmjJfryUrdc+WpK7zoV81+AmvHTxU3mTEXH+K9K1IVYe
1VDRPaeVj1spw74EXu2hUB69+W/GFJccFjtN6icl5/OFoi9eCMRpHB4Gb1wWB7b7
zdQH6Y786gS9ANDXsCAbSyss0gNaiQ2rb1A1JsrJVXGRrEVc00OGMgsuv+EeZ8tJ
6h386obrExmEV34ilY0kQR/grXwiVf9OCrd7gFiKyp0erIe21M3m3kPauOgPVeiC
2aGHDujaPYagjfxQzpdpVGAeohzC/6dliG2vdXS4kdynV6+fvhuyl1XVUQ3g3/zU
eWCdx4F8yf4zw8Jy2GElgJo0qsegmt9IiT1H+WSwlRKxo8Vp6LhcmzUfFa0qs7ph
Brm/L6WASsQnjbb4/cfAUDJsj3KiFfmEkCBRRiVV0e66wGoScyIACife1Ma3/BMv
IpMX9xz3Pu0CGpgt2ssdcV342yAv3lMT/scy+LDk2u9GRtqMjvPCITGMQt2KedW+
NbYkbjqSXcU6Htg4qWMBweDuuprqMO3TBzCuNS9PiTxLca1lJkbmApczoGN7UV90
tFWH2cmHKvsl2jPBtsFCYpiOXDfWvvcmHfxFreMhI7IvzwtuxgPs8KtDkFpEuZu9
LvJDYST+yih9D7Z7L+r45srMinfewVia/D9l7iwI7NqrxoiMCutzHuXLQx90o+00
ulX/NHFDixgxGzDUHR7WXM5yaSnPeVCBi57KRx+WKwam5YWe3mwXlbdUNR9vDlRf
64HtJdISew3g7jZ6Pe4FNUOyS5Nih9k0F1D6yXsnz2MpsbEVzWVQKRBx9X4eTeD8
tScCm4oLLMlXrlaFi4IZMFEu5qEQNzBsQMXLaMsjx1gy61RWvJPbMWxzyXdPzC8D
GzalV6g2kLOBvPcGP1m6MicckH8FZUymPWNUShbfNuMoZAhH1D0PbwbgVVVrdg+C
SRoV2zlxaqicpT5m3AzoD+i/YU8u5pqXkH6yk9DQa14hPNSIzS/6lxtnVY1ykCW+
/La3beI2qK9NNwA7RanzVb2DIeC0lQliU3VJ1OQJGqbYb80EbRAxLrxzt+8Ua/L5
H7qM7K2KNbMLG+FkssaiiDdRmKv3kYcOCXfF+80uTD+FXv7Qa8x58Jfo44p9I7TO
h5sL0AsOLscVyU96BoC7iKJHs7FgCgZD0iXdn5eNSMbu+RviXxtTJ19ozz5g0N14
oAQEh5z2CwO/VxBEpMantxYrwewPjUya7LxFV0qambk1oRNYx7hEJp9YHiVoVcNF
e1YjPYqIZduXAXClIKzHt9sSy24LG3zmVui3x3DmRGifnUoCoTmjeN4NsfY01wF6
UEgoToiPpnRyr8UjPUBNKJ5mbmYGnXRHugmTTtn/MxpaREOx7NxOuQGUN9qEQb8A
FLlDRx/P+J1uW3r/CzwMKlRQp0k/y3BPuHIW/SlxNbDNl7jnXw+gMdp7yDTnRXSe
UW4uRvDuusXelgaktQakwU/FaeBnf0GIM4HLg8SeZSkV297joymQ3WorFK1NoQAu
etfc7rPaXXRJ4uN3yQd6To1ENI8nWSP2xv7ChqsWxdCWkjBos+CsbF3/3KDJj3qq
Hw1ZBw+RBtyS/ZU6IQ3D1lKs3u4imz55eOv45x1sPErJNDvpzitdbTF5ssJ2dOga
e5Bi/o/8KHx4DcynlGn5kzee1foPQUGrYlGfq3RfOl7bulvwjcEJj9WrzoxBBIST
udwAEkg91UsPtIK3SfkGnpJyXAcgPfz+Pxp2irbkLygC3Ml4LxtWgKBXui6FgxGg
N5MA4Ux6rOxUvs+YO/EbQn8tMST7ElNkIw7Xx2I2cMDdYWNBqL81/BC2qzgGSoHq
1S8CkjCRpo+vaFng3/GCeP7bt0fYqTp98xhhkibmmzN02iLEzY7Su168cAmUbPJj
yimW2EAHZrOtQ9LyhY3MelRbQgDhCsWw6FoQaMLMtRE/svqVlegwg8Q2o5Iuoxqq
jKTe6u8AX1a5gk3CqBax14meeVeRP/Qw2h/59XJfjSV4q2/FcWASpoXMeU91bgZ4
Hzs26sJmZ1tDdWC8dinDPmdRh32DKqfahSqO+DBQ1PPFonBI8Ge1UwckYY7Chbex
PcEoSaRr9T5kAKWirDCq0JmHmCUeSfoTuISwOfk+AV595iWdYYxke9RBg0L5C0/i
MMJT2Q2tJ1+toCs8HPNF8dA1I2EtXxwDRYhCamG6xCk7EFi1GALcSQIvQ5S1xPgl
5hs0NcpC0TdNv98pgMzppF0TyxWw+QCiTax0ihiwz5SIXe5+3X4XWBRoB13sa5sS
5CVIhJTIHxR+8ifivleRVU3hX1Y8WjB+S5d7Syo8MaOBUWb4uLOtfYUo/NqK1sYi
Iz33IkD6Ay3wfWM5BUf85pA5S6htYPJ5+y/QT5p7mNbHFmjWUrl8JqMTNXS9uMe2
E60UZJwjWIt9LBu5hwFIz8kJbWf92GEpcaKAQw3npCnBPZPg+LBVoDsauTFoVHJh
SJQimN2weIJHWtYe+fm+J6tG7J3nWTEqaTEWWRooLqMjkD1IezKr3JNXrMPXHtQu
CTkAuTd9Utyas27bx8jozlb4I1PSOTimHXsAjLMIntmR9oayt0Xp2A6oLsaRpL4e
n2eVuwoNsNMb+B52h1aVMNNgtMNeFSAyA0fyUFI360uqmPutXciBvTLHfvfVzWdk
7k/0C8fYBgK3xAINlPiA995fShu+zaw6UkhxJZdE3yyk+jfMi3d+8usSgquN46pF
FN2ho2xrm/aZ5YQSaQpGYLX6FZtNNCdyfD80OYLKs1hSExPsXffwxA/jeXlIGNA6
SpSNPfYPLKb0zhOuGiFjIxbkGpkaZvQhxvVQgqjNU/X5zCTJyHGDrVXn6hyJyzdq
uadIike2TLiQKpxTPInz9KDnX+4AqndMsxZf/5319tqvmO0OJ/1lCTkHqroXK7gN
xTLDLOBSD7NnTi9446o28lE9Uvd84usNCMgiRNB9PCZ5RUPfEOkXsoa/3S+IUAG8
UwYeaOhmsoDS81XYw0LpOft3Q9XqXq1L3T5oDFwAKkFFr6aSRnlERBp107pMsMo9
vCfJpAqi41V+CVW6zZh0vgT8zubHNptM018ZCvwplTnaEFOigrX7eto72RySkeZJ
lKNgSfqxOmw1DNDJKDKgpOFh3IGZ/9rmTgal0ANPOtRPkxlm4/5EwGe6ZUMAZOUb
FSsZ7UsEm7ulhJu9pwt4zD6OtW87dwCjdibvOgx95/bj2B7oJbMzBOFvM3+DFuKV
pNpTkiOGSfQRKhHSmeHrnel0RvxziI1aUkr5O81R2KLutnmu+DfpMVAupvnxSQur
kpcaotyw5OKsExNinO+SyjG0cR6DJogaGvQGtcWml3UNlfjB2xouurbQOt3JPNPT
isUIKpVNY2pYzFg98Ff5yPAHgpVgRXj9Da5EK2Nrh//XkcMQFLCSb2XckBj3mkFt
dQJmfxkvCC/ZbVDxYv19fk2bGCJw1zxLX7lF/jwwYF+cHWHCmTL2AXId9kffEoKC
6ntQVgzg2DEFC3WiERcfZyer6Nh9vgqRQxl2152vYeDjodUoeOfDlJPaX4FSp1vB
0idMOcmscWpTrtplfD05RNUHIsfHeqGACRJHBZy2aG85Fv71td4NQlzWIe4ivJPo
huoO2vHtcLshtHehYnM/3Nt0NBANEK2Nqcm3NQKb9vY80ZshPw52cLN3mJLdxUwO
kUkOmZjmIGUJ/n1dhSjmTnnR6IO19KVN1nEWcU7srH9v+vgLEO0JGq/7S15RAp3z
y2Gkgzpikkpq2CVHbkHcoH5F4UitonXr16c8NCfD9xMBNxmvhAR4OCLyqltJTtFs
N5PJzZfJWZwdVkpsg0HAPKuQXMcaSjXvcOKB9MjhflLqbMtH/lPkdcjYyoMD3x0y
YbeyVUmhz00gzQkG6WZgkPsTI2oMzbqq5eM37cA/KbOL8dJ0ZfZQ5nz12HhC7Tt+
xSGQWLA3awLnf3hsFN85z2/KnsOxgQE+iO61KhlEeqvq2SUf2YmYhuNyiA+C23GY
IVgkBb9PTgalA2e34a8z8tRQsTbuSuZL2I9Hs9s1IF4LArPyfjx00KZi7ioZRpdb
IqxsHUI25fcF1XwUVGeMU9FbHAcvV0YLMxyRIxNL+zj5Gl7YHbWkzztl4mL9LUP9
PoKgyzgEMGXiPlGHxSXZTihP+tzH2Lks3MSmK6zC97I6hxe0T1KJkK8DAtiJnTnG
RR75FGf3WsRQ/qtq9jEZHX5ToduoumK++GLIipqCLoU1YOgNbrrFm2GhmQjyz9vy
csJ3UzBSOihDBDbkpaG/HFAwe+Vzws42WCXqHWQpcY9vxrbASJqDjhThb93Jrktw
BNq+u5K3gkyoyLtkBm0jgq8/8TqWei2RXWevz3M4mwBT/zhBF27IhsUygYX4Aas0
pTr7dcNzxAsA2+k49kKbtZmczyxRqmw8hTvqCgZzICxoHRzpMCVMor5T0SKFVhv1
51iuZ8ODzbAbc9YBkokyfMFtBLliicJJVvgWVLSy3C79Cur9bjtUztD7GiI9sg6c
YrPNBksI/94YQOikab0srMI/nPR/JfH7wxnhKrJ7/0UV0PEGnwNnyWRIoFFq482d
I6cAP1pk5S8ZOLOTqnNuPtIt0zSbwKf+lx1/I10SXJqsc2XTdRGIcxMf28g1fXiA
WeT29YigjUgWVe/u0iS4pzk/oHp0514OGCHfWP9RiTmxGyrM9J9BKuzjbDJ/P2wN
fj36SPlOe90UxIfsOPgBcsnE5hMvY4wRisX6+MsqTlubjf+wiAnf8mp0Mut0hx9c
YNawddoy+QgNXEmRQNN1uLwlqdpYJTm7KDCAdQauXwXWXl0ebxmEfwS7Q6VPh/mv
x+OnfFvYCZzKJGuC+PSbUPpg8HwHA0aG+LrBWhVqXCcoyY7hMHDfxK3PdawlmExw
0TDgTzRE75aeqrIzK3PtJF0f1iveEZ+4ZTJpUqA0gsLT1zdCASQwHUvTfmuEyeL4
a/fYs/eiInUXIj46Eyny0zoEUyXrtkYFJkHl0BwCG4pgqWKB9tO7vr5QqLrEKkAb
iPqj515oLQwPNfWEHsldcgWSm+DGBuELvp1O7xTxgrEiTS6QMmmQitGWwNwzNuTc
MH7WZFBqOwM9D8vXwosi18o0ZUAgds7rTnONTpbP5NgVmiLKZVoUd4Y+65CP858L
2tmMLkNiIHbWpHaRSwLsnZ3aR1mcoOcNTT89hUwWco64BZa918h+Gk0b6sstcEKV
U+HCPyclhT9xsC7rEyl+yg9RI3nF8eX+AOJWzG/IojELiU5kiHjQ8nTkz2f3hf2Z
ASuURXNSWvqau06lqDk2mCWQ7fdHEftlsxV5Ul59eFFKpGUAogP9Clr+ECQ72q+T
TnimLsCsMVFf7hrhUJd7F1Oh1lEY0LXjSdCyN9aW34SgPxsyh97T5b//qv6U0p8j
e87zAoJbK7pMYOcSngs2rDgMP8y0PDfwiIBS31F9IhbWVwe3njYIXGLrISblttZy
2Mu//oTZ4bjCQSIh4LDVjYrt3hZ+PPq9EnVjORZUdYBIXZJapgCQgeP42wJCtERS
ObELa5EHCx+XisuZBBxcD4uN5Nb0EPeqIwQh4pF/xropq/EhkQPfKCUyJAALJbsv
O5tHUAL5d3pyQOj4Gl5wZ6tHK3rvbvD3lPUbu3UUGBNSHdyRmQPC1pDmIt/EvqOk
SxzaABSzZh+GA6qVd/q9k8vPhbcrnwNRN9Z4ZD09kHChN1zyQwQNP29bi6cwq5e0
taV+zjQqF4jP3vErdWeprhAgEaRd7ntsxQtDmXAsPzbdy27cvj1FdPAs5SCvp+du
OlBnvDaFqzUvrXTLsBzahZ8pPHOG5oKEhpWUjzgBn0scRYlSw8xxC1i/s6GEc8US
RSItZ29stM2DVJkcKNYmYzEBXCk4sU+hw9eBX+lhnrVZ1ukZZ6OIspEXMGvwIHMl
bPPoYUPBINl0XPobt8jmEMw4HjdzxWfnhVLDLPjzy4yiXwbBK7AM2p6zm8krGhuc
bPAAGT+arU5i3rIMtYQ29tCf9Ok0e5Q+Aj7u8/tyGXwiZz4RhKVtthVt0WGtK3qe
Vus3cOTXBcyZEaz8rLD1Cw4V+yEbqCPu0GxMNwWd3pE93m6PO2+SfvObdo9bfbec
xndupBE35ocsBIZCV9phGHVd9zXjU7vrAQKRp8vgmiq8smotSApYqVhATqd+2zLS
iFeHhQhoZ8X8jQXRuZecdkEnXsTLOZ+KvzLXBdMegoW6M13OCz/opiPQL2HsgJKm
XvNPpWw3PTZ77dxYvBHCoLtJWt7n6qZDVg/h0hjNezza3SRtlCm27Yt05Z3oKPHG
vv4vKp87x0TZ6TBZNxD2C/48lVSiZQDANyqCQaRk9pTLuXv9Cc4cv2M7GWjXqV4r
mCOsG7E/OlUhY4hshQa+anBi+vRtTD519pBYeqfkRJoBblR3ao4ebPRKQkF4k5nG
BkqdMMv3uto0LxQYnATcM0lUnNFSy/QnvnrvQGAaQgnhVxNaBv0MU8cZkzdlHfQj
AaMVFxHzIiuSitPL5HSsUjaxnCEZiL20om7dqV1psjmhCJPZds6L8vVRpyoRpWBv
O9NM4MKRf1ypCvCaju+FFul1TpA5CschgSFPR+TrE1Zkc2oBO2V4sfGZ+yBMQlfZ
i6pHO8UoMbVXc9RX1sqgROB8jfAQt/fsibvLzlkxlXRzGqRiC8rZa6YCOwGC6tUE
TeIsVnTVdCA69oA8DFWCuSNuAUpEbTX8mcJS3ig+YHERJJB8CsGwgQTsee6g65wS
Tnc8xQVhStyMxrnV/PPY8V592hoot1FalwTuzLBmxPY2lPyPeY3SoXp58NhtKJ1h
sefHYfSsUXvUXququWjHyI9dhI7enFChoIkyEDl9pDnoCDWDQUgAaNVF416zOQXB
GN7lnF+5QJgInEOcT9Xe4iJVQg4GEv/yDjhMqpn2cJdmFg38kg1j2BDTQfzyKpVn
8dB+tT39iknGyKt9dAjYzsxehzbg3eXSXy26nlpc/+1gtDY+S9EknRyIAltLpjpF
99YBlPQTqEymWEmTKicImSGwU89R21+FVMA1XOipFfdk4AM901VXkTzj+nDagIBI
qxByiZfCwNcounHK3JEHQuKN1ZkcdHk5Pc0n/RU3JExVTe4MUWZhDUBXNnOV44O+
MAxYRkSt5QKtFi/XCz09MXh2eetCjlVoW4h3dpb2YZa+mJrbtT2cUHdLstlep18H
iT/msk0p5Zec2Rmz3ut0WywNo9PE7/W5ak4w+FtzVyaUp3J10qUgxIP6FMDziVvQ
hBoW1XRBhmgIOxCyFrypzlIojX5u6+QsTyjUkFvd1AlLYsliM7piFONRqvdTkilM
jhUDjTpuo4GR4aAlomwGRlZ8yzJuXy7lDRtYRBNdZDG217KFQobVqqORyK2HwMUZ
J90k8xXbfHrDaILTUTJ5vrIjjf/qqO+0ucNMs3X6+DafR9looxN7WVA+2HKXetCD
b4lkwllHGBIsn9F9urJ3P3wbxUtkcl24gPspNVjrwqAhh5lhPeg69g0TpLun2ONi
NhHLynlB+pTgSKJgcrNgxf5Nn0Ghwh3mvqpidbbmGim5IvvrFbqf2gEhj16fKt+r
Z4v21uSHMLlIkl9Auv2f1/J3Sx4iiX9LA7m7Zpsyl5q4tcB0Puuomc6ouJjhK392
/FaX/K0nO0OBh8qd89J1DJCT4ozpWUtrTgTRsq28n0s+PuUzbUGepiAJWbj+4i5F
kT6g/gFw3rleODpNL18dkA+OW8EM3bAJA4If2C1gI942w+v0S+xM/h3XqhszEvLJ
yWaoCO3WN2pRthPyB4KRaW/xw0fGTYZ49Kv/HP7WgeKa03q2PffAEO99+Q0+mde+
TQgruWtEppNfm3M/fQ+JKzbWMR+PqEhuWVf5pg4j4P3QpdQA5yuu1fpQfuprUazl
flyvK7at6Y1uI5CYfT3RpYuehpQ/Vt+B9BkwMqqpIcB/wflAH476Yf/U3fxZpEAF
g5tgFrKLm+g5FlBm/i/fyuqjl+3OzfKWk7n4R7+j611j/FwKRhoRb89F98wxsPs3
MaS+IlyVbcOozorO7ODTLcEbCROLtEEMSqVbvKpzB0a3SMtiISXu3NuK/mGxg1tA
HizuwRrBbefD4lOlQw23X9CAtFknh7DVUjTO9WBsn9ZDLWi7drLChamP4vQzi6EP
8rTJL7+GkZMb+CRaLU5OQnN3AOC2P2ZWs9JWYETZRFfeP/UohtYlHaT2iliqxqTV
UTfzBJDKI6KopjPX4UkwJL9w/gfJuyIZCH3Hoo7ZlJhdOAKBZ/k2847fH1EkMRdk
9kJTb+4HL2SdBawyRPabJ4ZqLEyQkpHoBsbsvAC3e6ic9FwnHILad2hN8SZJs48K
y0Pf5flTJdYG9ErQ9u1BhlQM0D5whTUKV8Q58N5uRkwYjpZZPyDIT9CbcxTXmxGX
UYHLwy91E+qptoi1TQSlyFnnPa8nfTixDIHVWs8oNdSIR5HnGvxAI2ABRURF1UFg
Qxo8Im5uIdvOSonDANkyWP+0leZcZTcNCeBHs/wsoVNnL9M4hrMl0i7PCPCpAaOe
AfM5thCSFiGQTduUe28r9I4YD4lOBl7MFX06TmgZWQKU2opg6J+FX9XGDu7bi5dq
+LzPIO3URPS3t8eBNuHXlUsKUP3U4EawDF1ymzG6JoNQRXTCsi4QIHycuzVElt1L
TcfUWrvJLQ0xJdgLbdrckZuLdMQfqGdaROPgpRk2XRq9LzzJY1+wOsJSOqNHuG1J
FPhrFEqvcoxaJBqOVjVBgUUDqNUNubYVcGQlgGNM9IQyceBVSU1EHkxi4hQ60ljD
i8IgZDPGI546MZY42AW4jkamd2JaRkqP60bdfWjZSNnS0jB0+IerWqSJ/AcyEBGi
CusVPZnoEI5dklkp1EJBNablnEHdo6mTLzhPPXAxG+pXNnzgYki3qmTLHSibfhAS
K36ViigRgbqN0Q1W/2Dox4PHUQdDifQUg54SeJe0lh3X+qcPXS0zAXAsmsET3Z2k
ReoCuaP+U8Ay502m/g9PmK+ik69eEYtwEvLcj1+qrmvzKQVFPEQuyjeeK/zP3Q7+
jWYPqSAuatvF63h6w/W2KndQUygL0ezhgMIOfYh45Ovqzac+F8FLl2TywdYWeBKE
ut3AiZJK7/MM8tCtJ39gbAOD7vszyIxZNwnKkDSGGTRsJZwgiBB+8ptveOgykefg
W3vN4ExWzrS3mrPsfd+CIhMSMJGVBauBrXN4FjM7m0YlvB7SvAN4Oa065lEwHa/F
j3nSTVxTrQTzY3Y97RjTSKBjT2isNRys3W0+66SSt6vBjpx5hazOX775Vbq3cpp8
vHlcgH5BszkpQ8QBzrjDEM9VFXNC0ee4nuA8yUE4s5lBnqvNE8YS8ubDZTIi2VIC
/Hydb2ZxIpp1DECujFmjPqicHRsWxWu5EJnEfpiZ1WbpUz4HqXMlGZVWNJlJ0rYQ
Fa7Fbx300fx9fXDQ6xZEkPomJP811G+1DYXTOl1dOKopf5oimH/d7+caSbwvn3oL
Ssdrc3YdoSGTvcrSZIsGmCm/qPPqWPl+gcY3UsmGwasHFqiJlRbcYKA3PZb5UGGG
9pX1JcZYxiaNMW3UZxeRGN29O1F8STZy6bBPwhsmH3qCgPmyfrkPogTMk7d27PRr
unEhsJQ/WaC2/tUobE1csK3MpMtmgeCqIYIQouaYRgirs+MlQpa/LkeerHt3kdJi
AKhiHxrMdAEfuiC0eLlvG5Ir77LrqqY/Rh4/PXwqhli2leBAg+TrY1i7LRaavaqO
Y82s2jYyzCdhlyO9qUnfnXNGYngUNWVLDHqkRi6MGyJc4cEQjqASeOKWVAxGQird
qv7GyrJ+8IuUIhOfyhppcPyHksssgwKpt28A1cPJs4GXDHCcWtxL6rdUL+23zBm9
+kbhfUTjhMopYYebg+v1HhUpIr3GYJzXzefGw9uejArsQKXyk7xSpt3bC0TOLA7p
v4/6xgtMUl0s2z9dNmXsxAkUy9VUPTpu7ochyVOfCBSsmNzKiYRbZeLLxHynebV0
sTnrxLmyhsFNs2ReUAesrfOhQ/9aoXVljIvTuirOA+utEn9PlXwpV3FrRa4suFG/
Op4Q1tw+VYctaalXun+J8Pa56ICi6IMi6Q8KWPfNxV3iV/Jw5bdUWLoXsLuIoCh1
gVsSlyshX3pJy5OYzq9wf7nO8JnyguIID1TqvaRr7Gw=
`pragma protect end_protected
