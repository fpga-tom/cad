// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
N4saJoyFv8nzTncCFTlBKv7xGIa94aEHJKu41/tnJW8JQD0s3tbKyYgYY5Dn9zog
HMrmDsPV04FDdVJuSNvpP4XzDZy0hji7c03U8xLlWl5fgtYrf+ERp7ra41PdATSJ
s1JRSQhsEmwNlEJ61O0byjmHBW3oleqhGN3vRh+2tt0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24992)
ZjWu0Vw4DVrHBAbTSavoWGu3/f3ho+qMOuRfK7nC+6Rr4RJ28pkOfRlIFV7XlR2T
pUZChwyqgdblYf3tYMgUsiAhMh44wKMH6v8sleV8jaGtynCwfF+HnelgXOWVWUYw
BOmLexHJ09eIktDEarIODlAdQPq//dApKKcss8ub7E3BpDkS1iQl+zpP530luREy
TjiGS8TLNl7f+MeY7563TmKh2g4+h/jiZJY7L3Li94uQ7bSr0swpSQznSHcMZcTU
7f1qXe7l7MSx1BwDqGCGznZx6snC0N7Ivua+i3oqvgsJ4x5vQ9qev1kt0tD+/M/J
Kluws9xX76dofrU9I2ZUMl21YUZh0JP+WJJU5YMKQKF6ck2HKJrR3UcR+YFdf6iY
cbcgeBJ1ToANR6RYDHDCKkZrt/38UN7o2leYYoMMp1pjXgN5YteNBKMQWzZnn2wk
iUrBNe/xNHKKUGkt+b8ZXG6bDXSgvWecQVNMA4fggDKYdUp0rcQlihkTla/JESC3
I8DBn3cUf+OdZQMtw4eqkMKhjEMxzMsDQho6etPIrTAMygcRdpYOthOg5446A+FF
GGaNtnS0br7AVMheC8y2FGGuDoQKxbZ0vJtEM+ACHaHTTrNarBjXZSKzSe3NRKkr
HBQt06jTkhXP6mjlbbVgTOux7VTgLwEK9LsW5vrEKNPTenm1Oz+0LE9ApVQCGblG
X30VAOxxZ4KDfJcTcL+TR2F4K+FzsVgrXAMGh1WO6C9E/PyQUe3XFXwW3DYoxVZu
z4+x+ZDcvfGTqFm1ugjhMv8+xpd1hUvNAnaXxGBf/FHKBujvSnYgboHMQYUaSRqa
mnczgqf3ZNkPM5tIMfYqLq8hCKrecb0V7r5huIJbTPAzJ4aM8JOVKwzi56C5OaOu
Jpa0zNhOFidKN2wHktUTbNJflYZO+obccXQvxYcRdKrBDnBEEdLmVHXHKnmPvgzG
BFwqFTHhlCzI5FCPnDGJR/l69KoONBjq+No96YbCntHsesyfKQHJ2Gq9OICFqUos
irN7xV2y0aCpj0y6dTILgrazgxytcIztYaUp5RrHrY32nnVsiJHggZkkTgpiB/Mm
YMo150rgG3+KGxOZ5GUvbZFfm1UlGQ5nzlIhLTB/+mJGGH7g7m4Gbe/v/aj0fkjN
qXUJMcjMB7/fjxiAwzdAoh16K6EhQSZ1o04QYHlfwqc7RknkgkzrW5TBKT5D97IL
IfteIJU5P0C20Bn0vU+HpN8bKiS+/8XVliaz/QGxrLHf2HHlsuI3CmQUyYzmyEaO
qBORRhiaS2vfFMtn+t98l1WHVk1JonYuWvHNIwTQDqh9WqWdgG1fFRufCQ3UtBBr
hZ8o85zrmLRUGBfXVuerb/JIEMiy85FhsV0eeWEkNswG7pJr2WPfE+3Idt/K0shI
ibWGdta9CqoXP/o7LYBT9W2Vc0muFLQQtO82cBTKDIAnc49XyNcM2+cQzMxOMbLj
Cg5g6OUdtcoQUqXwEGCxQHnJuQk+VLC/5Tj3FOla6ZvZXp6Y3JQKbL/J1th/QkAN
g844uk7mpmZoTGxX+gb/tZdcdSRMWq4CpUGUJc6PDb/I+hgup76VINNAAq3tn1r2
P51E/yIfxF38Kryladz6dlaIH86MaYCxomwIa5DmpIQufrqkyCJN+rqpLPjXXuJF
x/l7vp25fq2CenfB7e1155AMtNaFRPT63pygABmljF5D22jPqAKj3Bq0iSlKi5c3
vmjyase/Kze952bfXhQMkS+mR9sRsJTqNopek06mg1Ohi7eFcfHmILdSn8DvIBkr
MVaW8tEy4Muxk3C/ygMgAzgdBaLZVLjiGKAjb1ykg3XE98m53CRhpCK3QY6YIZqd
xkf1gs0wIQr4Ly2XfVhZYbXwj0hoYeauMKtp0W/LA7OTRGKKTMStzKkcCq5x0n/e
0aM3TEPdkzswjEZJ1QSGBA6s6Xmqip9HpqXE/x7fEb7p8jO0UON377I1sux7Qk9H
BW+X5kwyOPioOArkl7KcmcirrBXKb0R/Li1aMnWGgrQiVyP1fiKqbjEZ87wpvQ2J
zKN8WGNxOjZemdUYjgT6JYOxwdq2HZsEK7Utzz58V71LjIshcLtrXYRBJ0EHR91l
ewUaZ82pKAHmgtHxDllShsUNHbmRsCGW09s3WbkZktnxjysnN/0nrwLw9GWwjEi9
qAsL7Oi7hMyGEbUhhbyx9u6ZZ44Aw7nSTXUflraxlv+pasXFUw8G6BV8NEOqZy6I
lxAMDrH4XE/tbi37FhYPy7IQc5TPu5pTQT9iPU2n2YtfMko8Z/a3wxOd7lxOGfFF
4c9iOnIglq8UiXsLgDUAqviL7ECxSpRCRcZGou7Sf0XKloJwGRCKdI3ZFuIt/wTW
0pe2a87DcdUtcIlnnQzhOD0m/5Ba/ornQd0IN/p/YpxNlg8g0QGQOvpQCH7oVZBM
VlP+ZHL9C+rBO8dOM+0UmAzGqqyXrbluoX2wGwIjW2Ygur9XrJaooUb6NjN9oWxc
VjIjUDqFIpR/W+CrPIwmivs4hajm9q3ZScIcd711V6a7S2NGGuX0V71C4Q1AFMrk
p2zaNRQK1X/gHKqRu64Mk1b8aYm46SESd/nr6PQ93HFnJWPQtyS2KDNaPGUOjw55
9CFhzzPu+o9xUD+GoF/fBwl9pKAl7bSpgJkFEGxPhTm/wSGWtrs5LWj4Dk06qosh
f4z6OcL02H/l9M9HS4G3vIxf11pGTAzQSzFMoxEydVpRW3s+zXdyUrEE2cDCvWQA
LBlyv3a00MfmpbuVJJq1UxtXzSk7mvVgneYfAakhaa337X/CdJB0mshytyT6fjMP
JcuG7VpTyctrP/9cvww05IdnMqLj2NJE2wthZu9arkFkAiDnM4HJ/nGgKKFMTjEe
BqD+9N8H4v6FW35aOiAaIiI6UeuePDCowwrh0uTjJ96NKepR/VtOJ6FS3WXeo1x3
V961C3+M3nER6/dpVf4/JScH9WxH/wdVlbVE51GkSBvyHWI0VibpTqWEolzElOG/
30WsuQf4B4+ZePPivbXassl7e1i9fmUSc1jTcTJ827sJsVt7ubd60cUcTbsENz/2
TlXzgwN31sSLj1wPLNNq60AxfQqogPrdKh6OViSM8FS2MzhlA4q9N2ok/PAEePYk
ayfj6pEpBaIwy7zjR+P+AccEtMca4M5V8DxLmjbVBKR4pMotNecDBeOfOxafeFvo
8hV8fOcljUF00AR1qXTdfyM+i9nC134+7wwwOB7qWDES/OCgf0haE0RNXrx6n+Mf
vLU72Dk0GUAxVtX0AslQhFT4I4tIzAu2TCIDn1QonX6UzQWZifB+wFFPm31dsc1a
tB+mWuGw/4soKtnzqE4I2RWBkEb1R5npMZLlFc/8I01KwSRtJCdTEnX6GVzHmktd
wibWoL8tmydimljZAGw8QmR7gZHOvfa+PTR3Zi5J8b5NPTCTRuTmdjjFS/91htti
tNX9SAAUeiOaYkpUCwrlvZ7Foe3d6OB2XwU2KAnMO13sgveZbg0l/vB1Vi+jYL1A
TnwU76WLw4SCmc+o7pnnisqqmBIqLGwDmK1/Ris5FV4Ifg9+HPC67hCjGm4cZKyA
PI0IdQCMWKwQXZfF/+/71bcPjBQz6RYVBHXN++sCyvpPntKoXZQMHKRRPJS75oAG
poIkmK/n/ZEvhmvG/VOfBcizU6sJSbj5jSPT/71vdMnVhHRp352BaAoZzbJk3Gve
XgwoHHdR2IXQd9vep+WD36CltJtsn9v8/Ldr/pMDFBC4AhOs4rYOTHiCf8/0U5xu
uikdgPbIryHsuIADjeOIUkdhXXKrv46ryjxatfWWZ1U5OMEKIdP1+CZSmVMB0DRL
frb/uDK18KpWUvyHKlPkTQ5v8c6yPmyrOUFoxxToOfHG/X1z+bglLwzMWpcphDGD
4EB1q8EMZoS3mIgMlz0XhYxRKNzo1pJbfqE0m5x8MpV8uOevvVjqZNCVoqBZAVz7
hQtEEmOkSDXnFSZDDPn1NEfx2wagMThckLUc+6K+4027l0rVUdOrPg1Lg8DOwMHY
0Qut9zxplKt3hzDjQx/Q8PxaQDmJlvnaJLYg3uJJbV89EJGG/4wiH56JTYjxKC01
XsUzwsep6FGZweUIS7zuq6+MD4PlSqAFSHwqj9k1D+8f4czMY3IBeL38WMqosM5q
ZPjs6uVG1T0acQH2cmJZ7geW/LGT8Bn6ISgOXNjL8NyFQqz7euLLhKEdcN/JnVKo
xPBZjbxhW/QZP0KoW3tyezzqCkxtWXC468a2ymaiI+4jkQRGSGP0rPLhSXpt09Ex
Li2OPtRMPWHAaw5dPaCFVAoAzud156j7xviqTwW5c7GmxeBkWGmeLpX5/KQFTz35
fflg0sdvtxTwwBi1X1hCp5ebzwub28CxlcJvwhqnD3b947xYr645T7M2fqdEr7bA
exKObvy69yTlyDGvNE0BtU2nVp6xuQjIrr+0I+q+qNlp93MbOpm5d/XApH7Xomna
sD845RLVweCewJ+I9XVXuk0L5lpQBRmWSlew1KamYHNL2pGxZUVTwXUCcK5jVOBw
fGBdoTTtKsOWjy6DXPJnKMm19NL0jMHdGzmOuzMjQJvfE8hOChv3GiDVOG4z+0pP
IBDEx5LTkQXB8/HD03+zQ5PY8nY+3Kmhvo6n1eHWQOEDcUhyG8vno6NtqfdEVp7y
Z2NaDFIAumJ+lVh7KZ7dPFalqRDKflKXvlqMH70UcgR/wKaM/AKikvgdXOLaI5Gp
Yp4xNBq9le3edTvPA3xJVMK07maz5zdZNt+isXTCiCuxyP70Dq4xpV3wQHQNdXQF
fWy68Ba7Ck6W428y9xUdWH3FYpovtVZW9Kr7ommVl3RqHPgN9I4DfLZtD3zyT/AR
hFSVjDIuD9EBY0xTV0hw/lyf2EALeLHDC9ic9wXmhFso+4k5/wa4Ru2K3Gg2cyB/
l2t6DxI2V58tWZy802fyEgTsRMHZqUdjOguOGEnjW0JbamLV7PW0lHZQy3Cv+BfI
gLyads2bEdI7LQDsGLynVp/rHa005hNz375bUKXGomBiIvyFv6AaZeXzwPSfxCve
orDbby/vMCuWjv7Q62s+rlYmijEx/NEoYpipaszaFeb36mbDhpskIfY7bx9Aimrg
GGfHSUAmHThu55NNGtWSyB1J5u0+yQ+iXrtZobzWorwClGsLYGgcPxTGME7/w3u5
033DssP+WjUB4VoQh/3nW/4Cfk+4ChFuGaY7OAF9SI8kmocLMDyUDN7vI4R0Y7yX
iHnm7sRRYGvc+Ws4/vtCy9eTkEIjPqmlSys+xYKMNDe1wE/k7s3OmQVfsGi07DkO
avXVXvUJhO6LcvdGAVLncYdldElhj0bxR03uXBCHLHoWl9xMMzl75YuccPJRNWxO
mmOvj3yt5v+P99cLYYnKt2RiSS/q5Pdg+KjRfMXsnDNX44xK/mOsZK7h49fC90lu
3rkuQ9+h2yvfhMZOD47mxyrL57rrv7VLT7bETNKFuTFmKbbY/1vVXajWbMKWLU6T
fiAl8jM6eelZaz2mXJqZ2yM9M7UgfTSSSr7obFrWe5AZiiGHIHGAgqJ8c2T5AChe
eikop5oggCNfUw3vhGbWG3yHzZd4av4ZUOEeCJ5CdpD8anOu08eYhrih5S9uDLDS
rOEWHBCd+bgpKPJ+r9PUbzBo83F9QLivT4D25f91EKi5z4wwT2TdCqsChuixc8Bp
WsSX2D+eKNOZAKMizrxWDhNkFcJZXs31QoDY25GTx3Px7HRoJ4FvYr4Qu7Vss14o
b2MQJ+lqJXSnQCnaqAH69IF+rQczfaIF4F8IffOFwJFsJMzMX1Cr7coSgTuHzuQJ
A+p4OMslL4zpiJ9kRp0UC+ZtbwdVaD7zGHFxjAHkPthxMOtJxA0u5L33FcwDXZvW
smi2ZLc3yZXBoIAv7r04c+ePQkjqeBtr17L+2sqQ8/WcT2FJ29SpitD+W7HVjV1B
OU5gzU/Mq9/Q9C3i4Bf+kcirCeWrv5Bwt8Zhf4WrD/h/4nL450ooRo683SYL9zqr
yuY2QhYiksD4p1sgSxMZ05D8wULL4ig/IclAJREtO1mu5A0TR8Tv0K15YP6ez4wz
juc4WqnxL8Fuzc7hgHs366nedpUEkAI4Wiktx5hrT8oN3t8ZsWpwXZF+0ou8Mhtb
7gYZKimfgQ1Yqvfny1pv120lJeBRl5lDWqTSjFk0elmifpQhJ7LF0bvZxb0Cgb55
BBgOVI+bYHo5w356uPlp6osVuMQEZl4B5xyH9GzYJBxbhD09u7xplYAIQimOSKio
UekLxBdHVP7rSeui+pQchGtO3fKPDiXlIfoIdL6TttjGvdIHBCIkYhm4rGAZ1/c1
Axtbuqad2YKj0bjezbIVgGfOWAJxUK0q0Zf7XSi+pEkoFdlHVo8hlwlDfNRVeCzD
NtWSXF3lJ3ParaoThfPUoWUC4Us72+1qwLHI/SSrh9gLQix0t9o8kDVN//HJv2ny
Y5yajVB0gjIdAjC/V3VW7szfxgbI/XCSggGyDNdNgJuipjZ3b79QwgK+NgQZ7MM4
VjCUqUK/3VdT9z5IH1TNsu2wKDdYU7JhyBF7bx6c9T1DmSd8v27snIGGBgysRO3A
4O/E0InMdyHYeL7V+U3SvA7Ow4KW0hMztfBpe85BYxoMKqUUeZtCsqRnqbIsVEYi
+P5ID3cbztGaY4rP90dDLIZBVs8Gedek7ae7vh5g6K2joNKVFCxe2aIxkN0Efln1
QIz9em4ZRQRwrhmZlmJlVCdRBJTz/Du7dDJy5UcNYw7Jrt5YthqW7frU+Pejyigv
Ju+BaJsV3trChZO4iXbJVnhgL9LyTuT8wKTXPNd56XrI4HIGune3Pt9rFGcKOyqI
RsXHIwEUHS9pP2/9PpX5vRl4DgdZu+EYapFbb6T/pb7f0ljIMF/NZwM0Dm8c4bwP
Qm5NM42AhckdRjniI47ZVdC0C7iR8hQ0Yt068aP0Lx/JfkzOPwMp7aL9CfTGGrUU
fSPbJYBqon8GiOfd+xPgLsSqI9DlO3p6zg8deNJrkVU88saC2ag+1rtRrDWUIuln
TH9JnrUBlQEbdhJ8E+8JDHb+NK+GUxeCTPufWjqgdVKlwLT7iigqAG6FHc6NlEPT
YOs83PGFm4wF8X1IO/ksF0h0asJN8gzLRPZs8DQMQnj0W+N9Df2SAZEQgMXyM6EW
jyA72v66LfAh0Pd8+Jpt3ASG72iDfPozLXeEtR9r/AwsHjlhFBPU5hl+fRHOyodm
5JiUCIHk7FgeVRRVaDD07o/se4FmV7NlILjxFeWBk7a2VLTLke/4HG8v4rzf5Rgj
gKemFsacMVFnUrJr0Ef6iQ5DeJHmIMdi4JdZEWoQviP3xK+0opS8EMwyMu5VdPqB
cRXAdFVgl6DPk6DLHjd/37uzwAfoJ+9VRXhtO+Z43/GtwKun18nqfEhFXXoM1A2t
BjaVFdf9QTPYEgTuM27JzFoHjI8M+PTPFB3quDd0jCZnYNE18Vg9aW3/P1mDlkh6
KTH4lElRTfj7Ua+V84IaL6QPiFQ2PRsHeKNU+yJ7cMYCKvuY3FEKY19euY2waz1p
Pwn5Y9khZdZUEPmNXsbhTcE2dnCZXIh8laLV4+0VAZGygXuWWUJ5V2elkr5fMZ94
wRXPckaeFtuy6ccurE0n7XmaiOwdJCKVG7gtw0ikFCDgwV5GFDMOO8pAv1oe/bhH
fokaL2JBXD29PBdxh0jhQ4vYpGLPr7S+BJl1F5bhx63ashyFvitvJnNysUFmgfse
Y398o1trUjCZhfl5fk0pf9mE5TN/zT0YDLyAo/qQbbbA31qRX6LN+ULKriPumdl+
RoeqEdwzJYTRE/kjTYjbHdiwJyxC4hDNK4fAutmx1thwJnuG9dWC9B422XXs8GKM
ua2SbpDyiN9wohfC3X7hcnVh3dFmHF6hG+XBWPTs93QWwq2jwWYQW5m1621UlgxC
ZYYLpH5acMl12KW9EL81TzFk7nzQcP2VKq2xYLXkCDpS0+snGo41SlyDDIFegu1j
esTCGmptf5JWTPI+b0BG0Vsut3i0u+YyuZvpixfuTF4T/YF0bWvKVfmCUHPvHLGa
xpT3ekvsJZaK/S8GE7K7tWIGH0s/VkkXEHGYJoawwbhrLeBrg0kcZii1BOxuVVja
NPyIFubY9nfvzOlW9qPuAAJ33r/VOSB0sN5RaPncv+YZ7OY9JhYKds6IQ48e1V/7
yA+RQV/GZjAI4kqeI3+kqM1LJyUBcLpheh3NUWZo/ZjQyaysHZ/YNGRV4rXt2R7A
mpiRIlaQMTXLJ7XC58C7jS3TARvI1s2ue6etT2PaQpOnNh0JdTo43j62xWUppehz
xUuL8EPbat4b+XJtN3Rgnl+AHFd8jP/bfV7eaXx+5yoE1rLXTsv4g6yCpXDZCTzK
qdJPHmFHVDbBd2EFMhSlISyRnjgWW7Zh7/MS1n2NdksMOJzk6Vy1nsL3RFYdzCyh
iaNNU4EYuhQH7qVK/34Z+JJRxeeNzIF1Cct+Y5lq/NExnFyyDW3CoOa+DuAtMvEt
L/RzlW5bBOCMd2cV1C0BrxW8yOZ0MvktYyyT9ddpFCImBzlBi62jvjEuuY7LbyBV
1Evh9KbbLSocH5KI7crSankz+2xSPkBmyOCTjVMjSV7izBGe7gC1BW8QHnRDVUAD
NFFvWt2I5fYB3mfxOErs15fdDaNQxyWa9Qdoyx9OxLvGeS9SeaBVMkSLnQGlTB34
rMz7m8s6gU1xhAZoMGZseSwSiGFtgSnFAjDnDnTQSxQb8tjh2kIKYe/RQjYZxMMQ
NAXcm4LPn3mpvJLiObe2NWFOBPgAPqm5KgxsxMg5MggBD6IQHuQUqI7hD9uDdpEW
A/gykxtTJq56OK6hminv/gWXoucz+iIFBBVDyxAxVI6HY3siczXAiasxR31VCePg
if4JsPJB0pxgus0MXGQchgnUI3QnT17FVDumWis7jNnELCeoT9eP/MIAj5v8Ikbt
/UDH9K/83vodjOBiRxnMeSRtYAmYQ/jZlklcEP6DKAUSrWiAUtbe6l7Qdax1yK8L
80ajDL0lbtidXBUUh0CrT9c5vwQ+0DjWnD56TlDpl6KGIafHbAyJnEL5TDMzgl5U
jZE/9IFRYefvotwxdpMp1xacvEbYNH0tims1CGysauSHKWdURjDHDOL9F81153ga
//PbGCZLfEecRjQ/Ye1PY9yR5t+pTklGzFmx6bUOo+DkD0+EHNsxLfgmmy58e4qa
96b3cMuD0s7PnWvX+KXYg9BNDtJYzIESULZWT292zSKxU9no14I/4wnHLM/CCeut
hew2Dm+HJ78FoL4AbM1OhqqKQSoLGLIcNUD5Brbw0LS9mKQWx0c3H6c+06LAmZw+
rOsCCcB/HMnDIEsaIYO7Bqllm6nJ92NLLX+0uMt4YTSoLFcjE7yRo4SFjobfrFYm
YeRL0BXBjVDET5y0TaDgqT2a3jdBv3pBhanhbSth1o6QQ2jMRWmWMXX9Kt6xi3fA
fro0VssAwS3JN02reYqCFcC6Sf8GShqSbMbjcfAZCwzhX1qSI8J8dK6O/FC47Mje
fO/2KqaM7xOUuPRzG2zy7Tzdda5f4FP8ovVIXLYb93DSB1j0mJWq3lf1FAihJoNs
4Ogb2czH58skUKvri24jBQLFG3Hf28SwbmoaFjZqtptYXtsJUjA9iAdWs8f4ZLqp
P9OG6UCnMe/JJZP7b1TnkXBQRQ+AMTFjK7viWycXgr8fB2Si0YbAJxNbFBjbYECb
HyHi3zgyd+J+bm9z2vnFEIMC8H5GkhUDwLPG8b0JhKrtCOuXME8ojeCfpGYeKBpF
2xvxO02aoMl/AvDRc9O6x957+ntlEMHtRiuFwbnkRLAbUlyie/3KZiuT7DvDPFxy
mvQXnJ2dWV7a1MFKyjOYXQ0EI8ZomoJJMDWXk1RtVGxeDHCO+1OowthnXXoxermw
SvzXIlxJ68OcN1VRblxSCaG6KWknJ9wXBxTu6bgWORnXK6uSAHi2DJ5+tFWV67DW
yyvxW2czZJ9sHylSCvABeIfH14gLC+u6lAvsOCq3kZfX9lo+ZGH98ipj4iYTc2Pq
gbRPxBdf8iqTLUHh+gHZ6e5cFefTR6TYz5PVK+2OHuHh9JbYrBieW47YWSQQu6VX
0ptGKwR5aTjoId25lh6WjpVwIX5zSRUgf6Lwbd/x2akQ5VypP4iRa2gVf6LlXoXX
rASqtoC/0U61FcgXohNdafjOaEX6utqQYh3blQwB6eqHiR6Yc0FumKHyutZKmRAg
1ebwWwMyH9Elw3QY4OqeE54YpkaP55lBTin/FToZYGYVxmpDuGenbY4Rn8CVDvy7
JiKW6SMQ5USs/4MdUtUFKIn1urPUTWjOLw8l+qk+H+xH8wE9y5xNBhEH/ivj2zbR
HOLXd1PE0MaW46p63KWZCncuICmIweIdKEqsaRuFUvy/53klEAbTxg4L0yR5Yve+
tjTl0BRODxds0qidD8tBghSoxzW00X5diIylAMAi1WLj7mUNlcZQCD6c9azT1pTB
2m7oRMYUHHdBQ0EMeGcbTGEc9hTCBjdV7BtgGTM1SeZSAhGwGOpo4W+U64HavagH
YzZ0JoFe4FzCbuYrkZuTYRKCqHmi2Q8vTgB3EVh4XH2K09TuMlvmkVAYyXX1lOrz
m7YB72stYriWSsAAmJoYt44UJmh3fycLH62hcoMoD9K2RkHJrjt9gGFNg4rLyEfw
nS4pcCnCdGR1s4yxLSB5oT1ceZaVyqSWPMHfuyPZfZR+xrMKbqhivUjUB2xl60gN
NQGSQiJ9f7LDMGt7gsCYsP0VDCziknHPUMOIkPj0o5wWOtUrJ4YasKJVtqbYb/pS
izsID3YmGlF4k1bZmiuoL3IkSuWl/1ivBgPbSGe+R+luXs8x+Y5uHQzzzY1IFekh
lSZb127Cy0M3wwpeWehGX38s1mhKP/i+//mbGE6CB34D2guwcWR0TLo7ZpXknriY
SDrRKnvbb/tl/eO/bkjP2KZ8dOu59xkBto7OKNkzpY9ytFKKxvUX5uX8Fy7wmZ8v
/LhLbqaPLeLbU/yE8AHO5FPTyflmgaKdLNEQEUEkshr5XZKS6gh+dEujH+zIlxJw
Vzaj1bDOKd4WTQr3lCITcoH1gVzlhonYn6R3cEqhIh3FVqv6wv3tj8f4bAiPsdP8
T3uDEChjzJXgSXWFOK4PsHRuQ5p5ZIsU+GvwEh6VU9OmqRiwEEWTqzdknMvL6ytw
T6jOYbLYTUrK8lrqinuaYq4sqP5ZyNZO8d+5RPLcPC5a3I2VnlsJjGYY+NfiPMX1
5e/pS7krMvC8GDq7KiIr60CP5ioDs5dmEOg2THXNaPEZwZIZWDR8j0J9w6mRbiaX
zz47YIt+KKrXOiw6PkheEH9t0SGGBWDESht6aBtmWQBsBC+55RfKj0KKXwbXV9QL
EmPYm17Vf1uCa76XkL6mkJMgOx7ySbYHNlXskD3jZCDfqY8++VOjOgR0PKitHbXh
KbO2n8hONgcvU/ToyPAAMngdWcI90QyfZNQdGpuU/9Dp7RRR+BypMSBcAP1FRir0
5ZOYW/TjV8/H0pp07n7+BnMFXLofjz574NlcwhvrkJm6R+bdgEC13s2kxZZKCVRt
5/hTZpSsAknG7SvKqYT3ogkAF5u61UHbH8a8SNNJPejlBL/c1xclGUgBIJX7emoH
Ya0kIXjvBRUNc6CfKR+gQ7SA+zYcfOB1WiL8fVOEn6UC54RYDuKx2FBzxOXbxfRt
hPxbVCVGZCfX99WnSEduZJIKzEAuW4qeodEyPUXZeDc2nIIxhfmMZYhr6TpOHDsk
yQf7RyGBzodJpZee1lC+TA8jre1OfXRO4weGXv7KPsz9LhK0hzI5Zl+0ZLekvscO
01/OR9nZw8gUNY1SP4NeiXIp+M9Epa+dVpY/BslM+dCU4LX4W27jlinp4CmNrXxl
SAmUDIcnbCxuATUeAtZSdYg+J9dODk2mfm7dwwlLQcQOF55deyis7BMFLJRbqMgb
SB1EJuQ9P0pZLCrsfSOzmi4qjAVp3BEw95jIc/2jeRM7UqvVTmauXi0Ntr1bZS1c
uxf6HshMmE96WmtdHms1lR0FHO96cWrUQfqClW8JUwQuTs6k7b+ebZ2d/wLVSXoj
y6SAIkcTI/OoDAp/V9ermVcdMle95yXpd/Z1QUfkQmIbCJaUJ9hI0UEe33lIQNYV
Poc3VnjWz22wTdMyDQvugKWAU2kQt8tTqf4LzpCqnGIkproVGxqeqXVMgyTkoRkd
Q+4lz9lf+C2KcSzmiY9z2+CBGt14ao+FlkX1zaOqoFxnrkwrgWmq2zP4uwznZ6wo
WuC/9Kh+mMIro+rOwW7UbMaa3kDRpTFB9m8gTQMR2fhzieLzIUXnHFns2p38/ExY
E68iu4dwj4CykW/f/1N9hrU0Qe4hjnImb4ZI+S1zixKPSR50Nz3K9ra9fwtJDdVj
XU4YBpyZ3oeU0czJei7XzPWpV41Buz42b5tUwn01u/NEjGuPJOfDTdi3SL34w6f/
By7bQrEu1SKNrnKUORacaJOU5npZSOhmPAYVbaYI1e1xyS5u90Ly2QXj2COfVDeI
z3qtFbu3EV4VjOD4Q0da/1jq8cYELYZKpkHJHbV6HPty1AolA8ysy24FwYFasEcj
2RKkzoSbDCBHifSi+sneI/e33jEHvExIlGvmhi9U7AUcPNUdbzqNc+dr3BBuPN4O
DbhCn+Ftd5A30nHwAA+I954zpit6AFHFv+8rSKAYsIEhqlgh5hQl6StuCXN5vJth
gDlTa46DrgWSZG2MXBLv8QQruKHfSgZ7O4Z0B9oP0OMw3Yc9lc4b0rjSu9fqxi1v
b4hac2MJ0j2N5bF3ctwediI2t2m5egk3qbUlpr2MTR+rkah7Os7GbZMO3eMAcxLt
Dt0+c9SNuOBMM4jctlcQ7AB3P6MXLliwdOz+VSQy3qmxjbPa6Kgcy20sfxmOD48n
pmO7wCAhwr8UAYUYNtG37bjM3Ezew0mLpv+/572L4Nbo3k3gVbLRmhzlkWjWOWBX
QFYI9t5mrbiaTSfydcS82+XU5wqb+We+6V9eoRZ7jtT7OQXNu+n917T/9ejmrYjv
IMvwP3t9CsCOOksGtN0FEZK7yuLpgyMeFJt50QkUifd5rkR3wssU0ERUeuU2c5gH
zKM+f6O7/IZxtutIZ5W2GmpfC1ApI/NrkGAUJf2HthVomb/MFW2gjrRv5E3wPc0G
XrnO0/5PzjwKAnU7n4+McVHpIakKujgK7iN+7vihdARco4LNVotI3TO/gkixWFJZ
tBg5DqRr2LgFG7LjpTgIsAlSZesEuO3vWGVC7/vmH2u19gkZMcbWF+FVvWuSWRTp
JonM3uVEdnHc8At75/ZdzERjATU78RZEfkmxQTH0p30Css9C9yFS25wnBcjjycyc
Ea3xF86H9egTPzjVdJgzu45E64FyKviTUO4e64x4cg4Q4mkGSnPGtHc7Ko24Lv4f
6Hhe5PLWne6lUXEmhraS4F4fQdDdwakPrhkgDg3zsiktzdF0TajN9MmiGwuBuX7E
OJcsjeIFsiCwNxmC1VByr017ocWit1I9MgXC5NR3+8p4xPbLBc0QocsXJoQbTgtH
wSMrX0/MArFEPJ7IKdHQSCDBf5/XSiWilQo3aszApvc7NiCtDvvxcsyrbKL/0PFq
h0DAvfZaEV56/PGJ3/HurYKAj+AvDZ2MvWVKmu5m1iKu80RrL9w50ex5jU6u2olS
qJbjUVgQutckRq5NOnklFzLe7E8r/YYh3JdGTATFdPXwYqoK/Wj0pxW3kCsfM5rZ
i3zh+6tfmL1m75M1x1kfYzPXi8dx0G5STQtTW007kzNCg+FPYL9KZkXUR7YSPXv7
xNqAGuC6czuwxyCWocuSJ1+bFdSqTgmL1AkFn2NV2jZKAeh1OUkBE7LcReToVERw
9Otx3hVqrsj+a2/CY5JBTUiYwaAqInSm2Cb5tDHm2fIBNW7Vv6/m969sJ2b4JMhg
CuwW9sPinrLIszVZX0qxP0Qitgb1cZZ3pQx/70OjQfjFC5KF99vnlGl7sdLrAL0v
8nd6zldVAZg4KWI4LTOwY7ATnyz/LwGews/qpKxHb3e3kV1t5BUqEnaCs0rE5J5x
7rvl+Y5wcdpyDILriM5dUgStBUBX4YHVVeg8+/9bdm6CLgBplzQFc1mrksfAIQSd
ja1pAjxwMXCyGSthFAvbQB9GgDS9+Q01/5Rom667AmZtZ+ndJmaxN26N5yvnNR7H
Hoz/t+Pc2UPcqoTe12ZyAJnYo0rDppLmr7CqhA/ocL6hM4PbV6565sE2GalnaYPq
1A1ff6DyIJ4ObVoIgJdexoPg+EUhgODwHQ2YoE9qrKHRuaopW6HFuM3E5LO2owTn
WmeGENjGlQ/a7AR05AEigrCPAmOIJA4zKpOonf55qyOrW00oMaV+UsYTC4J4ou/Q
9Vny3rkN0pRaLlwQ0itdfHhIsTEdGnrlpF+AW8VI/0zQoF6DtYmku6hTzr1hCLHi
DwfZynIwm730D8MxEwvqmCHoAXqO53xgSxxi0bElhpjLPHHTBAKTR1x+WktoZOpM
UskqtAfds5mCKjcpOLLK1PDyC1X4CwswkAPEfbc3uoFzipkWuuceVNibuMr0dUpX
NKmSsfJTrjtxRYkPe1Tjalc5MgF3eCmMfF6Son8Bn58Cg9FbhRhSCR5wa88N+hRX
DMwJZMHnBXAX8onxdm1gGm2Zj70Si6s3BrMs2wJaCC9sI+VTvdOAJTd6/NpPXxRy
aHBMuKgoxG+uluiVDJ36DODB55vCGuSO2TbW0kdVhgMOM5i3wzC6GvAJFPtGEZsv
u0PEmRFMcGvvT7WeLOFcu2Y30VOyxc/NUoG3BbMeGnYxwnnnMwZddC1f8Gvv23iO
p/iYDM7tNmcjFC+HaZrMUl+BMf9LPF7bUaibUMitSSwxxcEGc4q/C3213Rz1nAcz
dhGKg5k4/MuMfkZ/kj3YfepVUn++DRUkd4NQ0xy0yYZoS05pIm6Rxe2SRGNqGdyK
WTE8cuc26eF74U08+JXSqgFZERVCSd9fdw8uGRlwmE4w+vo+UC1Bl7ZMHygXN+FH
PvebyQi8P/hHZkHvGgCkvFcat5PGiWjTVTcH5O/goiMWMdqSmPbvG6UNeyYzHZTM
qNYP4Sv+zlX0t4vkDGqEPMBK/yzRHacwnsuJK6qeSA9EoqpY/9crYUNPVkZCfiW0
fDPHphxuztKH8thy3vHqLWkbPHKFhPG3zVDZ3OzZp1TXi3w9C0c49HjS8xSZbRn0
Py/dDVd15b3gL9uA4BLsEUMVzB68nrsWxSaH/Gy4GVX73ibexBnNw49pl3kb/POP
nGOrmTy6aCyQ7Roub9mlClMgp5VJGeW+55zHRahsVQldhTSnHIVICKcXHj6HQ7t2
NqHAMoyCOaIJ97SnXS6+tSd4Neb97aNwaUUDR9Ml7O0VPajJXliXVjSWP64Cysn0
QRuH3A5DWBsOPBV6oT1V2aft9Y5xWrFDWihXiuO3Zz9jot4qMhDKDiTwFqsqY7Ov
kt80APCmU8mS5rg1DdOP+4SJ0kZBSnhHxEWzKQP+V225Ip16c52PdatLG/ZreOMO
+MRSDC4ALWb1AuQal13ghJv1dcgskwkAs6S6ZufJq6PLd5A8jpgzDqkXwE/1VENv
tjmG6llyi5ae8SOxZIr8nWopqhkW03w/PjXVjBKiv7NrAG+9lnVW+GQIqF1X0n4l
0HHODyQLrq84ay756ONx4YAftwmiiXdePjOxOudCZsg21FHvEGRKtkY24X6/PmRd
6hCOp/8n61NO4oQihLPVyY5tQC0XNDliqiN+MAW7IHaKpmhIyeCSu6gN6LNycS6U
/edpUgurcV/UqdHxGc2/QrV9pGJhelGP062kgGu53GgLM34i6w8eGS8m0qw/a3cw
eZvafGvsDpkVw3aRbAonzw4lweHa1IGAN+qPRf0yTtZbJRpMP0AFnwgvzosJ9VXm
bMkPDBC02FKSCAIbiTsnwFrYcERW/J9Wjb4LMmYDwx2JyIO+Obau6mUBm2mE/LvV
Rwa8LNqvob6Z3rog2MsMH9MmnWjRpYK2TWFHNyOViONsAPLsnwit3ri/y/q3TnBD
IblAiYWphPmHVTwMG3c3EHnxmdQ86UgAfoqHescn/uVeRkQSHKSBJr6cqvDb8vPx
YXTU86LoKdmrTNM69ewxKechXNkoynrveP8eW9Gl3/W2Xa6KHMTnot0BNRpdZHI7
QTYBlo8nX138dP3xDRsxz0LXPfmAeJNg2BB117IdNt4O/36IDqXhi2PI4q5V0Pir
ovtF5ygYTMR+1OT8OWDSEAMAb/0BugqRyg6Z3HNsJGjoHAlAjvgTywB0vmuyiGOW
+9OH9ymVS5dt6vdHcJspObOc0xlD30rs/Npe0mBr3FOM8zTHLZXCLbbVrYZvIq2L
DnuNWuf3dRAfuMhpykIbwI2J4AzqstvVehk5zeXHuzpCdFJJskQEbBNHkz7j7eDp
ztYTe8zYH6l7yvQOhwjanhqtHR98+WVKUsP84TtBkE3b+WWELiXIWqMPpMp0nbxd
Pj93gQTDL0mDOkux41nkOqr746wtnWBtkVpznb/agY4dNmM+Ustx2QC+SJcAlBwq
Zx5xFkKrdcd+kdqG8hz2qNLL0o5LNuALKNjR+sv1Ab9Dwwt7C8C/R7NLQUq+suTU
3dI1FobpVDoc9316OckCYR+nC+def1Sc9wDHpwZoINaQKEHfGluom0sPN+IUe9oW
nIMJd1jJxR/cu9sOdJ9WBOGUaJyEw2utNsSUmdHaLH+LyBG2EW8FUdnieIbxbhfj
9FSoP/s6wHBTweQGP5lQLiUOi41842cvUK5R2XAcOZxi/qWYf32HSpCw0E+fd5PW
WWRcW7GpDzegEWc2B1+sHM1MuvBKG2CY4HYLG6TYRL4Q7ReWFRMJPIX0VUTnmSQD
XoaEykOGnWsk1g4ezRUwU6AO8zDs64Ta3YdlgS6xZbGhVujfRLzBVqTVN03n+HNB
T76+VrWtVhAbmZu9RYnRVm1sxDJbBYwgLu6mD4GO+t9YF/r/uLqmHn4XgAk8/uit
zoeWDlF2EW/qRDF5DvSrrNQ1p7wOvvS50tCk/UjGvUuwoUSOcKvYJXCJ4DXSFbZM
+De5VAp0llMwDjuC3382EAhdkIkzgES195TH04aIqjg/L4utcuCoCf4ln1JSocw7
3s2xuxCrEQZDP8FppxW4rSWnwcVLUWlg1khfnoCzUJHECpU7OjV40Kkrt+q1H/Ou
C/aZgjTAaAD6M4A25tkPxMa0XMKRmKSbA59HpssrGyxUQa52UBqgbZNX/n+20XOj
P2KRR19htBAu8cvy6vKDZ6wj9+nPbYvx+KMsf1DbeeRTqNJtjv1A3FZyUCAwA8Hd
so4z1gejdyCiQFtrn5by+iOXsWg+WypTG1VlI/gO2VJRuXACXih8XKceEJi2zwpk
02YxtqrUx+DA19BPx5LVb8LPQIVY/bRl6qivsaxOXUEfwqvyqgfOcwYXUziaGypX
cWF1iD0Rh7T6EqiHKlPG5PTzpcsldsoKcUYvU7IwTQB8jfQ5TbVvplEFs9fSCC4B
6D0O5ejS28Dx304p398E99gyDHgdvlDQY16WYk7Z5PKei2lUcSgi+K1eOCnCy+7L
AE7bTukL4xbIqy40lflppO8ZJuR9fHBf7yqn86bIPwlvngcZ3ZBJVpGUKvEHuahk
TSmxkRN1sxoweHOQufqyQt4X9lrvnDg/AiQ7fu9MLE6T1sg1c72F26tC40hhUfvC
8BypZ2IMBd5gklczL0//+cmxQlYzshH6Vf5DBKXZ+v0itCmS14nS7T0T5J1EyDoQ
m2X2JTrQF5MEEOY+aCkUhi3G4HfJDT57U3P+ySCgTpmjNnNiAtBdYx5yDu+1SPck
wWte+qOvBq2fMqywdFYwqWzOLxJC1VKuUgTNYIZqwik3dVow7q/2Uhfely/8oIj3
9dw6GGd5f5yYg+z4LOReIHBGSqf+zM+Ao7tqfJUiacdb//1g4/rKV1bHrKHhF92I
ODDxwkl10Q0iSwUQk6IMnzWXA/CSr0+yA9PGnmFQOwVermV2uQhrFNNERVeG+Qww
5zlGFNRgYU8zE7KhiyW447nrjCHdJ5JjTaigueybOsY4B+EQyyYgUQ2Y2gEGKgxF
HtbxzQC7ByGqD31whHr1u0fmrFzyFt1cxAyJWU6MmPsERA5nonRULo2Xy0LKnIkT
19WjwgALSb8b7mUQnNDev8VE4N38JnbbLUbmntpSIfhmr7fRiHQh5YIhMgnn7N4L
SdK338wwKP8vNlg5wfrM1KdtMuUNMu6FMGfYudkyAvOiy5OBAJw37srmx4q9uo+c
eO/D+Wkrw59xtAgc0MS+tyDe5Si4XxfOqfCYWQAaBa5XkrbxtaJbCvmK7QSlQXtv
pNZCSbgFfdyTLLf+UjxZt+f/iK7rbK7YG41V9yg4T3wQyV8gKsFLz9hGn4zsMiwT
5HLN3r29cEsNa3DC4JoMIwzZBcXyLkH7kz32Q3I1q+QwtLwPiwCWN19adcp8iR96
3ZyrUOm2i0FZMqfQpVPV5omnoNng9PugulbB3XM9Btf7Meq8595DzsJoXLm1qqwk
iYdjRmhPA5iZfziKOusxb7Vp5kAX0Dnsq/IZxKYk+PPCJ9AovgiN+KEkoOA9qn2J
j557ruhSZn256TcIlN4t5On+AxPfCNKsRPNF+LmmFbf20Leir2PxYOn8bmyB37dG
FQnKuqyHjMo28nxgQxD3MZ9GLS8GiaunB2VgwJzAyiqjvme+zO4CFuJzeE8iKUMf
ON0nII7L1ojYWUXRAW/bDdfXiS2ih0ur1yJXEKfKYcFzGcE06ZPJW1/yoUJXpSet
FJPYipd+SSdACdlDnaUgMOfqDNrLR4MkxTu1ZWbWs7M15HP/vILHoaTlPHfWy4Qp
2pD3wgn4oOgbCaDQQy5uFK8F4hlT+DOIOb9gpxSBvFhN6BEqsosCiG3gL/3BAQQo
vIYD+tEy3ytHHPRsmlJVSDLQeDqC7vAmiaUBjNdVs6w6UD0lzgU1t1uwfSQhoCb7
/UXBXYt0HpaK2SAgitWCPiXIXK79l9hxR6snKMQRcMRIr/yqwHlU+kCH4yzFWzkO
QC/Mis5i+YUWS7UBz5RduZ/db/nb787gbnKT9Ue9Dpokq0TZi5PhwCKuBkHPPb28
AnBZb2zG38joCs2TPUzcfpRgZMrIPvh1nq0sBdVuoDCcto9siXFuH7wCCKchu3FR
toO1u+zXEuPtFJTJlXL5rEMq73aFau91XB+Ln+Zl7+M9Z+aBSwWD80DftyXMKovd
AZKZVNLqFsE6F4jvg9KaRD5F2fIf2zPj616w20mubfYkIW7Wj670Y8t7nVcR6vk6
9J/ORu5+eGBeNensIFSdVq73kD1fKbbF8MTGgWLEJIsU7+qR0M+ZIX4FU2P/JhR1
Sb5r/OeW9ragfQejHi5gJEwW3j6141woXRCfyxTGsEH6mYo4duXiNCMjVq1BhFGp
dJW7QuIw4lVqwoSzrLu0M1/DrSpM+I87gdM8TZ6/83JRdqNfberVay9uIvUnNiwm
iQCSSM5skZ3RCBQjSNZyJ3QtYdkBYJCMc1CMy8myOnz17xeTkhBiyVPBdPSITvNN
Y7rZVf9j+K/LZRHQurhTiu6PFP2uXaJopDnCIIpitTfEHOxSIfJbZlshWBoCBWRV
xPSAYoVcxumBDCm1m5nO6lG3QySYgToOVAO105niejw7KVgkCeRL03wrIwZ2470n
gonpAHuQtz/azwqwbsr/glgp69lbPqOf6/evakojxe2gROkK+WcB9wU5yfVQ72OJ
/qGyVEYu1w2Q5mfocAe7yoEq0vCRrIuyXfn6rj4JK7xYpCa5CAiYi1Yv1Z+kFzQO
9XzI1kl8NWUD+6hB/JZsc6xEI8v1EaWXBlkBpI6CMVXSfJ0pcMi85gJlE01BfiNS
CWf5MBGuc3JDouBIl3X7VEVK9C/L5LVbNpknTCj4fdLup8VA5dxwImtIv4uC+IH7
0Z2XuwRI10Y717Y72+tqc3yGeeM49DISq2Sq2JgR5RFupMUiO8v/N5vSrACThbTF
7eTHgTGUuClyNz1jFrkHRkgEuYDWywjuBblm7Z3MEYNRo8XpinU6nqvzdtAXNf2o
JcItSEyA/hExAWoX0KTf/zG1QyBT+DNWkRjYLiICkXPhsM0SeWqbbTZQKSJhogVo
ICNoVaQAKxcujX2V/1SjHThnWNojwxrago5vczeImXUtWVlcjjNrwAt0uxqqH5Th
X+jlixD0mriOmfVNyLWKISPXjw60/dbZVqw/a1oqfTiucEjCQD3EGKa3ZBLnoRLZ
fJZOb1e84qMVEgIgg0ECb68zZuj/YdGdIuR1GZSBC+eZEy2fwfSEloQZGVbt6G1K
I23+fQl21LFsXsntmT1HJVdnX2aroQwENBQYjznNJaxb8ENavQmo/52S2Z9Amc3x
H0UC6eNdJgdLCYtZzIBCnj47BlpBtGxO6STTo2+Tc8tTcZ4ca2dM/YumMWfo2LhX
ZRiZV0lQBdG4rSmjXdjLb56ldGL408rApYFFNezA6UPesWQZShQjCnkU1L+AVxMz
Udgw9xwbCvDLhApacHbrrkcEPEtTv1bCWUQevN1k/BlXBMYo6gOt0wtVMJHDaOjC
i10TgnmuYgzmEI+nPTjy6zY78INSPumGDljON+dcxf4d+7GY3qbAdker+P4m3jcF
hDUqB0j7HadH71L/tgzpw5l77kzdHMfJk9/Y1WoOy2A0co7LAKe6i/8S9f1Y7Qmn
PCnzjGVqc+pIoq7ifBHRfkauYK1l+16pmY7+NNHfS/8NJwqMQSFJE8+SJmGfoSFQ
2LpjUnHGCp4PYgr+9VYYmOus0OXVBn6CSiR+7BfAC16OtHwxQRxC1roQYt/s8EAc
v0SiZUlb0IWBO98UXy+zu+42toIHI94mZw3oEvX5Sm9vZbvc+ZtQqFmw0bu72bWE
2Sgz+kOxwQ6BguTamWT3pO8kusFHOS/aeYErDW14+Q8g51hHCv0nfFoLT2T/0c2F
vJcFSxWRAVFYxOcSgLLs/Ho1KzPYNh/gDZ3hjW0Y6dzDqlvUINzGlv0z3HQ385al
ZJaLvt5R5oooB+T4c2yfVrE0ucuYzUli5LGIu9zeZSZcsB1DWkZNGZvxvYe0EG6d
anSsyKttVZC6Fmouufgoq22GqUce3EYn5WG0aLHEr2gmLARxGt9nCmffcr1HqXXA
o+Sl7W1wFNlpCSBjciUzvNAHFtSywa9kVxpc3T1uUL/4BS76uOv4Relgo1IkXjTv
AFbuZGiGVzPAPjaXdrVE2HRb0XoXqrbTKD+TPkeB4DDGN8N5yqbAB9TwpslHVW5K
sA/QkHDm/Xhtv7+4KbjwygHUsff7oB+Cqlm9aMKnrkEQO+ON25oPd9v4lkr9r1ZC
ktifAWnUuBuSijHZEvahnOSylrxLL8vQjDSvJZpFr54enagB0dcLTkCmUnCBEaCd
SSDqIGsb3rMAvj+2L5dYLB1F1+4vEKfnysfWkbdPRf53Tq7RErhEKiye480QohNQ
yDBw74+Fl03bHUWKjdX80e12WVSbYujIdIAONacbb6diH9ADVu9h/PIDEe4szNvT
RAsGirADuXfXJs8EyveUp80VnVuuCOgVnWU0s+yqxRk819dbCAYUOt3lF/dkKPxc
tP//0KFPIayyVI3vo2sZIOYS/d601g+jbFkSh3Q0RvjxlPYp4bfqud8tXmeEgfw2
t/dKi9+XxIKPWj/dJfZGvCk/DYVVapZCNGIF1koImDBlwDFEUHJmlFU/pOAUoZ19
Eh+VnxmPOJKGjAh5amYFgvqN6NUAu0UH31JSkSo/MY7QnVC3hybnsvgMIU1akAg9
nzsJsjRCPWs4iZZchGYTtffWN1azNa/4rKm9z4GLu54OTxKO0op/el7PyCg3bXbG
remO2W1aM/xAHE4NybR16RRVTifsHfVEAjCyPBM5nmmSmaPlnMAauYS8tYngQp+B
yQLyXX6Wf0sd5iGdxXwddJEBhlIt/hnyL1AyEmeSUXOnYeBZM8CuCTH2r2WmxuRE
1LcgiPmeQr8IHkWpRsKrpxFQcUIOFa3anGiPMaCkSEX1WQCB/iPkKiEibufljmQ8
hNmsc0ksUYo/8CYt07AIvHtnh85qTCMmPN8BWOdxPseKzVGHLD76DOoXw2nJzT0t
ZN3raXb2DkyF3QIjqwp6Mhn1tdqZmvBiaaTBGNtJDcw6EbDmoJ2t59BXR/GEDViC
DR6RNKP8QslgMzS2Ud0KhVsiaagYdYGvRgKZ2znlVcVaC1Znacir0sw7FR6CytNG
JmPbpJhxiyzMJ/pVTcSJp9sIeVgYQmRwmi1qiScl4NqJpXFjfNpf1vpw9X2ivffs
+5lXyIFJwhfhHOXOnUypNMf9uttB1MY57EM0xo0jg6F373MFgQ91xDO76J+HtPGy
TAf26qEPc8A1mFRpmLtbIg+nWsO//uCYqFkxGJrVU9JxdP5UsO2duCYJaJsGy3QB
AaEaA/A8QUQZa+oBZaZXEQbT6+7f4a6BcYbjAxE92NwBs8aLa4+P+vRQhadwJboa
NmUKFtTS/7y6Y+iMOwOPeUXvV8KXcRwGFCZe+35r6KxXpgiUgTwKBgvjQ4vUc5ad
VE1GpmXTSyWsNpEO6Rp7FRZl1syQr7WFgBNTYvxW+OplGF+X0JsJnM+CjvWOaN5D
U2RZUD0tltijIFq1G0nLanlLVcf4gYtnURKastjWscBmvDKK+RWaRQOBesai4onl
Fna6wYCER4G2AW7/jA07Pkw+NARSNDpdS23wcr1tj6k0CEKUrvmGsTz4CkpYFFqJ
X515yNWtaifY9tJEw3kwjvIJguvzmSJKEbcX7ixkavoti7+R94AVqOZUJ4i/WCvk
o9VZI4moTzqb/g11QqqeSndS1dOmtmmpQIVUm82qbxn3ETWqEdiS6JIgg5wj7T92
ZzjgkEQsx3dN+cnPBlCKbOXTeXzOnySiinZJnviU77175SVggFE9k4UIKp16aNLL
bE0k9kYFw+tpbvYDfuLjM6eUfDL9e5gawRSdNGiXNk2N3v2AERzWOQqdzVa/x9Hv
Rbz5Nk/zUMua+6+2MkgAThOwd6IirJ1D+zY4cxP0xCE01QJLO/KkiBuDML5HZlBp
AtHMaEbwSoMsSvl0liFFTAaaI7b3Iu520ijQTXOwBhd/64G053Rb2NbBpr2LrSyt
MO65XK/YYDTbPMuGz0yVT581oOo3DTQHOB0A6DXlnl46R8o9zvETTCmgGPJIbAPP
ZpoMFd55bwGNOauzDQrpnsdFbfvu4bUOYkCHqqQL6fszGIPHI1WBcWsOX0pxiuv7
E9ytGsmVcIiRIKEzygdNbU9IbSZ1VkVjTAHWHezmNJOzmMKjsHA5Su+MS/cV+Sew
9YArmrNNUtyvnP4LdLNkFrgo3MR61K7/gICwAOPb+lOwGC500x93X8egnyoBje1p
KaRhSIKDtVQvAjJ6eFUAmlPAyIF1bn+bSsAAHTfDh93qCeFpEHD6o9dCP1yOoWBi
jEWpzCs+LHYdIJ03i2eE0zoAQdPQgKJu7DIogdpiG59BiXjiql7KtQnV7fweMIkg
SIZ9unwfVhUSFcmPoVgRUYlAT04ALlmdATqXMb9YOTH0lYwaQoNtGBVUUQyMBOzB
uFXkJDXoHaOIcWrnbDtldywHRRWEjLIsBAegSHFsdH/w4Jc1NDYiQVGkiOOsn64e
fykXA6x8QdNpoQBG3Qx1hi23oseZ5t8M6RgNYl/EU8N3AA7hRn7CWq6LvlzHFrjM
SyRGAoN1SgUJUbkAXQF9xCF/eoG4G5CJtcQSiuz153GXdFJq3XV4kTAMtDokMDuR
Fyf1iyThzphI0t3FtXUi+vNL3v88rTAWNVQ1nQrt83en0uNaxFgLP7rvIaLry7ss
12qosg2a5T5CZA+X3Qsy1PWjFtCGc225kilxVwYHrRhLIpmJfnMNX5xSCozJJW/v
9zRu9H14l6/LWjqy9R+ud+6r1nd2bfhBs9DdzePlmQHprG13ylPNozyEf4DGspFD
1/BanM6ddILXQvxGjoitsox0bkf7QMKfsHc+GLXZL189JNCQSatgw19LZQFeVARb
hNbsbr/CFwwgc1pPjWLG4erJxcRCNTjJ1e8pmE4gdWb9nc7CW+uJ/aQRMosXEQZ6
ki42oQirjUJoM1X9d86aDjotKL/XkvMXZmPqv2dtNoUl4yEpLJtbqHfFKM/0eWOD
yazsbP1uJdvjvbNVmsBNmdUq2TG1vwPeL10HXrxEGvwM4UjS3OAuvxDzGZ+576xE
Do3LPoxVQKI8L2oB1ELQo0BSfI8piPliGB6MXPlZMjB/Dv/DdDh4jm8cz+dpJ5CH
xFvA/6y9r0AItLRMXrdY3NxUyXob/dU2YdMJzG/QIu0hg9HXP9sjeNfYiDgsC5KG
ShnTa5I5JYzcN2v9z2g0z6hNB3TUsPr1baILL7bYB6f1Z6gDv3yGiWzbMx3NYD10
KbKhpS7eH+2cpAYwzzZKuPjXbJYYW26HCPASd56Gb1mYH/6b0atptCIRsXX7U+gA
8DBSjOGy8FTOmG7WimcqDHt2PnGZ21Ua+PlwvomXtP3xnw3qysIfFK84Eedh0AE+
J99h47YrUQioRHW3VnE5rqWhlxfaM+E+lbDeZQ2AnyiJFfoRluCci76/bxL5fuoW
vR6mUMklOjjV3U6EfBgbl4XFdwJSUcNRgig0jkywR9FLTeuYPG4F+dDwauXe+bi0
1PgGL0Hi3pJcHCwXHL4E5kwiutwtQGJQT8F1YIANVZMNYG1ZMKC3vEmRo3R2Tdqi
YzRDkpkylBUgl+PotpYEpev+tRn60PhmT6YMaXngDBwMSGA2F2G39GAada+U1nWs
T3jp49qGQsphvDW3Tlpl5YcTMxHExPAeb961eZKWctMuXdc0w+FEt8xLjiTyF3sw
TDKe2hAr15l4R3ie6r53l3dV6MkRg8jynb5TOqYAPkAPNHUER/9YneKLpfD/7Pe3
Ea3KywTlkqfscHTI4ogs2hm+nplLfNPRG33wk4BbWUshmTAtcVaP1houbpb6tI8d
IziQFB7ENuI5NYcYKKKrTUsO0kVzJi37vbzjuK53JuTtj86KiFap2J9ZNg1g7+/1
HXEmNphkIdkL7+/Ue+pbPIJykm64kDnjEcVQO8/R/MFPveTwJmdquLPRjgrvdqRN
yaEtW9OH3CCNnGgC6XJ8uPjjIJ9fgbHpF8RoheWA01qEMGReSWNVysJMLH3uZ+xH
iIdcB9d4MrEFnoWll+3dWtot27Cq+8ufCxMP7YFLeiGnbUywQ4OO7YBf8up2Q/or
0DaFPVOT0HGVY5oLcJ27+9nSCKPseHRtcHGKDSl5RWpew9caII6D+muUs5xkDKJU
gwtmqV7QHAqdsKfDzYCP7t1b6u7xJdpUf6x4dy8NMNpsqszBJB8ISpC7qOgAmGrs
FmCU+RzdX7x4GykyFM9HffBZGbp2cTunetKl5gdYjAXNZY1oHEHLV0bTatrSUb3i
9zRmIQUeaihpjM5qxkeeK51s7lojGpuSrsBGrFuBqYrROax64Ndz9iFTbrx6BDaZ
B2q/hSf0sd955ffNWyso0rMaYx584vdI0fKdXMHiFDOm66V2q6WbDaarhQavrg7G
AxS6R1JnrrZGnIfSBjpfcUl33AuUTqfrGID5+lBUX6E7DqzHoOuzgPqB9dyUfYx6
8Iuupp4hVHZ9B+5HA+1XHayTJgjEvKlKvyl2LLlhPLvs70L1s6HYDihh2uBdCD0/
n3a+YX3xUOYODIHsq89qYkBxXtqhy75qI3QXWTI3TEp8F2/9Z0aAkETXnb+UCwi2
9wWHFb/xT64leJkLQhX+5AeHbyhWRDm/RFfZpHtFR4rNd28bDVWB2sMDrUqsYY4V
DN9My3FKgkVAYu13t4QFc4mKGTKTv1FaR7bnfm/ekAdXxohYOXdbd92T8LxCTTOd
++fB6dsk2uLibi3j60GMmhIPE7BgYz/EEE7S4BH9/SykC+GUvGNSkCoE4mYgKy4M
hL575hNyWtoXFDDP2IENq7Hg/MdjrmZExSGULuRv31FnNn4jC/HD3JncHnA5mmfn
Zmwh6GNkQi9nl6Wgp6Xmx/wIb4FRgljDb3zSFxEUhDJPDMmygFLcm/9OETTGcDxo
EHL9bTJ4aGXQcAzklJzZDVfdIsU3eHl06AwMgZk1etwbN1phLIODNPmA9PLCp6x0
ywZybbARJWYrTNSI3LwGlT2os6gM72WauFd7+lULYm4WhMvx6Ce378RPfgMWEvSz
mvenXEIRuKSVNmmBKxNHZc9Q7z8GjzJ74IBnQhIRFjWQJlBGmMilBLH72k5S8RKS
INwsR29UlfCg+TlfSGQHMOi+ys4dMoGm9a93gPa6Z4v+f69wARCODDIDWaRkrMtF
vRaEZoJ9aik0jqVZWxYv46UcMkuRHGAzNnmAZhqQ4bRcR8GhDINy6oacYnitrqxS
BLF20GQv6uvo51HhbDa8UiDTacBvPZVH2Mw9gaifrt2g3reZYfY78HI2u02g9OLt
SN468g2C6FXlH21ikyhvdTzCV2oq628eRUdqOKDuIvrA1ukupu3xapRg3CUWRuG0
mKW27c7Z8TV1Ky3KrWmC9w2ZFEIFAnsjEVIly4TVj7s7pCsXYo8PybH8ZOQ3k4o6
aAQEkGY6DBLL+o7GmXuQ0bYwHuxXfVfiisXMfju+NJCyC2gUAEM3BvHECLsN8x3l
k3eukdzebOB/u60+VFm77619CeQSfVZpmhjmeu5sU9aXaC2wDP9crIbNMdGwUZ3A
U5XJzij+DZuqUkphJo3QYeLPWh8LUGXJcr/bipVyojxcrs10k/NnZOVDR7Vra9Oh
/iL5RYQqOrKBv/DvketpTmeqfk39I3sFegLei+J/zC59GVrZxIqI5b0MiVdx4G64
6yBBOdjhYEKKqGoxLKuJ7+R6HsZKkJEKEUCfd/ukC6KkDBgxU9Jj/5gG47opzyIx
y9eRgT6BZ4Ts4hncaqzisplV2oiMi2IkDhCv0LcKh1qa68D5HZsqTzJLOu+rsbE5
7hA3c7eHal4mvoFTdNhPpGWGBduInzWcqwJsqsnpazWI/4OpYqZRkHLExm2Q6xBd
eK3lcmaTnOnkurLlv8pcR+0FOKqvD1G+j2M7itVQ53+NnH/ggcds7grdjHsRFOWH
1jclo9AWd3vPlkGyrGr1NhMBG6Ji/k2l90puRRXEAKyyDUp8GldqrkqBMsERLcpq
wuDogKaeF7qOWmz0io4g2hWGFyuFDsBoJUt51ZlTbh6zjBrbler5IQQe01v7Z1kp
yiWP+eED5JlwhV/nM7rXmwGaerF2sY/rVTt/fF53FQchR+pQKFNzAFH7sxJPAbAr
8aM97TjJxdMJOuRm88/ikwDmZYrxFMzBMgWn13vleb7K99XZFdN3FitNxCnWNBUW
8MdGkrLt+fOHGOg9YNhM27HSQfSEdBEqreqZ1T9hsl2W+924AUxJ1gVsBfs+/PRj
448RGSHmEzSyTgge63zjlC5X12fWC1vhibiMbFHeKdkqad/7Ry5b6/BmqMLMBn1K
/QPwJuFE/bXV92ndl3M/9P2G7mnpWdO+7lVh/+gYviSjfMZnLnxvkDLnVLAeK+J8
gDdkOMJot5gV0vVtBEtzyK9vT/5UNao8pBn0QXLRANhd8ycDlVT1gHact9yL9zgA
T76ZH4xqe0TNUVMksKhqLO6gJu72sAj9AXvNNQU7/SVisSIbEOsoZ/5dYtkydVPE
satCGRF8+hagF0zmDHATyXm0q+UZlHtkzuJt/Bsj6+eHFmmeS1FyInFvzEFTl6EC
HfV/F5SswJXo4touk7lrc/QqK8kb8BbtRZv4rxSKCntuJb45WOCwIyACNx3eyUdg
FlmDexf6RqcZyvaTz5Zfw7VV1dFVgzmnjnv3aqFXUbiWfe2UImDQAWOjChQCCl5Q
JGzrGXt/2lL1AHDSKnngYhuqpNGAEaKnwfm5wXKfA3jobkSrOufnpaHZLTWap1fM
oHFz9pPUIEvk2TqsOxIPZTxrv4EVzsWckwSWzte+TmEvNB8UtxBUVmwoPDqS26hM
cqY9A8m0vje8pzNthWwAA3nM/428GwO09jrSRaGZiXsT+9kQLirklfyg6Ks5KTVE
iUkByTz5r0K3Ta/SRRICet3RviVmSGVs1sXN6PQeJ7xR2k8IFhWWby1xRn5DqMIC
vOYuuahM9yYo9nj81Bnu50mfiZDElN2YmsbPhd5aiQl2tZiGOSldQL6KudiJRlqf
xNEKYF1MPIgj++ZP1+4gHCjNpOq7VuSsYIf9Edq0wDH9f+0+zfMoxNB+IBE/Nife
qOJlt7U4TTHdePGrtv0GUhOxWZSONKnNlDch5fCy356eh/YlyzWEvLGxi3TGygeK
JQcE8DROTTR9Tbwu8ICA0IEoZ09K0FoI8JpC/Aot6qKB+DVSKmYiwiLBT6jxU7fn
dnJzRVUaNwuJFsyLypd1U4oCW2TeQFhdEpeiD4m9d1JJ2DYcDPcH0/D1oP/6/iqV
a+Qwdjpx5Ne//etUtFJp4ey2cBB7ByzLl7TGzcurje7fbfBQVWSLgOB9k9BNrvno
cthFlGCob2o1La/Lujq0sI4BDgeq9VxK98HSwCsver/RBGlAYF1vRMWWVyFgAzHW
phWHzHmvbEJhMDDe7eChy/qicnjEcYmweVTlPXc7OrfzAwnxukdTEasB3uRDWW83
XiDboxaxz5Tjf6IBE6HltkQiDRuqLa0+u192XTYS3Ceo9FVxwlukvHSXx2wuMx+K
vIrxDGFe1ePHSI8kV1bVDJzuCdD0mRlptKux0m7zx1MAm19JmMQVRhtmsH5P/E45
5OKkBnAM6s3FzmGf51//Rg8ZFJVILRrLbw3kkXVoMGTAiziWtyhw5YvOJ+aE3Far
3F4K9hzuTNqHf6Oll/Ri2H9+jU0pcQyB91RmTXks8zqfgUAwLi20Y8XJtpddmOMW
iddfoC4q8gFoAxA3lovsXV/rHfwYO+Z+civWOQI1Ot/QO9+RV7nnd5cPp0UPhGFZ
xjjmDmLjPIxcS/tFZwv1LWjn6jmftsIdYxVbmJ6RLXfCKJ6p7bqBXNzlp8F4j9hm
O9FiTjbLpWZ32ctRsJYJYQdaXMB7JupvZn7IQQYf/AF6ovGeAFvIrWF/Xgj3LCe4
8xh4QEsWti2EqU1WIGJW7bovYG1kkJzZT8zvJ62SiAEpZRavxiPVTAtGDNeZFmbR
GYnyzjajG40la1pxvCW5gHDWLSWLBW2kBVqL3r54ysr4tkuZv35tonfplnr+EuLT
5SX3v5teHwihPdFfuppmN1JRfXoAIG24TsqPnovh6W1lHbJyI+5s3bdDn9P4iAaC
aOF+MQJlLscKQn9YGhxOv+RKqzjWnLY7ncZucYfHyRJHh7POHjFp19U4f7sSAGHV
StDlffq+14+M9nrOFK9C4LolQ6OVb7xCBfs69d4/KXOV3mRU8zyGJGweOMQfnPW5
5/qGMiUaICl7m/ufB6iwMa/2gRFPY8fnBuI8+gB0Jc/hqEaeiYq8mqiwy5C+ABE4
Fq4d4CDeMuKfzhchOK9aQ5FQizKET/xQwzpB1Dqbz8jM9A41gf2i1T1/qysp8viE
JLka1hswG56MIjwbijxwNepnYYe/Xr2wBOzsec6vkE5EA33MRJ/MetkfGE3XkOzh
ZbmNIrlFYZKd/xibaY72QDOvyjAnOK0GanPYfCER32hRr+h3ASq0bgFf/NXGQBKN
WPSaqpUlvsTCh/YMq0AlmziLY4AkV6exTGO7EQ7N4qNchIyy/m2djbmBxjugMSaD
cSSXr2yPkWHXQBk6oL4gvhuLMFK736ISz+LHsQHLW1NCNVB4IJjow/1wnUlgm6ph
7mQw3zaElBcCyUID5snKuPglJX4rPF4NyVtVx4c4nS3FwYK1AZJbWZErxnUWrHmi
GP3jNB1mXkYHMOwBDyFqojctWvWXrL9j9w+5Ni2peDzEqF3lU5XA3aOHv9YUy9+Y
ceUNU6zbZGYTY8sVpyqiHJpL2Lbsj4SpIvTw9it1mRoae+GYkRHLbm3d9NLYrCGr
AhT8ki7eBKgWVG7o7m1CIevP1KvYcWEs9n0AW3Mu5QgKTQyK9spFE+n1nnM3Fy1X
lEARLSUBK/v6cA0QQgmLtKrv88bQwo5AuGhI6ilSVsR6QQwhBiHxkUWjXzxMZR9e
oSMaVy0ha0RuWynoomi38YHy8Rlx0/Fa+yM5KeB7DYlOHgCQB3AP/PEHbLdVefxc
SdxsMzji3YI+MEjaPpY/GcoDQ3A2bcel7OFEQQyaqG/vXGMQ2aeLuQ0K8kiyWd1m
WL1NCbd42PKAGxeXeXvIxBOexYcHD5xt9h7TVWlLQAYe0FWvSaIhnmxn3dgkcU8X
ipHeShN6+twoqo2D7ccjLS96H1ZpZ++15TEANmZ6oYqjRGEfUz3pS0Diqtq3UTlY
Bc6uQgkUiI77VnNlPA8VpuXwkOG8OwLHN/Cpm+bPY9I6dCRXpe7KJxDO2OrujtM7
KfMmyg06lwXiJmrUlssE4kLXAMfeipGpSNg0uV6Mj4x7uxbD8BWqB0APz3ud+nG3
bJLn/NLLeeVRgJ6bzY5zbEdo8UvzcE7yyLH6fTnOg8EXaZwtqdufL98OiqRgoXpx
6AgPOgEQrCZowH9sLsj4l4T3iWxjp/uBE6GDuhziSD30sVoYk10oWpH05NmrusBE
WoAhHmGbltfJBL1KUI0UOn6dcT4pJzB6AfnMs1B5wIrs80UrJuTrdnjkTlo5R4Wq
c5q/ZqVWvD3SONSwdXNu46ZQi6+1qdl7pYsXKylEAlcKHkdA5VnDo6Otpl243By7
cOQ7DY1yHaVgvBTEr+QHor1ZKErGB0dit7wX7PEfYBG90JmjhIo2HDRHD3674dH7
M4FXs3dYVtCXNBvIX88MIiRrWZf6iv7ygMdrr67zXj3oV5vgqk3xZ1pMsm6YCF7e
IX5yAvDab+dYPvhH1MpgJNadVL4uARlTApgOCxGCo1Yw7yCV8m1xa2T8i9+2qc4s
WhZA9a7qHR3l44xwF6/Fn/uBWlrBLVabMGAFdPrBQjqka67wsiW0AeVXl1Arwtwg
bTiL/5WSefVvRnq7veiwwPIyhR/tznI9vUMZ94hE7GhsmGLRe12mChcQVNV/9eC7
rhKMqIF2TQkqn+NkTUgYUkWqCClJiQJpiM/qkQHr37tqAK7zLOyk4zySHpbye46V
YJvzMZnTcesVch2JjDOd31+IRXQgiuJsPJUnMb/C4+E61jJlai3A1CVILQgE80AR
8knFfnttGDcZny0dCxYA0sL5IhW8i4Uri5GhFztHtsCHNM9yd394NPN16pwtolWK
Q455VpbnSuVRFn2+Ahvc4OTcoLspZDVPsW2CZX0nsPoP53sZwSSLWS6nh1Tn4XRj
mwfneqjoFh0Y5PBSYa9QzVKnN04oSPeQgXtciFjSJkGjVS+5ijFvTIrasxX7JG2n
KDv6X+SMiM81+p9CGhtO4dJvNTyZTsFAxI011Q/9gKI7LTEjOzksJjpv9QRB7Ksr
ZhX+D87OCwYJ2BJZcR/urZytGDoWIYjMEWKryUMSTGJt9j1oToKAPtqfyF+SLdyO
oHAGTznI4QlOnMVOOqki/eMDB/3F4cPIV+gln36W5rBn214NJwVZQBagH+N7SWWX
K7CD0+5ObGAJVLOe4mQ4eQcT0/x/8Qgyup/NEj9RsW/4+kdESBV7DcsHpj4ZbteE
FSbjjE88jLZFQNqv2CpRPcJKxpwvmTdyGJz3CTITp+7OUETeBXHMfkyD/WtUGNP1
pH75alzCOS9hLceYhFIbhMigd04lKAkHCRSu4SDSsIMNMffqjHP+o4r4kC2fgdow
1l/Ik5u3WmOVsEpZtQ1mxsyl06GThb0aFBloxQgf5kOd+PAqHJ830Opj+zOhRIX8
5NsXBwEeG6/kSYLXs19MLQpL6kaBetFdKWZQgPGSzq9dY9eFYJsVWXxRvdwqoGJp
HuxR+iClr/f9rJ0CzNu2EGUaecHIUJJ4XUn/mFwQA3iEUgEKvnabkMj50ZryLw3c
gFwaA0YGHo0ctG/XqBnYRR6RHvd62FcuYDb23y+K7hEQDIGd/7NR4a563pITzdFO
f2JJKRRvswHCEOb6kDvEOso1gW2l5wK/Y2IR6f0h99F1H9TBXUfqT+hCy4Qx5Qtq
1hvtdkAoD+rZZwwnYZ2lLGzNmw0gjOfDbWIbWfvet+O8CIEmsjnFDisoXcW5WZ3g
AV0hFGP3rosDsz/rk+f+hfkToYv39RieQ8DXmc6sOEPXqcRLN+9SdNURnuEz/50S
/co8Gad56Kzr6ybMlXIitUtK9q/tEyZ7NpISWmSbxHTew00cI07A2PiM0w5ZjHSM
oUOe9VoUNwyBuhSY0Jbm1nuRE/GlcT5orVBeJDi7vq5/5o3sk2RkXumItk0uv3EX
8F+XJOOCE7bHVeAYSA+yfOQp9PQS72LfWmBd8ARNLVjBqfdHATTuDBYnNshYEhf/
ECM9jDAIoVy48+8t3q6j1lntOeR7NV2ebinfPm57EJrlz4EW/dh28G3bQLDczHxz
qENeyEZJGg2pOfW9qtZEgVff3gRxTpTOPw4jaNIMjTmqp3KbZ5BQjjLWRNWKGhnb
SXuaOLkqnol9mrW07504ogHDW5wcXFxs2PpUqmWKCB6L2Clwx0Au2BEIRx/ZnMew
vcbsmyI6HhQjQtg99SqCppCTUKSTDW8x0G742ECgWaBU+Hmh7ZdmcWXj0JDUVlv+
Bv+86hCB4dnyYSy+0ZBXJueCg3alEI23/M9c3GHmBzxA/M3O8GXU0v/7k0xGc9Gj
Zf6x4w7P1/EYA3S7U+yo/hMQAHoxFkZs3JXrzqb41+InHyA/NRBHJwrxGE4Th2SG
Z8FNsD7yazr9whbXvFVsJVPq9h9lca/26vDv+c6lZzJmPwwxpZ8uWlWCjEqSVscY
7gUZC72I5ohZOQ7LSWr17583bepGCLvfuH9RD7tjq73lrwdoORRljqmD7NeT7ADr
SSTaKgkOvZuxZCZ2UWWMgfzFHYcc29IUHSWwe+56zHx8YYgKtO2eGJHAwlXNxO8A
r5P6ggSmKacFfvtQCTciWJYry8VZK3IlDgCMqYTAaBHbRPqP0EHNeaFNBXjGRH0t
CPp/vAPByhmp/WgwPpqyuQvhtNYGE3s+Qn8LE/OA3NkFvBjhqG5bh3MMWI0kNh+J
wMtC9gaXMHN4w8FOIos3rP2qdqtuUHlpTrYRSp6PyATQhzB0dgfq2DiDHvmDJ4/w
vPTAQl3w4evqEoxb12A+yFKg2bITRjlSFJ1NB6ASL+yx8lZjMvNAfCVyGE01Fkuo
817NfLIY4/jHOwMNiQZiYCCxdJ3vHSNZkxo+/nOy1Ew=
`pragma protect end_protected
