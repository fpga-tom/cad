// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:53 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JxZqSJf2uXTi56zehsJ+nosgixhik04MamklJsCXoL55PFXojvs32uaVOsxv5bb5
q6p4IOhQN4phJipH47b0ff0TMR93yZby6W9uKHd2i9CFkzMyI8rVieG65tgKkHiY
fadwSEthA1LE/mSR4uBkc9xK9twyIR+ltUugq8wKGO4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2288)
7kIpBdVyOEj4ondGEmLjrXhfT6njljIg1IdEmWOV7FAcMh4imXJEAJ0jmsBex0+9
zVYDCzPjR0GvFkKP0N9oorc2jFNEqFdy1O4LfQelRaUwaRBpMy0NzXsI60izddl2
bDm7V/0FXuG6xWRwqTiXG/N/iVrMp2FtFkTCk4vOR/MVB4nlQX74WU2h4V0rvJ3t
nzUk5g25uXIS911YFYDI2cnAoVL2oqpvlYaL9nH7M7gt7csDDqT9wlyaFUTGklZN
IHuQOiTIss00gZm3Pl+wk7iQZ/MX0m1pMmAuHurF0GTMw2/A7qbKpUOEcYIv/Wr4
sbeXr9IE6EBFcZcv0hp+oTQbj8/ThTJw+hIvdGOF6u6bcoxXglIYet9crSpbwoXR
fOCLZJB7T7sbBBOOS7htcAY+VS4XfglsYn8BhXUHuM4WyW5qqIoGq8NrHiTkTtNQ
nuePjF8uFBwPR5x7jOngbPk3uMAw1xZj3kcC8j/8mcUrko9A1EbBwr0Hxy5gdql5
IuGdQTkmcJfzj316oAhk93jwxWVsnOlcVeru1Cs0nZUiEPsAoMqrwJ8aLLQNgnPP
8+fadXEb1wGwEfwEf1tISbAHUXC2aRRgjQvtM+Cw4lzI534sP2ymixO4t8364Ila
qR51BmKjnF7d4fEOFxw2zutt/my67ZH16ba4/B9EOo87HxEIrdNPT5MHP/yFHtX9
4qXQn1JoPzS2UiK0RU+XPtPBiTSJakxq+nWVd/c2MLVKevWdr+h4oLYweR3PPKxT
sleUQ33PxnP/2u7+tjvq64iLo9GfTkDKsWn/WcJyClcFDT6GSdSHKruiVsLXtLsI
tvG1X2iyS6Qccc7R+8jsRPc4R2cIweRzwXrca1Is6NNRpzo1ezuO5yXPPt62J5ws
WohXEfRhpGVepNTyAnv0qL0CCIYCtNtVWehWPwVzlupvLAwiywWoevl78//dGPan
7MkbKBpkah668bakp2/rDH4plXTKqHrsAe6CyxnCT5xIDZfgOYHaOXTnXNsfBCb4
X3buIQIEKyHISC9kG8TZYKrNctUGRfRaV6t+fgriZC8FhSrt531b56YWJ8qhtuAb
brf+9EWsqrgDlpED9K1AcPcCLOuc80plvh7g7PriYqEHGqJkEBTv1mld1ZweZaRF
DaJEpALS8+x95Cu1HbG4r09LP4kMsw1mvHD477YIHzFHMRskUI910XwuIMKyUfiJ
SRVS4rMLxFfi9sDAE7TwLreqm6VPxH8A3hC18noXF1enDOm0nfMusEdfUY52Nsb7
ksI01NKNlB4FMufEBgAumI234RwkyqsC/7l3VU3z78EH0eZdhwTMeV0iqMMXouvK
WdXrHcZpqeMdtMnvygbWtI9zojeDQtzhu8vc0v5PKM4FzyYtSlfx9Ns8/B3iTBl3
PdnZd1hHJsT4FPkFISX8Qbg5g+F6v3WtrPgIlf4WU/QX2IXQk/+AKAgTix1K+m5a
xvAiu5H/qj9t2TDOsAcyGrnLbJ1uoWj1k2QHznEp/8GGKfrea8nwjEsWfjgJ7aOk
QkYeTskHKgCYJl7YGaaO1TXFceXtozJ6yzc3HLvhjlVlbg/h8HhfB/oaih5QOjFT
3gITjjzPnwiMOwpKk0MtVj0dF+um7CSKuz0MZQUpAm/sTomKmt77nQL25WU6x38U
e8KgdoxDLtgzD3uiijBYDURu7wfC9qNoP2t6MDgkhSmmy/hMR2ADx7S3phSOn7ao
05IZFe6q+hT+lRqz4sMShfR/3WsoyGdjw4/AJtNebRA7JV/cIu+eF919Kttvl/xM
qw1C5d12gWnAMWseANGGfL5qd871qdoMFrAABkChFHRUn22oKFRvrHJZTYsWVTI/
fGnuxye14TSoFB1sy7c3wtqOHitVmrj1nGHCd15KJyZlcHfGmzx01xuAlnbwBWv2
8BqPNtQSv2Bkztw69BzY9e0rEaBs/FATtzjvjH4ChtHs1iNoiRWr0kE8K/jYLZYE
ZMuYZnd/AjQOOD0WHeVcKGTtEl8zj43axy1xrrP/N8wJl8ljXs+mPWMRDPJTXAqp
ZYwQs02O9RGVyZ/Tvzf5k2UyI6KTlIak7Wir+Qb2CEGuzfwr+zadfFdXD0hUVbLn
Oi35zjumXvhK6451b3mQGkRUI+SiUh7COR+QWfw8pPTA8cnlYhiE4S5yjeeCee8Y
WMnlgVQxBGYxiTZfNVHLXM7t0Se2JQO08JjdCzUvDOl5PS+HWdeerGBVM7RQrZ4C
oYNMagiF78PO816smqJfzIvoKhTKBcbNV2bd92G+pNCMxHSUkdG4Lg4WXbGczsqC
6k4B3cn+b0VacuOBKQCHcv2ctGErjHxLD3xR8AasiS3JX4dU1duEN9xp1lrDkIZ1
e5RFZmkYYm9mRRLd90c2trrXz2qzuh2HTJ3iAH53QKcQBHuqQSBFt6iG4ayzh9l8
gdFqGJWKT0qwpt3k49x1ab8qHGp+EOwKUnmhyAfxdiEF3U/EAdJI9WVD98FhrCfF
q0iZSjuAyMFkDnIaXpYWQdjR8hEZvGrbA4rw/g2ZJxRdZpqZPyTsNN/MXhLA5pXK
r+vCl7Q0jXVDZKmghCsiHwpb9oedJAEzEfJ4sDdiSQVx2/oSQtAweQR3NQtfUt2H
rh98ggyAx1Olj/CQVCxd2Ufst8VoW535wp4FYOYqgqB61O4lvu4N+VK/Z+eTNT0n
XIi9gkajsFDm3oyLitHVDztATV96OcJZNvgjm/4MUINEwMXjrPUkbArTrcOqhM5w
NR3taaV9AwiPNYPHrWS4aTsm0tj1D2Vq4SDCZMS9502K15fX4O/KnpG7tnW+HPif
Z4xqboVWBmm/QSZjgIi76JSCOIflPswXxxRMr7pSsCj/QOnyndl8agNqK7Y2u8Lu
4lxoyS6tfePRcuiobDDbPxzZirb0dnWRaGbG4hv6FZJLvbqyS7hFr5jEUADylLuL
fuGCkPvRoBdYM8axlhqMySQ9NqpgSwmUDXYggjl9OyriJ4ENVAAyFYIKCy32vMR1
QAkqvcS0QYnmQEBhgboNWuQ/MvQUjXQfWeg62BcDTWk=
`pragma protect end_protected
