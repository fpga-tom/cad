// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Wm5tUogD09gtdGkTxpxMQMpLyFcoMFxIV8fth8l9jPQJFhVMqcpyojQFdlk90UGM
rNVV65eNgb1YbqZgC0v48FObYNiK86Xycoz3M5N7h0YrD4QwgOUQhN4yuQ582j7C
TRHevM5O1OtuxPXEgv/g/XR8ZRgUrYjYk0dRjj4s60U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8272)
7R9tNTtA4fM7PQ9q/M7FMkkgQ4ojpT8ulUjlqE1RcL/qGsW+IiKFVTu2fLLw5Qz8
1MCZeVtQsPRU12P4EEguoHJTfNpyVhKLCdqH/l/WQafS5SswBiqunhtNiOWzz8g1
2cjp+qRuGXEZ8Ss6FoH79aW0EUNN/wNu5SySBvUJ8wF2C5hmYLtN6Jmi5KA5yJz0
4v7o5K0n0t99Eggk9dY0ata3xR0FQUROCXMYXpE3GBvp53o7DCUADZpFLF7pLdKp
LxzxOELwSBFGOVHjVbIiqbjWrdQVGyHKY3T1IXofUdCimlzt+Z674KCOYYWDP4mx
vOMmSwuuJpIXQEZ+uIt0NQV9Px8SLjEe8IUCKAqS9xGC6w+MVG1gtOMVVPbMzDRS
/YS6gbdyfvIBdsnxtTgAF7CemFLBH9LxE2NXrGT8DuTybyq3DhWUzNtRJUymrzvY
9bJec8cWWEqiumWocxdMcc4C38zX3lwt9SfPJpVUXEzMTG4YyHXUQMFzj5cYZDA7
Jx+mAccsLesslihb9yW+pAUhGEmp4X0bDMptE3vVW8rFA/ihn03WnVndA/Lc41up
Gwpdwo14RO/Z6Eozt3imVXneGme1XSjr6JLmW6vCPTLLND8p4y9bD/Dukm+JTatI
cnEERlQvQ3JF19CdRXeT0y+EfL7z3E2tYeylGnaLgPwJCzIum7linP8WuZPTEmaE
pbr/Baajkbw6GQRJciWSIwXX9X8yvbnalACOLipWyQ4nieLT4lob+gkTf2B7EomC
VfnKHFdV81S3IsfxezBoHhrBEEYGnmUiiWrBLnpF41XeJX0/ACBi4nxkGeZSJLdy
Vkdk9l0BDXH4yoOKXlxpdBB8OV+gg/tDhch+Gtfc/v8/Jdcxsa2YfwdVgus3QvxF
cIgTeZfTpHyGSxYkZCawbLv0z30LCroJybJGIREmw5+oaKpi+SuKzEYVs09G8KlX
R8CRBOwqdSnkOoa8Th3IjCoI0omYzop8TWxnkZ774NMfWXX26Z7DTrPh5C3isOW0
7Zm92pfI9t/j1eKxA6EAQYE+w9p+vQtislNY530uYLxEtFDDVqBRazvlx8J1K4Eu
uWOUQHKrJNDxz5dSAZ4U4cwoV/lbrFTuwfSWuRe/wenCYg+Ua/af0LxOqXhgMPxZ
r6G2AYHROTfK4/FSxvU6Bb8BwBRgJHaLMryVqGSslcPdDglOEO31Op55/LacvT3h
FH5pzbAEGoSEeg/Rge2AfjYRvezvlxA9ZD6r/tDDSqrSeV/MKjFL4+NtAXvEG128
dtMz3qMwQF7Diaq8umtrih7I1F/bdUK7QUOkOBXL36rfRNT/7pMY1++kzjKQ0rZw
qs0xkTqo1ldrq04cyPhfKAY5BLkA1v3JiVuwAzNpb4UfgCk2+X162xrew/XOfAHS
ZeOqdcXMzVeg46UBuW6ydxPA2czKSXXb8iZzkoGB2nTjcw1Fvc6IK6kNcjIGVkvp
jLLGHiZY5T64xDo9SoNxqB18NUgl5HmpQcdcuG9QMBGoxwEo6fdbnXAulDEGAI0Y
1CC8ZElNF1D1NOLlOUXUWThgrQIgO2m/K7BdOY16I73g3ffvpnFoWKngdOkRTTtG
+P0VOLvjILVaLs1YJ9+Szh5TKKeS9xvza7QkghJ/jXWnvUGjM0GheReFFN4KpT9M
gfETvQl/MX921K07oN4XUsm+GrnhWiTHSlIH1of50vZFQjnm78cQS6+moP76Dy7y
gF45RkpkdjcpFRwm0Hc8gxViCBZEYQuLUspSgjpOdWiYJZuxQcTbbgvHC9ObMLzo
kijCCASDsKmh8tWFIVXFk2zs6t2CJ8GUtb0S+4jBUACHGdyf0GRBrbKbURLEM5AJ
go4DY+JMB+Grrbj7fv5Q3LuVBgevx9Nx5893cU6ZZyxfl/N39fvYT9p5m0TQANWr
apyXnCRjkL0D4Iv5fhnAemwLW+f6tfMZFhhlA4td2IGXMPTfmnz6rUsxBw9TmI9w
qNNyC15+bJWs1+FMXyPcRn2sHV1BqlpbKoDMRYQLGcYIuU9SJkbWY6KO6eZHVgsp
DQo9rd5flun8oPW1KxZerxC+mMhzNErA7Qlgc2H3Z2J0SGloDj03SQZCNNzx4Rz+
yriaqfD1xfKH5gsa2vkKfbq+MXU8q7Htg4k/y+K7ngHpLv0wKUGUJaHgQ/0mP0Qc
99RwFJHg9LgJCgv7qYUJOd93i4k/A+v3ZsI12ISqlPwUqfYVQP9B8Nx9XQNk4d0Z
DFAmjcR0w0EDux4isEekykATVw0jm40RJ1rj1uvN37v/5v7UkUjF2S18fMSmIF+U
RJpalojkt/FuFyyxEe2BTL5vvfal2w14Q7NCSTOXswKbirg8oLSgZevttexHhwGr
FjkeolVIXChfvj3oxqmE3oJUwrpl2E9gRhBS7Z+GrMMW/rekVd4UjZDlHQw8P7H0
g7unrIMaEdjo5EN0iJbHiJK3/ALFBTZCGTm/ungEyeIlT2tNgQ2P2Ufekm/O4IUm
iHXGC7kn8VnYWx4fgZ4hDGnKp+901ghhpwHQHwn/kjz8wxE+68ZL4YUxSb7jf+31
L+k8G5e5NgQZdLTp3m9kymMjKrysOH08W4Qu6OEktV3Nt+KNd0yKZnWLe5LLMERG
JJ9GhYcomeqDF+yfCgJfrLlmyQ6BGHCoaylGfxuYohxad8brIH2tCRDMuQ58U+Jy
bi1UEpXeElTiZStsxk3dsz+yHGJx5txthT6qKRsyah8fQrnuG6v1/9YMObMPNddP
Fwmmqiq3YQzl9XJXbv51+qLg3gXRfJ2dYRfE/xrHhCQFCNGMTm7Se/Q//K6PYGl8
DRq0JQXLHXyJAD+YH6bwVBRH6fKUAS5kpvs6FTW+7pE6v59PvpQiKIABOoI+fp4Q
oGhyS551qUwlZ5kVGm3+s2wVuN3qxtlsAhe43/VEqDbmAJjndCfxRFr2JcPMz1mW
/NYSgQH9GenZazZ15/ikuqlBTRCDluUogKUgSCGZ/1EAdvt1Og1ZuPcCHeaSADrr
m6BGPAy0vcDohqTK+dT4Oal7pim5YL9agLiVPl1B9wojmhw4x+5kwjdGhEGKYmLl
oHOnALijomMRMbKWjqZcK+jz1X7NGnmA1y8KUmAya/gJntnZKZlceRsLnUVVB9c7
x6ad+hWCSP+tgy9XRA9STNk84Eaq0/W4WW0lk/NHmNjtTBRk19N8Ebm0/58Zv2kK
it6jJt6gPibEZToDDuRxPMf5OdFmcfM9pNpXPGkOQ7i5DxGf8ij6+GmHKYXE1PQ5
t+lFu8KQVuJ1hs+EsWNrdRpgmYihVfJ2sLLFkroNk+gfyxp346u+gOrCazoIGknC
osB5884GSJ747svKEThKQO3supGp9nnx9uLNYEUX1koiG0Na7vyi9jr2My75tIdW
o3yiCKw+qequhdbyvHnUPJvb6/OTZ6lYB0yfUmC43oR84246iVjnFJKPNE0bAvWP
kd4KEV6kdDC6H6oflEQjuOrVNIQQQ0vlDuJmnEvakBuWuoAUSkTUZIwsdJlTfn24
6PDF2Pc9nDXT7KprfSMrnAvB6sEPBJFLKuT0t9CFb4F7bc7kJON3i4xB00D9p/r0
6xFOVN4YQCEmOmffRjk4zdDRnI5TelJHa33vJC51lPy3IQVJp8vwOo9phfCZT8DS
tM2HoKKdSuY4Fp8J2fvV05+f3OvD0A+qF/P3mVV9ETiuw7wQQ1NavM/VuJ2WsQTS
PIgHXgHbNQ1fVOMLLX840gHiJhPv8qxJQ5ahsteZToUHxnjfhet085TsxYg+ohzs
DVP9wGkhvi/XoVh6UEz/tofgfdKGxsXZlk+UTVR1nxKS510sfTbufpmntM0oCD0K
UwLIbNjj6Idd/K1eE/FZtQaRjhY4uydS2npplsE/5cT5KRVKWfOVim0akNN3pa+g
InyEKXyiy8fG57a008cbElmxLSifF6pVgCOeF7iDCRgmps7uz0SBAX27DDpeOdTR
5Jk9o2UYfz2Tln4pcHfeXrZUhmC8B/+VApgow/D8SHjmcVJJ1VbnZt72hHYKs8WD
w/sDGsdSRZieWFrzURjkRd7qekaRXfxDeqnnrweg5Jrdp0qqXV1qQ5slQB3EF5kN
cjf3D/wFgUjgxWrVCiVielsSU964Xc8IoMgw2eiCvblkRF/bpsrKJiB8IJdzh4S0
ezkJJzegw6+oZgJZG/pnHUXsAdIq+T15YxBZsJyokYw/ZBoqsPK46KSxkzbvn4nU
t6qZ2QnbGP2WIO30U6ZerN9AXGW8gEBuNU/7cVDGNWkMYX0v/bOpSU7L5jXYIHyb
MzSDLiSiyfLwhqrnHLiB6FGiLWrSd+feaHeZk3KZ/dS8TJiMXVEhaAg48UQ4VDVl
WgtNlKXFbPGTkdAm7Hgg8HEpnZwXzTuN7MZPUVn3z9ZnL5bKwIW4x4LkgxYQ1iJe
7gYXGPLi3WteJr2j7PrgXmftr3PN+TiZNtRb7n55dv84ieAJ6auUDxSISiKj4gN5
QfxqpyydfhlyYu2a2EqOiJy6TZSB9ou8fYSzAsQmyY3TLcob9P1BfIGRApuWxh19
E4eP7RUHfCGnWAzckDrMoWsGOxi1NTgGWAqr2yBDFIsCgcud65MBKn/Lby2+DGNt
oud9LNUjJYKMySvxr4mBUudFMa0oKzHi4miw5dOXvPz1u0TsfO+e08DiNM0NDPDJ
9wegGyGi+TFrmHVqBZOl/TH20jxvBuJCoyFowr2QGzr0XXmRlJTwHFdIHBue9XCu
ndt0s138lwE/7UbAwl8sckvB8Qj3Av0BwZ8+4VQSiFUpw1fcUCWNRqYSlMC7aEAF
s/uOqXcQ2dXuYJP2yX87KARSXp69u8bDkIXP++YedDtVuWEcucqRIeFW/R4DI2XQ
GrBV69lxMNeU1qzxETSn/fHs2f1gecmb1E3FX5XImhPe9Ac1TOTjjW5JMgAiXHbA
wsRAcXGOPurM+f+eUhr5hDH0qTrAIc4l2JKcAL4J1Wsf11KaUTWyYgq7LWCNGWZX
GBuFI4oV4yiAtYhfZD3tw/dVWMdGxx4zzDHDeYBbCtdldr0quE9yojhN4pVvElPg
4wh28kqKfRnAYpzh4MjSrAqGppiby4vBc40Lr+OrMYLMSW/RMJxntNt1DHVOLxRw
o6jjfVmKNm8Y/bryGZeSZT6PUwgNZQIt5QKCk/t0bOF5mbv7jIUa9UND+dXeDKQu
hxm4x9Vqmpfqd0yi2Akxc+OV/BmPFlC7jWrI/Di4l1gTdXqBgIqi8qsM/HIBYuVx
/EJTPcklSj+Q/Hq1yAeHkn4UWZb2fMq57H+6HsDRrixWj1bKXzA4lCgL3POVUT9Z
4M4A1fvgcTKuY5SYSWF1UgSDsSdF4IcRVKWAtCdk7swE+AQoJRc8DJM08YB0pbkj
+mKCQ4sOQJJJdHJhCy66zeM4UOGq1fpvRJBM7HJzfS0T4BBAEJy8n1M4tp5gQIcY
N0MB/Pyc57JhkYQfCtdkZ3Jc1yKlhFXeBMzN7FZoLj1JSv+RKhJSJ1mY9YkaIx4H
8VZwowVd3hG0KIz2xkdcNY8mlBGf7EDDAYdicVOhJbdcX0LSxcpIINwwO6KEcB3U
sAt+lny7Q88cAxwMoTt6f2R3Q3XVFQcNZtr0Hrwta2mh0VNVH2Fi8G3QSsafdn9G
DbsXd80eQKD+Qh+wStGaqhrJZuWRCSn2kA1cDcOhHmZJ0eVYrqDD0fSkAhe88/x/
ARuvSNMhHYgv26voZhYQdevSfX//sKCFMUWdLH2tHMoWP19rDzicvXbEkkWQLD2a
16vZQmRD+/P0vh4X5PZHOy3eKIKifjzkE45ERrKGassOc46yuu87SOs5UJBuK8p6
Wt+KnLh8N8RkRc1hVCDex9zJCRerZ1tWY4SeF29l+OXbqmUI+j77MQCw+UOHJgvu
M0/ts7uwT1N9q1qnIn3JyTnjoVRqX2ETHAzqnfwve4XwgMEE6BFHvdMQUNtbjDqA
oRRicq0cxYcf7t55okjmVfOCkCWrqnqiNaTheCKjAF21XhKrX2zwV5o92KXFSbx2
32KvjI0W2G7MgIdDdLc0dG3R+oYHZRIRe27GZrC8akeiTMHL2wGVddvXfHRs/JlR
HXtA/1/aVyB0sOIDFtHQT1RsTQeom5wioMw7aVpf+HI1PT1mLDKuuPufpTROaV3s
Q/oydt2fuXPIBwOdKgYv0bHrFCel20CtCI3yi4L9xHinnuzN8guTw+c/PToTM/P5
uqBZ39tVmjZ5QCWkNUmMqJAzH/YIY0ImAleBhjM3Q9p7NDX/S9yh7FYLtxuVhc23
oeJ7nNXQkVCYt8m8kMl3Q0SC/BcOc4sa1LETJdmXQ5Q4lScS4fd1p52CGTiA/V7H
oLPtOCTTSnXO3HspaGWZKXQOCg9IORDQfsF/g4TSFiKBRPB3wAe1sLZYjcylzGv3
PgI5nq1XXHOfm8i5lfXdu1sDriBEPWUFp8IQEInqmQkZ50idkcik7i4No35YX6Qd
2dIvz1BqaPgYu8TaEnX6zCk3Y9KH7iDOpAj8lKo4o6Cexx1Ca74PeWmWggBKtTCR
uB509J1X8wd3vB5cCVQR8k4MQq5u2FxyUMCQwwWU75fuzptF6DxZrsn0TtsG/MwK
DNz9BgN8bS3JKXGW1pRSjyiVZwENt+x0hnIZT5dWaEZEMcnyaE2gc650PQbVQWow
Qlm1Yi5sRYxNU+bvk6LTbLUghiRz/b2RJCdcti0qA9JxZ4H7lCK+pwyxofg8FYhT
Iq7rRa5J713kJG9C8dEBn+OSPV8VvQyaKYjs1QE54sEdtWYjOVx9TbydZXDPf+ov
H9JiKzOJXNw/iGwLkp1ywIWCENWTmeCUGIApwkFw5DO/LYP1JAxKEL9gmjOLAksA
xfjsJZRyzG2J29XIKU4oNwYka4aGbwT4/y5xlWaWXwV6P0pwDX4IB3wJUBC1QXJ0
Jc9EB1Cgc5VEr3I2Ik7JEOyTQrjPTH6uB90cRyD0Eb4CBBkSdNIwZjiU7Bkk8jPQ
pc9exx5zzMyokAYxGCNWCtY8QRaYCB+uoDeoWcY4LKUEkK0zJ9SAbdDQbACKgwce
GC8o/t7QkDJW/qzw9U9h3Qst+ZU8Y7TX2E1ezlkZpktRwhUDNuWzTD/yhD9EMW1M
qtFnuBg3wkU5iC+/sgoZVtCu2exExITyKCaq0d2TsFVjFLQJ2ILC0KBZ5p1P+ebv
++1oul/gcmwB+53Br4AxgElUWJjOqVFguOzhiS1bj+OGn58s4zVNeJdTKpiIuXFz
0ZdPapvW5DIB1Fi0EIu8FApd2En9qybkSWonWkTJgBz38QcoCUBlJg6Rw07rH1cN
byb65maygC/W9grZ6idW0OQskzpcVucaEdrtkl31D5nefTULTdBQCoICxEsVF60Y
x+DFPgPYuV81ALoFqoasxd/+0GTqzqd6G8o67VGmFtvzyxK5EqKWgjl4cMjDPeZn
nFSWqtfjotSmI/EVZz0BrTZAnQLbIqGCPGsQeZ2pIJ8AQnRNsjnVyy8PPzxyDSxw
Ja36Z2u3nNPl1m8cR7NGgFIkJbZq8zDBPipLDgTftyNR/j8JdeAwe2APvN96IAfF
6U6QtWgR03f4kEdZuRSiURX1ByPTBnfUrM5g65Uz7YFu2d2O0HTn4rQPgJ1HnLDd
Mof33GKM1Wk0mcVALP+wzFoUP2gxI2RWt/mXFlRClA+vDiPLyL58YZfHu187QWm9
mRQ1CnHBrawOUBrRXFH38dT+pSFFTRtjNJtePxQ85ev/2LrRis7AlHcp/fWlVQM4
P9QG30N6i3Rp66rjk1Ovn2rAUAQbbjAECku0NDJHT/k0Kvm1bDDv0WLzOjkPWybl
4SndizU/BTIawUbjCk5kmBL2sVv0fRS/ry2gtuJf9pZ9pU1BVlmp1mFor/DnzK+i
OZ3IxI/cMXVY2hIo1hiNp17MKnoAyxHaejvcdiNp4xWAFUaJyf1CBrDm9zuPQfre
zBRJvYkp5SEX+K56+MQZAz8QQPY1W7ljGSGxpiUPwDcTIa9bG597SCY5l3to4V5/
n4LFN0XKxiAx8qWyAF532joMqzb9LRrK1dlW+AWRv9KW8JoSxgsCVAuietwjx9EG
Nnch67uWCmwC2Ctl39wu+df0IvybnfaNHBZXbaAmxZUO+Ptdnhh9YokS8rHNYXW+
1gvqSpZqVWd5K4DijKMp5kjJUWVmSM7qH++XS0YPtIJ5OoH8GTg19jnp2piXJDI0
NUAQydPqJ/zYfXh74A2gOfNGIl+vmuzO8gLpCivAKVwWx+81OvK4D8dchlyyyVgz
A6gEpxZd8fgC4o4S1oqNeh63moJzuyDn81TY6Nu3Vyue2dcGW8CUx75/N/jOhrqk
13c8rbaihhQ5oszB0eTIfLF+NDL6hPXP4jGhK6qOzGT0oMg8sLvG4V+R6CWSvk31
3PkOqyJRG+3FZqceeydesGzc2eqQHagSonv3wM801dxuYn1IzE7pQi4KzYMT0Bc8
BsPsjkp32EcJhlKiKVSorcJGBlLUsV5C+SCKka2PaYSX0U1EWHU15wNt2KbEbvQS
mX1r3oAybvTj1ILs7O9QyO9RURYlCfKb0PWFTENTPdB2sfb+G2AFR574GMzH7Ml4
Ua+dOQ2sKGu9UBelPy3XEbWuSZJQRKvf+FVW+c8WNIKC8rQHiWjxx/cxxeEW5/FQ
qE3eDPuc7X63WlOVUd+CZzpbTJ9nf5EVBPJ/37qvz+MUIxnzE07p0dhtIJMb0bwT
3bp0f30r+NB5YTzJ2rRSwri12oAUjwgU6vtpv+RoWcLVNoHqlVqi73uUMSBda1ws
XcPOz5XwSBBOWnatAUl0OFy2lTVgIKBhgMssL8lL0ddq9KFwdCI0v+DVRTW4HstX
Ej0yP9xIeq1beVSOwALICLNmgP0Fdjk+lNB6Und3tGBr2ZXVwzEG6ESCmWhGkkp+
Hu98+uz7UwBIn5WA419AqYARmXA4AnUaokVLKHG2igIWZ3LEwRM23yJUi5zOnCb9
BDm8+c6oT6VO60GyR7j4dDndXnlqrBc9HLMWmGNmFS/F4XT7iQeKrv0+rwmcmXHE
RKDS9QeZ05gR9brnOQL1p7CdXwYauItu3tQm25PFKHupYslM/eCQpprTVDMHLXeg
xVAIhf86sp8f5Zykrr5eTJJzU4FFqJxAhDLfp/Dc/h1Arfpry1eiWsMwKO9wonoz
JtXjZwUVWsSLIerrgjFZe/kPeQBvUxAW3dlNcGs7Vg6bxTZXz+8/bnMj+Qmya5jG
7ZcWxthyrDh9uLr8f93cwmPMHVtCXQbRVqkxqfRym+FnpyjIXkHY5s8UGMGd4lro
0D5ubsaPOikXRJ4N+UAcUxUjpE8l1W3LqNeBPtTzz9xDJRFJooECP1JjkXwnpWfF
ImwShcXf9IT16MagwPW+0FRJvWHffKWe/MdUqivPg76k7xdC4Y9xCg4jhWgREbR0
wLGSM4vihP376EZycnDZ/Hk84TCbWZx7nkXrvs3ZYSJplfAOehAfH0V1fJE9v311
NP33o0CtJr/0YF6zejdOInVN4r7nd0JD/dkDF65JtITeEo1joN0C0jxrqmHW/Uy5
dW/u93N3rTYOw5lgTwTooLLXbYlNK2jXS4zJV7zkc6iqUjMyFukpoiQzAnl/iD4Z
XQTuUsU9h2n5dkpY29H8Y4cBAyeuWnj90wAOET/LpNnUzqN4CweGl8rFTfueogar
bgVke2RIvtgn6H9LS92sVeSEFDAAXNxipkry+A7ElN00k4TXwP4LgStgAMhGkgb5
MxFVva4EVGnME/B067Q+omeuQgBlUftgEP6MP/awUAmU9J9IFYNAl5dIYa5yDOK4
CV9jE1lg2NJHhA/wx5Dsd/Q+JHFGvrfrtC8nxMpI+iQjyUljZcW3FsTIk8ZVmfeX
YDPrRumylrphfpBe6/XmqVUYDVIk/+GszatCzEtqUxmf9jec4/2+m0846nZe9Kpn
S9N0susNIqNFB+y6Ob9vzOF6Rp0EnU8DePqzAualXa+ugRnI4ohjkd2PTinuQ24C
B5f9ZMw1XnY6//SAW321UJ+XQ8QNzu0J7KTlVqHaX1Tj4lUbR5o7zQesfIe42tYw
uen1xyJ96gO8TagfWtmW4Hty85tyjtlhEefuIqI3ZFw252TH32Z4c7sY4y+y8xlO
hgK2LIrXnU3HiIyUFRODHKRBe4WB1KTgNhuFKUA3OuqTYje3CMf2AZ4t7tYD1AzI
+pEMR/gR8ZvR1guXeAwmjv/8OK1CeMjFb0SAC0N3ioHmKJu4Hj7OhoBw1Z4cKDcj
8yAe76gcgBeROAmWMNQB0UvZ7EtNeueYOrVEEGrvIq6DpVIP81iU2JRhBY7W7zVz
xmBzZ8uQM/vD/PlTqHGm9dGU0XKcb8914jkTAAhWmWVlw+RmdY12aIsXY8xTQqtO
ONxyWneE/+DXp7foy46q++joV2uScd5FbPHnhVfz/nGzs+bqd+gMaYDNez4sd4U0
kL3XSG2jYfdcNfN4fyrTSD1Jct79ORrHbRpdwWvq79KvYqU5f68CzwMOEgrtJWA6
hoBxRkETiisvloWRLTIMqeP6bWv3zUDHIPvavoKa8GQDQz49TyCe2NbXLj2sByy6
Bo4MRfpW1PrqhhgpMp8bqvb6KyFdMu29PQ4Td+SBB6ZWJ+c6a3PvvIS//GLxrbZh
XgdUC46jMjFfhKpqVBhTRzDPdZREyJkLF0gd634SYR2a9OR5iLZ26nEL2chqazKp
Rl5gG11GsPUpdOxJEPhxExja9Fs6uvHueIx6qMW28sqhN1My1sN0KQ9gJOFxQCTK
fvfKUnME15VikdY6Ie3BDcPjoEBEWKMQIcDytYApKuWbB8n3nc2FsHW4EkMnphMx
bLdTL0IoLaJWGAB9MhQI+ZbCtnxB/dmaYabKWo4X4+Dz98tfp3ax3i7iWokpElPv
xfEi1Te4NY65bkx0vaMVwMsSlMcWmMIEELgY6zd8u6NlP20U2hN0ZNvhba77k9nn
C4tkpkUQ7Z1Pjv7D1/0SkcqptQQ6nk8AWdVaT5QscXDHmkJO56XhVuj4WUJCc6db
pyuHp39uzR4/EdyOMNBxkg==
`pragma protect end_protected
