// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:31 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FihWlmUPRFxOcLr35nH2iRUiHZYh4p2HFnzT74prKAWirmN0OsLSXs3DlsPo9GNr
UNmVqhqXSPVDXWPzsMm0CcvUJlYjNrG6BgIOwfRf6CiGK5PeF/+mwg8y+ToWyfFx
NiZ2JOHxl6EUz7DHjiBOyPwydikgVPDglJdxM0BIltI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22624)
yQW2XoWsZ+79fUcxuMuqi14ic7wdAeFVt/QPMURRaZCRPl808moI07w5KQwG7dJH
kEtzjcZhJfUTEayQPgPaIkpBxgS72r30nmf1urGkwoDZNxUufgBDx/IQyPbJu9lt
6lzfc4jGKf9fhZVS1kTgbDyIU2z9UxEVMmlXafYnPtZtbyrJEOb2m814C7gWZsvP
hAOQY8FzvogO0JZ5Hsb6RniprtpP1YQhiXfRAeZaJ2aSsmNwnlAed0h/mYEOItot
KWGpCd5xwIr3xaSmALbM6hoINtyFemcf1K00CkcFu93ihHZzEwyiOBpTZT5k/hS1
4ukBD0qqYmOkGHc0eA5vNL8lfBdhfKHFffNRyLPhYs+hT7lW6H3xe2PTmkIQTkEq
poJnXHXAncbeSYg99YFt32AB1qVlGaebkwzBE33+8+fxlWPYiQwdapY5PALOa9Nh
kzTaYwO4EHWQ+gh/k+QWeKI9eFPZ/sBUCnWIZnwNhQ+BzL+jriwDFAvhfIr1ipS8
qvpqGJIlbuk4TH3lS9kFfqfAZd4DkmEUeHTKcM4MZnqEMEf24QaFcblvd909DiUn
G1jxYSgfD3Cs+Ubr/dtkUqZpZD9XkEM+E8mAK37sk9FTToJ+RavkZIucAiZxVw+d
RLL1fLnM4taFzn9AETiB68sBYRqS0PxK15Y1X9jfydSN70H793UnCxJ+f0cA9jWK
f/Z83Cg91QFjKzluKohY65ac7MxTH+J5Fx7qZZpYk91XZKV1rEplVk6EBm4DH5xS
Hl4P0/za5DWwWW4uZG7ESOeOfs804gdCuMngffN9xy2e5AeHinwvyasqprfeZgfJ
+TO2JXRJovlLLnGI69DAI85jdXFq1Mdz+CqOQ1BrHjTWpc0oI1bASYmJMoQE47X+
/9gnNB3yWz5hdBpJkMxAftPxutIOrSoUEQD7mDgVOkAHLFL8xk6c21O1max67ngZ
i/obP+zNHwRKrrNy11iu5Ai1OronwvbBL7vRwA7kkEA0dJCh4I+s2G21PpgU3CFx
d5QlC5mqJ/AFvCnWwOKUZGzX7ZrgJixBgQ8GyJRrn723MTQfav70nuSNx8NiHbFD
AP3m5MChU228AWWUHu4KCLLXXNEEmsF1FFVAFC9tkfODbd5ZON7eKX14pzETdRxU
fsN6K37J56qTBdGlWS64nBEqfq9Zcsxcqxwer+Qvt9hfBjWbBWnNicy1Hm5ZFbx3
W2AHeaepazVBzp3PRBq0UDZ++PfdebrFCQHhB/wpP+eS8BGiVnIbmrkCaIxs3V8w
YgD/cg+1CnlbbVmpVOu3SQvPwJztbWCaIHJUbgVPTuSrAkUdGXrO2aY9AKMds7cw
zk5rN6U0vMs1d6v6b83sh8V/8Qb/mNNqq4n1Nf1djh6BOeqzmrWM5Q+eRIFmiWZi
SuCgLCzlmkxGhPUOzdeW521mo6k1XF0E6e8Ncy4/cAHD32FMZfTT7s4V4O+TpMa3
LcnBDNaXOzFvybmmOFN/GKqrV6JLX2l7cy5O9JeGTvu9yoiJSUCbRDmMF52lGRuO
h16Aa3GmT4HSPHsELUp4d6dHDcEJrS0HEnyVzDcYLPYEahh2xhjQNSyql3SyUIDc
y9OIVwNfMxi3QBdqd2SBrmi/XxoEJ6rTmbnjB3HCICOa0pUu9G1zH1jlbKXhC7Sb
Ywi4hG5XqaeIvoX372iN8FlkczEhPHTa2fsLOD9/NZPU6XrDJ5wNE3HtdY148fHk
3eenjT5XqY+8edyOi89ORnkOjlQtc8+JOV/yHzy+ZdlT7HAbMCyUAqM9BR4YxjTd
e1JVlA77yt+QHUJNkfNyr8QOpjY1BfFCRI+p2/dT9XBbwmCKqim8nklDc+HID4qb
1jIuBC3b64MbaKpyO7nilQB73qBhed2AErehhEwMNPiy7EyrOx7ihuuW8Xzl8dlM
J7irLTpf/X36UZJ7aPb7Qiah+NRHGRXVF7GRYiFXCC18uG4FpY1XVEPar2E/quKU
BrTEykL1NhVBZLIwXC32wL/9Ph+vBeOzD5kLikXcQtjJpeqlDS1p+SM4TqMknPo3
R87b9owV+lQ+cXny0Gjlel69v1/A11iragLRyzjAYG/nIyUaWKbmcD2FFqSOnxna
1pfw8HPTqD4UC+QDzXhOwc7AeSIum2amm3e0INdWmP56Dyzvsq9uxgy1Judjod2h
To7zcmh2p9PzCAQq8mqKUDSzTtgg2Zkc4ipbIUHr1GohPIB3mvb9mI0Q96RVyxmO
XN2qKDa7V+2NuhLI7sTqP2hnu4KIwxPLRez9zzuX4AeiEm5tmYGTCfV3xeuhqGnj
pMAG/bXSpT2TaIxEfhhoyRDfXOcqNORst8BkofH6eUC/7bOB0ahSwKd+H5EN3WrN
MiF6W3uZjm3Jc5OA5gq2E/3kVsiy13smzE24I5REto9H0rjowdCm6ArGj0xxDRYo
Obf0JNDndORRQ4O42U1CSt+Y68ffC9Nu4yQa5E1OiyWk0ypMQDvN/svAsdr5Ftog
0OKYMVnCev8qMXYB+fGicnWHJvuS1A1K1ciPSOAjnSlElFrWNQTkB/i/MfHIojlO
93rN72wyzh4NKQ1cM0sHiKCMBXPDTNoQ4jKBBZfDeljqPrz0Q6AqSq+6Zvntzhx4
ccUdhAf6WDDsGrvOsR0faya4yxkNbpYmhj0iB9t7ZuZBbckpA+Ryq/nPQLjg9Gvs
pt/Y/EG9qyHEA05mVGcdj2VyfV7NJhGqFtp9HBDyHFDFP6R8nLLel1JlmbEPdG0A
S90MK6Bnb31DbceXVd1TTvVFncFMOxbt/HkYSWYQvUvh7Sld9ZgygvytID51q/Id
49qx2UJTWSFA1jdsKXR6GUckrf6moX7KaFgbEK3D1HllYA7nd5JcEsSpHAnW1Z/5
g4YxmimWTBbug+NzuPDJk7uR9OUYM63N0AoCFxYOIYMnAgZe/rKmrcX14MF5aObX
afZqTHMbb3h9rRuzp4oHh+KawTALhzKAx40KkKUYjxrpvvv8B91Raa/ARBHpYGEa
+URbuailwaTyJMwgBz8Ogrz2B2P6nC+SQMmZIAbwlmCjFSos8dXVtZRBoITJvDuV
APk3V7KP/ZZ6tbPtFjwxt5QPqSZzVxisONr0JI4ibL5hRA0nH/bTY2bFcIE67SDB
dilxA5/qfacQQ8xoSVvUnEoIwhK/GPnn4k7WGAlc2OHJS2o64evnnRT/TNbfq1UY
lJ1rd+XPCN3oWkdABsPDORAA6+tOMXTrYfQqqMuukfiRcU+EjXGPiuyEuXmoEE60
FOdjOCzVuJ8tuHQt/PFtUgH8kPwAAhh22XWAjn09M8DatLSbzpDIgMeJYRa9LLEq
r+6M8Hv9apZ26Zo0mVSuxRjgO6KzyTolB95FPGC6h/Xi/RPUaqMwfeh9V+C/d7Qy
sr35whttsO/vfpjh2vy6oSLoU3HAt9iccV3duam4CyPLsHcFjXcaHFDdBdBrGeEg
7E3zXKO8SJ65GcdvqqGqApcDo2fZ2RSoXJ6EUucWXJS1uqYGSnj1QxxxM2oVfWrt
hKO/dRgb7P5HfVZcipXAcc2LFvJUTk+EB1J22X8IF0OunA49sqmFODamBzQOKvni
X88gCsU2xNqeG7c/iDZgQ8RjGerDQzXuRLVxWN72SH2VsVDHld04CeWQ4arRepQX
mTnK5rMkOMKG9W3wyiz5LvNNhO5z4e+ZgSLLb7OJKHL2hL6X8DlMgWOJ2pwGLuIU
v6+BNNHG87oWtWfNlIATiP+Y3O5CMpIzmxj3ykkiLQqlZUQYm9UeB+wjNq4dSNnP
f0ppxTaGZeSYGSBPyFB/98FhxgCmWbQCvEDIVei0EI73+atdt7je1U9s8XVujOPS
yjT4oTJBiPRYvdeuaLEU1njHcWWI4LK2ud7zVEa4FA5iBTgnI5YkIpkRZiolt0VR
Zx1u61+vzYpOMNRO0SdxLpRN7YjWOoH6YZaxRFx895V3VHObilfMORTGPpVJrhIm
OFBTghhDBzbBjyL44D3DgPr9Jo+uPPLl8DIx7vw441FepUsRdazIFlaOS0fD17rk
hNz7SgKKbmliP5FROis46Mc+eT8/cnoHvkIxy1mYSC9BTdraa3PbCBjtkULGo8NW
+u2xCCiws/WEgywCMT/Iza7/D6Saui277tAcCbAuAKT6QmBoCzJAH8e0bCly9/Ty
AInfhDsLCv8sNnDhtKOEP4fG1lv+tt2zH1dFa5fRXtEHj3SKbXxiZMR4JUbmImq7
6CKC5Ze4f7gyOGnUf65fL/5plTV+KesxCyWGFc+UH3tGvKpCZU0YdhEjFMRArvqF
j2ZZ+YXUuyn3FE+Bqh7FS9sPRwqVtqHw1TMLPUO14boolTkzCrUuNxGfnreM5djd
XkZ0Lf8QPo6nptmsdZnD0LFpptO21EejfMau4toxy6XKeYNO28JfWc1KVb3G9GMK
OXhc2tyGtPGfX/koggmwLGpbf4KwoN9RjnMOPtcIbLkjcovMZcofixfn90ggf11r
MuCt5aczGcgv5A0daivLitz4tty0K85F+qCymOBxJJ2wiYHRw/fTUhfgIXZD9GJ7
+CLo5GdDpens9Q+anJkGsOjfniZRILv+Tc/MXSIJv4F9bud6/jr2f6pCU+n9CC7J
iFiBRjzy210p+1DsJBp0+7i2LbtK+Abg7zPnr8/vtoQXv0Df/2z74y5QO3DEoiW5
he5xM8K82XOE8Y8rW92SYCdawOnXeKC7RUw1lltRVZss6RBiWAJkjN7YjlJa4N55
x54/ZeuzdFJFKVLf+qvGd74LNXfIXHz9w7QdcedSpQjZBEUsgjCHTHK7PmWpU4C2
D759fAxuJCw8dLy595bZ5kiIqy7r6m8NfnGTnEaCkajUoFvhyPEdA7dw+g27usrm
M1J76OHQKTHnt2HzLZ77RkHNu/aC5KWl2zVHB61s5oCba48RDPZXl6uYGr6fBFal
cN5fS02wKqbF75Gzwv4z+0LCR2wOV8cK26xYix8t0F18LeQ+4EYE6v+peAdxteRn
3g1wJeNdN4+h413iq05ZA1Ylt6YLeEc7X946TGxNjR3xa+7HXet8kTUsSSxzrrzD
pWx2UKaXG7u6roPzkI9EQ7kpxZOn4okRHz6LJPaa2nWz97xKDWHW5xwn9ccL1oT3
3re8L5wblZjQ96sfdY8umAxY2d2d68m9q1twNxPVaN4r1IKK0gxHLfDJDQqM6W48
nmRrDZ6uC86/Jenf/ZFY8UgqVPQBvYn8Fw2YEHIEI6Lrvz8MC1QAiEwmEKFUJk86
wai8ffdYZs/w5CZitNgVMR55CjDPfQpszzC3ybE/he85bVJPrsoGEMPU083HjbXW
YTCchNMsPD7FMywGOW+OpApC7fbz3BOXaXEj2d+xFW1NshwDQKhH+M3qUkdIAJWm
OWFjSgJN0DX59KbV00NvzRIIn6033/hxlaK5bd05VSKR5ZbJdKTFboz7hUHTQ/ot
AGZbn8HB1y4rxfoWWEBo6igNx4q9g/GQI0PVKTjdLKAc4KMS35z7wKfbwue2j7WJ
SFIwtstYkBKxNm6YJBnokui0iJzPCLdEQHIibxjNrZoDupbPyKHSVd59yidA+dSr
yWSG1US1ZMASmDV43/8AwB6sn/W03adN3F1b+o6wYDqbdv4Q62WEg0CrOyyeIyMz
/wHhc21SUwDrUEetSUnb0DEXBvjrS92jo3rs/hsP6welu3xhU6lOg6lqMXH7xuYh
qMNHU9lUFLYZUtBJ4VC0P2itHV+j2Mj0x5f9hfGJO20386zwolrtGEOMvUFZyptT
Sji94sHQf/0JHN9d9SqRpnpJOXjCwE+zDQc/lKfdoOvrWlij2eDbi0iVzoTdLG2g
Y7qoNd7kO7wqibvd8LgfJCE10DJxyjQn0bOyYaHMm6drDDMJZoWqMRmEJ/Mtr7DE
KLnTdJPMaUbrUPWWDly6M6hFEvge729ZheOsoy5fNIs//mnn6T6uBtp2nwoTMwTG
dMs2FPY8ejAZXkZp42YNc3HmJvhoS7vl44a/7bCuTlE4Y468tc9aRPGGJ1CQYq3k
tF748JwO+Q3THz+yrz/A8wOrD3xCoTZspuP5QqFl392YPuRIfMLJxmcuyXFpMoAV
ACbjvmCT4AlghcZAivPhVFIaexAVvlxA4q0DQppXQ4Q/MgwZLk1y5GJBZEzs00P8
Ar7hxa6OFdo8kV3/3XeWSzJUop37mZiDdQge585ph95WhMEZ8FaKZz5h+2zBGBOB
JhBj7U6RaLThHSqokpH87ul8j47d0nGOZ6gOuRUtvSU6WFWLG526MmtJvz6Cml+l
mLvCy2A8qfrllRK+UOUr3BioO2ZxK4Uy8608c7Djyqmm80A5uqe5f9tVldIMzFSC
uOjtO6W4UdBSgbBzIlf1j26iomdS5hgqwsOjOWohR5AbpxWn+N5X+muS03qDY0fs
fouyYF37iXuDE3xgPPwWGjsFdxrLDRs9kzV5KITgDXPw9PPxP9V3+hWcvk2u5ZJS
g0Rl5EQQyOUjDJfCJDAwkLXsRphFUZPXIjHLXgtcUq+HBkL2sZcEYMP4MZwScZ9y
wwWH8dFftG6OGvk2xQUTKpfZyFBlZJadvUxWc6cRfVyGXpre12fMIZQbitbkmf7O
Mso48+D5p3+tweb29Uttv5ycQrsM8oe0j6FI/z5q00L/Bnp8mmIfqrVB57/sK5JD
z0ucZHRMdHxCbWS+o7C/KXMQ+f1/7ektu62/DM8D7FJWmoDl62qboSapWerhRk4y
iVSNpjL3OG3LtVHbWb7/XDBl5OWWOEN5arnQJXRFRGWYulIaHHdLnlT7AWBgxmHs
y7miSG100jXqERaRjlPLPKz3uFTmA7OMD35DH1SWyvyYuRKxWvKIOmC02UXr4jkY
3ertRU3SfpE65a2FU+kBkGNOKK3BivU2zs60RWRrchcZNDSIG0+3M8WiYwrV1W+9
I/LOhbJXXtWas1Am8iSLTIeNZHItgKxCAkP27Knl7E6eUp1TYT8MlmulBWoodbFj
jlLwKixPFJI7fVXqzo/7BxJrRV49vsWl9cevrfFYVa+QOaWTtUqHFEaWXs2QFBf9
VmyHDSkkbWfJQj+fWK6jNxQI5YuxqPhUQsolVyw41GLWVUzFFwE2v5jrH3c7Dtg6
RlufwWMeRV53OSZzW+PVsngf6Ck12E0z9xd7G7UHRvX9txOXIeW4JArUZaaOI/6c
2sFs2Ek80zQ4B46PhHXnSzb9Pq0Qvb2SMgGphLj/aHslCjb2r7awyzPUjWUTVUvw
hi7fTp92viM5P0s3E0gKGnSV6g76absa0rZTFZysKet1UfiNZgkjv39W5QtAGbZ8
MR9syJFF/n3D0I/1Ca9AtKR8WDYVnR3Itl9sNNMqUAjJi5wY2/jPtg/A10flKWGm
P1zTMBzi5ypy5YhHn5B5AoOKCCOB4gwSphIsZJxbvxm2pmPci84F4abTFz7bw1Q4
3d+6Bosb0LXRkMip0D24kAS5bnxawPpgEQEmQYebrS0KSBOr3R8pl1+MFXG4KMed
+qU+vOU4fO9YcLiCyt+Tpfol2ZqA5IfQ9Sm6/8MPXHauC86fliC9nyjOhYi+/EeD
e70Ccuk3/eXnfVpHqs/l+MefJDyWhjV7HNH/gyt0Nz/sb76kM6TXIvGNcKiSGr3f
Ye19DcPuTft9fBQ5iAUnG5oyTifMYwdg4l4mmzcQiWo6Xa23f5jN9pUxvDvCqIF0
DHD4qw5pms7hIG/GvjIQms1po4chdcO12Em2BuiiEHnNjPqycHhMtjMVt5tA+JNG
3JcMHGdgcqiqY/gpUIVT1xbIMluBIm3s5H2z8060kd/qZBKHGAYpM9a25UmoRz0y
jLhs6l9jTR+T4mjPxFTLi/H4bDKBjoMOztuo8cT5kb+Tf6z/2trWyXxhOCvTi8YW
T5s9D/kMFWeongPOtKI6ATjfu1QVOQpTNPsHrp8OqHzM2abFXLo6/aYJ5X5963WE
Su/Cug3nOhsSyo55H2N4d7gU1axGBJuuOQ/AP+3olNNjEADkkLHJta+UetvDd6s6
HqwOL3W/BvcxSKQiivMkdUgDC2PYpgvDeNeqHkG9o5lIPl4aOmGFVpfEla28fWrG
fZna7X/IUJgdLDvJjpykJVmNp6f9RTUu01iYPVUlKQ9GL7UA7Uklptmm+5qlDhZN
g6oQvsB9NSTMaKQM0jnHejJfIQOlU3ptqRpMJdUwMPkDC3eVIOx4KTXTVCOSO5bz
+17efY6DqjvRHo3qFgKeKXkBWs94/AWLn4MPSPCJ51GW+CHQBIuoD1W3xvZd6bxz
Y8lqCP1VlX9l9+0FLmblqLCtZYF9QUFapuUuwzi11XRRuYOLn0Zlt8AaeCqHY0Dp
7zE95QyZbrLSu2JGguDQXORVoyHLykhGGPFzVfiinRuuvGW+TcyhtWax9f1yO/Qm
pRoJYFB6LOV59x01UcCXJR9i72OWhS0BYxtrjib+g6yy03s9pQMNyRuW+tqM/grN
ZNqhIY2VCzhhLU4CQwmqQqqIzwjn7fdqsMWC1c589A7RkXh4l7xoL7k2ndbCIMYJ
C5d9DHvi6dANWPJ9DR+7EkqnTz1mzRvDbTsY+j8GenGiEd9Dmh2c7NfclyhfxHT4
jv9JVplbX9kxB19XIb/PxbUgMbb1FPEcfOlODEP0aXOUP5ypPKOS8i4oikkk0LTC
IyoFei/LjJNGX3+qZwEX24HnGxeACmXOxFTVwQFlSPrdumWg2t+X5XSF+cq1yGcE
SVBUM+Rt2Zp/vuTLlhWIqJzlIxoBGOsBQ/0E4qrCYg9QZ4Id+VXCykAqBQLUxnlz
ei7iZ4k8uAeMAwO7tlYCp/8iJzmXSwDyV+wyhB3Ysx1Lzy0FNYllKg6lsDUjfq/A
hIEvioGVC+Hpc53cUW4A8TeWMzS0qdqstMm9WKnG7J0JP06+kI1iwgWsj9C3mMo+
+tzkRTB3JVmtDtcKVY13Xgg33ZXyQKZiTjgbJr6BIR1V46bGsMwtmNO4BdMmXtoL
oVDORg95qKhDC1RBkN/cjLJsN6uDys6FOmXZikX9CNpCBRSLi/VLQS8oRMrDb6tr
Qca4OV1m88ebMHA0A8neqAc5SKtKlOI24IOC5tWTXG6XLRTR6CD09iPUFHnNkFaZ
W88SyfExTYf/FGFVvU4Wb6K/Q/k4Oh+TjgMiSLK8ZOQ2WQ/kYNUMlcPYM1EzwabH
s+idl1dRXO2jniFYVJKtduebKJascu3KMzhz0TDAxRZbg8iyVi26cIpR1vzjHFni
Fu7eWdEym7elteWyhKOwPCsPsLZ1KAwZPVsuOUOvebys5srwBB2sX0lnEflaEX+X
lLlgLgc2LI3A1r8UxDRodDjdJHLklVmo7jxzDDMVYsgNLJ7Uy7Nu289e3LiSqj/Z
ZsBrADWMy9VvDW9E9FdLB/wpPL3dExAxOPkM5CsyUR4HzEP7hnRJiBrX3z5Y//J1
zysBR5SkhNno4vtaZOLEygaxKORlvJmVTQlXRcuR8rsPCGbauxsDR58CCXHcTDLm
CX+k3yrGLgBMY2oZeWzvh6SKDqJfvO9xTZUZ7EJAEaLOa1ylEdhaCpO2f4gcIzxU
KXcy+6LCrm+hzfJE9lLBs0YTV+kC2DPB5yd+GyO5EQ3rq3H/0z7+9QXm5eYFdRrN
gerlhXIJ9133vI24Cy/58XxDMmacHWQEsFXsY9xrI+4Q3OdJm2UCtk4d03nRQmGA
Ka8XTbFkDnf1wJWX6rAMUSd9mbCB7mB0hAvGyQjffLe+rhymyj22GS9P7XLXMDxx
EtWkh2J3R9JVdB6qOVCvn5QTxQmjVF6I7dKYu8HZ6RjXYuPtc/wdkBCL3OMgN8rc
WsaAYPlJCrOvq+8NyLb9gTTusLx0DHFNkxoDQst7dRmYjbnF/oshMRI4mWuRAYYf
ea/zhWmxFYmNYiPVnavroRKctReKkMPcro5UFTO8alwPmLVeGzNNOf0Wy/mdHoWd
RTgQfbUPHt5VK4yCjZtcUPRLcblEHrCsC1o00Aqed5BXw/NC9WZl8Pe2r+QeIozP
hhht0NfQ8EFQNgdu0IQuQ5nJ5USJD7C2hjE2SOI5TfAVk5id7ro4Y6KeTWDUYbqp
CtvezMxU13ayyiJ92rL06IPMszELF5u6wS3TtowT+BUNhE6Oq4DKHzaZ8NtP9W0a
BbyjSCBa2d/dw1hDA6ir2e1uCI7naKruYXskamBr0w+zWObOvp8vD3UFNEOQa5AQ
DKmUICyKnQX9W6IPOy+p6gLDnKjkSWqjOGWBlLrmWDW2fmKe/a07X+1M5lG7hsSX
hUmb6fMp8p75Ysvo9pYpdbpoEC/3Daa5+ZiSY2vckaBWGDZZQOGaV5tTrIpAAQOO
CWNzFj/L+H17xzTkH0VysM4ujic21zXGqWBEwTHNToQk80Iot8hxucNznTpavevI
xtyQ1ipUPXCXVYpRq7hDSt2u9rU1/FbgZTHrOuh4j5soCv3x7pGs4zUWVK4cbdhb
2oNpWwyGzqX9NNc0hAeGacGelydR/pMpXdgdviMAmjG+KlCcVdbfzQb+iSMUv/rT
cJDTFvZBcVvQrj0/NObIEQggLa1S8UvGvs8X006hKXgHzRB+npCRSY2pWQ2MyCE/
Fcd68c2lJy87b2BscB33h/mKcEoigljhgLdzs98Aq+gSEESqURd7gvN0QYOTqz2i
UxSCbr3IZkg4JwVxd6PY9o/osDGhDWDweMBDIAKkplgTr7GC+dvoLaJHBntKYQk1
uuM4UR6FBug2oT0uTDNjwWPQwKj+6vu3NopsWoGnZ/8HvnNCdGLvocHLqMaOz0rU
IWVfyETl9C7VBoe6UrhC5SPyT1XqP4rpTwI4SPMhbWYOV1w6w682rpcOtmTty7XX
QnFFPkw9/DJJ1AqdWUo+9c1AlXrm8TI8AyZcXRu9RsciHCY2i2lPGv2CaUg8IkW+
Jx03OBDGzIYJsb7Du+pKBJ3v9hEzXdM3vOE8wX6DqdtS+x+CMRSZMdgtR8VVd1bO
zl9ndIjZ4/0EYABBpi0wFrCOFoRnRG7rdPJrmkgko08WBKpQzikb9o1zSC8iLcmu
Sb8IDl5q9xY64n0MxtHPgDcZoH+zYKZsuVb1YUmwMVeQknMnDYxIsEXXPpzKAH1y
7BNzDwrRgBanM0CRyYpzcnFwTiuykq3xHlYCWeIPOPQvcSdCvnumekp/uIi7CiEG
46Yih+o16hKib7CClQEWTjyJXVKe+teDl4r3AYuMqy2QlePJCpcjUN2B/+VHCKDD
exrT8UNpPRgadv/M0y6qi3o0OpjCIJyzd+aNtrUb+6BKDpEaAOgBRLCOlA3ci6zV
1FJ3DJcWR6bjV9+xLBHy4fqXzAI1rP835NuwBKUeULa8BqmAt/xD7+WJXpjXy4Hl
bwY08+9C4Q4s4D05aHjfX8Ps7xxT+MaCTnr7+NHc4fE+Y2WqojyLRIvFrtEU+wun
57YAleG3r75aqy5ng+ewnM29BDSdc1vtvUuj7ID1ongCErtns3X/e09YRKBYIM3n
pR1ev3aOLvXPseLKuLsfD8Pg+o/KJyHxRi5u5VhmqUm8WUbjwdseDiDQZSozyQDO
wv0itbXZbq6yV/wxamv9Hp8Sd1ol3uzx6EE0+DxX4tQRLS4qu95lPqMWHzUL1UF/
TcRD7J8YY43Y/tt3y7m6QKobiWpJ9C9kQyv9gzULflUrr4NEeSuilG+6+Q4VjtqL
gK/3aKd+Xwjcd1EC4ransXl4LEeeR2oeflMzanVD/fZif9mVVuNrrFGnNLLHuN/B
zNGx0Hqmul8V0YMyCI/d/vOTlM+MC5XiWdafj/Q60jLAyT8fJMgHjsncdySJ4OtX
gnlPUkdqorqmILY/mhV1+6RuOK0Ntl6b8Ls0ESnyYh8XNN/6k6nZUKTZcxHTT4Gc
NpLlsyiBJel1MOoA1cTcHWRtP7dhrWe153nJmq9x3I5AW4jRrygj7oWk4Yv7ZLTK
+OtdDJu9v3mWyFZROMDSR2clG/FEjMpBDLjPy3yGHamoXNC+mZDuy417+d3mlC7+
yRsh8LVmONETPuph4nDYNbuEsGcWDEs7uvXdtsbi+0GcuaIgE+q2pEekJgsF32CX
b9isiuqxGo2N3z19Mv8jN95WTt8I+ZU0oc7fIOsnE+E9RGYmdXRbEBtmsbQlbTEL
Zi1mibCQzn9VM0YUBO+qvDTcOlD7Eoj3QVbfP6+gS4YRHLtNW+E9gV4H3ipOuOX/
3JweN/gegdB/bcvpbSqH+fbHC3bkDkjFRGGf5tKadJM9BWvZdeshk/1Cw6fsnvi4
kh235nD12+JptE44m+AmOHjxYTFm3SwPRHgvDFq6GvwwAN/2DoCv5Zml5fVHmKOr
Ul0zKCgXojlceFCmzncFbnbZPT9mqBPayVYpRyvB+faiVSB43BSPSykF+zewd5zk
3HlJXCCoRzL2rklxSG0YmuTEApNMgBcW6fkIpZlrTWrIu8e9ZZeNfJ02MkSDuHgX
2GeQYleeOUnBrwp6Ne+FatKeUjiXpKQTIL1i98ZvdUlXrDGJoM4J1N+NQvox4FMm
c1Fh/RCoOB8Nqid/8OE76u3lci9M3onfl9CjyCu731dLgLZVnKwdWdfG1TmL5ReZ
974IfTRN4tBz9PWgBZ6Z4SCw+ciDW+Aaq7Up7OxPgHrdxw0sBH9iSMwaVuUg2WIS
ZDL+z4aOENzEaQ7OZXNGyghQ91W2uBUoBuSvbTXXTIGTWCuLk6Jui1tMSeHbDg3C
F0CkAqilqFnv95J1v9YffGazF9WfjmrVxTJed3i8tUiUjkYcGXRt/i32hWLJaYN2
gUBcDuDh4jOOB2kr1ZrDg3XjUpoVW48h1NEeffRXP1XIK0nwurVRIl8jntjM+aKS
j4+yqergbSg0Fx/I56VUPk+kf/4dj0XqpuJPYQJvqV6pVH9jeI8MkQ3zOVdkGIUe
LnyPXtwI7DUtYiZFE7XJvpCbFV+kcgs6X+HEF63cxoVzl45osQGItkQZ6cphsj1g
Xl2FF9wyruFcsqJQ/xQjPoSKP0b5kQOzvFgKmvYTHqIMKKVEYm2x9/P1KaRDFUvc
TfNyyqNUF8FBqk0B08SquGb351z3DEmlGtmIhtF8X7Z7dGARiIfq2jnO1eXQsqdy
3jiwsdSSl5QpsK9WkSt59tITyHURQWOAN3FcAixI4IqzYg6CpcY2ZPwsSkv4NK4L
FnQlxs0ssxGU9xE0mm5aDniCI5nUaEN/wOKL711cSoiKDOGHrwIGfQ4C1zTGCutA
tnhCAOe9eVOmUPy4NT5sFP5qk96Hci/79TgBbmJu8O6KoU2h8YxDcaNLTcPjg4mi
xhscMBdYIOZuJYzS6uCcJ07BnmtVMy0nDbph/4x2s/RAvCji5t9BJvgFpXKexFgV
+wkt6IrI8i5jhOl2MJd43BoME5WE5TCNvkDBK8Wr+r7d4Hqe48og5TUWQhg2op3t
hQl/1rfmq6GL8Y4J3OT/YSmADBRhXtMQdVuPXN63qY2GfQnwiNF2yMPz3oZxILts
U7SGJSDIVgGNSu603K1YFf4Kun7xk+XFV6P/YtL/3nkQKnYo+GgzRIu3Njm9bKxt
AqdOOVjFsdhsVA20Qk9Mgwvrf9IQ1p/W6JCaUxZ/UbPADhc8XXpENbaTgqIQFmP6
+aZqUPmNmVfwMDQWkbgoOo17oqCn51pTUXeLaSe2Ga8tqJe4MxlZAPBk3dTD68Pn
PiiXLPTznDAebopVjZqicHZ31ieWWaeY5oBzHVRhXzFyvpld9MAeZUSvSBUGYTFy
XzSrKMvy1QgmjgRQMFowKrLt+cDABgg8g7ZKRrvfM2giU3HFP3l86gz+rizxqabH
ZT2OdnPphxT6O8A+dGxr2TKUH2MQps4tVTGdkmXKdTIBGTHMqncYC0/GWnx2pGSV
Z82Ou4/uMddLsryg9/fzuRvZJPKVXpUzUJCWY7pGBYGgpTmA9i9xjJaET4SIsRFF
25OIoz3ZgOPcxq2PfcNwZZwf89rZDWHZEZrkjm4gb5LA1f58ScfRasUtIZjUXLp7
HdyUI8BJQfNLwEMbIHkN6TAI992HqnA8Zl95N4tBIz0oBsC+lX4rK4AisJDVydI5
Ku/AMGfrUAmHZv3sO60uFS+ec+K30fQsvlrtX1gFtKaiWnAIiG0QGEllyGN1uZqg
YPToYCBOdeIgsbpiwcLLHRFV/fDW5gc0EBrUWCxei7+Gr963VGGQbY2HAqsggd0D
wtSXZPzVg1sRNluCIR4Z/0Y/eMb7AHFZYMRrcr7AAoA3wyq/GfhtIzujrMsotzy4
3le5wLwMSaC1Bcs3TtzwYeeVlSbWfjnr/2HQiI/8WcDVCJghEjS2n4CQYHfaQ/CS
g9WVATQ3Hr5xJPnQJrT55YDIDMHl8UbknJ7/3HFynWZVDHeVKLUAd/DL3k+9AwVw
fNGVT5o5auBPkaKE4f2gmNo6sQWYkzxggbFZ+6BDk1AkgLzZ6BecXlhoR0WtgaUI
K0ET9DqdZQYREglTuIvxGnrT6Xx4zsh5dH73vZcpxxLifUgjTgfOeXhYatMT6qZh
2WPGrpFiLntMuceavCb/EX1qnOjvGZdzOniqMy1ofYNBOQ0y/bT3vIRmhJliCVLv
HWEO4kYznfaePi389MCBn+E7W4sDMBwtTUKpjXX9FekuAvNn4EulJGp3vQa3YTXX
G9rsFTC2x/yjmQA+se4Upk9VcE7PCYJjoMK+6A2xWUzPITGE/3VGR22hp9ve3Ken
RLSQc/UoRiygoVs+b/OMeYPrSKm/ethOFJs25YLQXZ6qG77PXarR1V3iE96JBmIM
cyC7H3zkGhZkJOKtVGSr4eYgH3Ke6g3Eav8foHwNVeU6onaMVre6YfpNJ9B7EcG7
I8oHtpbzrPptBDME7OvjjUUsJS5i42iAX54w29rLtuvURP3Byyt18+5rzLUhtAcs
cLrrptXbTd7jJwZ8uCgPNbeHb4CW9/flv5q4QPvKyF5KcKM44nFRS2fzHbxNwO9v
NJIG4apmBxeFlcvqAgU+UMM8EDXd9CMQONiVnlUMICDp7pF8Uw9nJ2xwSlEac70B
soWLwEPr2HCaRn0yODZrjSFWfmEEK5wpXMlPybcZKAveC9qqa7x6bB/IFqk/nzFT
xq+IRUUtLkU4VRBEJbsx88Z9PfpkaWWNlTISbc1w9qsdFhHEQ516mqW2gTUiXD7r
OifvJfcS8EmwZ6BEZOcbZgV0k/zbSD+InqpvaBSzqXFERrWrRAmAx/v5A4BV4D5L
ShTS2MmXytHZP58ugjK1IfOv5yVkXy0fWOeDi7FlbSLrXeR4wRbYoSorSaHXjrA9
pgWxS92uM2lOFDmmcuqs7UAflxiRYsuh6bVNZv8rlmPy47h/53h2TMgWMBylI/uS
p/n6DZ9qWFLnkWVORR28yoA55l7QOhD1BUyVnP8XQdGh2avlnUqkOIMCkqO3rDK8
eheERbRsdiQb5xERJutw7XPkaYetB/uYqvMI/8UHZ1eUpRAXRIyT452uwkoXTgIP
TtmQYEIhwSmq+GirsbrIGv8My8IpZvCxLewfKbUpxs9qfy4Juy9V3wB4yxgkgfjh
kqO5qTrDmB7/6Eq/LfLIAyxmtN3WmmmzfOUkUYSe+6jWNJcoU69gIBBfWUjPQJ4o
v3ZC0d2ExwO5WDchWk91MMRCNijYhaUz3lS9IREItBzVniWGxye9j0vFGc1aj32V
oEparz3cd5d/l3ghajw287AJ353JRLPhK7v1JI0UF7AEKH9bElWo0ARuKBJb2zeQ
KwCfghkpybwvg9s7mBlOFqR/1fI62AeSkyqSIzHXu1+dGTWHiGHo5WHNkAfAiuBH
YISKwJW8+Qa/64Lwt1Mmjjdboqr/C/l9pX1NkmRlvRSXfuqqh7Z0atbu+tHZGfYl
XjuuCu5MBr2YS5wSzrCgh3VZsOQ6YIY/WJFHtZXJMEMMm1f+Bx4X6DLc5kR44Id5
5Ike6354N/El9UJVNesYK1UR0mmionZ2A9sNVUf3U/xc6+wJoCJJH4VEoA9ArWm2
gErsEeG5plCklyZAnc/XkYhJhsVXdez3gEr1f01D3V1eN5Tw1KuwB0n+pQ5tnXWN
yfNhrEQexdv5glvtXwBRLy1CPs3ZIl3mkd6J6BO5qvvQmPitdm05jiPQbF6X+8Np
BgV4cfmIFzq6cgmxBBI4aeeGVy8wm5W+lgOGiDOWvfbE2mTuD1t4Wgr4VSvPLOKs
/F9yxMMnu3+bVojQOHWLvgHIrzwdlQjuwqygtemlnrnXMnGUZ8mxm+fJvPFPY+J5
US6FAff8u94YrzdSIrjydk+yHxpnalD+ey8SYOWLwtnseeyMrBndweLCaqHygZuG
WbJvvcBPre+7KuAPBHTPbmp4NCgu2T+9nqLeF3t08jY1w56ZvIPLq4C5GGXD2ukV
y1WKfYXxDzmMnX1bZzQnig1OHAuBCdqTcYb8t4Xfa4nxqC3dBTfpCZDyK7yvFpR3
FO+DaNml3N6jS2t/QbmruzWxxaoiKsc6YTOkZX9RtcvBc9wNWHA1NbsxlFafP+r5
PvpSsaUS7fUWaX4Qa4RZcumg+7Gz8vJcSY88D6Pvw8T3TyvIlmVG7USs3Q2HeMCn
q+OuWH7ixTCJ5nmVbYxHMsFCuyLm6M7v9WfmIbHaxHT+it1hZUnc/dJABx3K0eo0
l1omEGbvbKEhKdzLXuxio+0CLs6buDcxROj7u/s3eobAqSr1DSYmqrvBliYwQpMi
OXhnmEysphBJvuN4amOI/1tTt/rRCxwRw06fN/JAJ5fnltkyIzrpqhINKdNogxKK
/vDC+oi9nLJ7aCM1aJrAll/Mym8u9jwwrYdzHg9/BBT5lwskqkPV7KFGsWF5sCcT
VJsWGwZSnTUMG3ERjVU1gzOw73Jwm7QqVQMhKvlV2ougBzXFkfrTtb1eRDEtH4l8
Co9WwQHZlqU6jr9xuSfkR1Kg0s57hoHHS0i3147aLQHb4YlFWpzLsvr5P6F+kMgl
KjgKhO1MVpmD/sXl+SXSoQhOqgPfDu5R8SHaKpWCm5Xg25I6yDNHkEi+CrBsZzzM
3t/kKSOf5NJXsyXfitBgsO3Pn7/aKz3r7Qe1BLBRiuZjFzzFuNG044yVZItvZ36h
+90Y9ebFIoh2cRgCMla5o065cWqgwSOSNxiDRxPXyMzGGYs32vy+NJdM/MDTBGyK
1GUyat7iw4x78nhSEUoNGO7s/7cEy1P46RhnWVMcxgUsGaorQudgrvYzuARuqZvz
9JkOx5oZZqQKD+RE476ETIzR1wvcoOAcm2MgBmGMMjnnTlUuY0PFUaeq97lOHrI0
vBACbnAsVjlaF1fgNWzgIAgLyiHZ/IsoTZG28ACc3swR9TBmWWAN1TrprPU/YkIl
HxfeajmPaKL1KcUcthj3/SA1vN4hfRQOxxbzLj8ASCot/Cp0/KKPOzyhU5aLooDp
g2Cg50+aqU/OHhcZO5Q5BESTUipQ8wOprnA0fPrFkMe7NW1r4RoBRIbVCGzFiZog
TTpNzuDfbtucoNQ4igpEie+0cmODHwDZnvkXXpbCE4ohIQEMl4IFRfWEUBImWrrP
muzlFr34qxUbQUD4mqie7MBnUa03Cv+kxf7MWQAIx6XLYRaddej6bAfoP+zHGImD
KMsdjNMV2YD7uh72CjVov1pBJnQjCDRjktV12nueKzq7IknZX0Cw+RUv+d4ThQYC
y+T+wxW3OdiUOR2gcNUgGBffgEbSvQD5uIvPO//hTcJDOe8mW3OPidiPTGulaBfK
tpNFSeMX+Rknw2fiQhf0X28rGwe4pJohLRAT7E9QHE+nhUAAVAv1AEBbzrmFbuVP
RzIcztb+L9Ep6T2OssPYBb8H11gwZL10wPA34Ga8huzldhCDrpHqYqxw4mmZr8ZN
Z25IsF+3dLftY3yz7l6D2kqHN2yjjwh4PY8m6OXWENSJf5hIhUVU6BmiFWgxkIdT
g+Yp5LBABnzctW7NP9AYH9TjGwubooYwQKrmUEOzgXhrF6BpSAnOgm4rqR5jWSPd
XnqIqZ0tQltFOT8OsOqj4+xAI7Vm6BguDFnwR7Nf8SK9tyDPcyq5HssPYqQCHzyD
CP8MgoYNbxJ2q2JxazPrUR1CRkiEoJUyu9pt7EfGT4wv2ia9feSsP0F4J09MlrNf
X/aCgJTfSORGzpZQEckaUN8wClyjH/Lwn53UPWgBau62nAMv5jg+Qj33fMqTblkv
x4tmp/ejIGDiqtO/kkM0XzmwrSJ863+JtaVg2v9wZwc+ME5W2uNx5sx2yCGxdABj
ci8dAXPGLF+2B0hwihcrjszbcTHuN3XOXSuEFyHncU00ogv9Hm2Essbf+ZT8UeqE
R0Xbb+XHbda0NNMD+tMsJgG36BeHopcmlloi8Ep2AkK9gtDje3cMnMApkPmAM3Gz
pA/y4OjZNdXbx1murJFcPxVm7BdAMp7ey16k2WCOEAQIErL5LQGvcs91kQHTEaPf
ikZULBrX8fq6Wi5wqgHzcSF4tCVwZ+F15utZ4YoPxFMhjoKf478eKSbE5ZcdGD3Z
b6dAooBaymKu/LthUFotOr9xJ8t962ujHtHd9M8hrNavClo8ruD6rd7qY18ck2oM
/vZKe7x6PHpuclOx6otWrW6qu9Fr+UNvYr26mikjy+qlNi7I4rwtMZZQnEUPImR0
WN108PaFkoaMLaCBvrENQC6br30tBvr6ZiQ5bs4xUQtdSMsbwWEg/dfT27SczRpg
Xhn6NDHKAlImZPuXVUPckOnnOS6D7eW1LgfpqFqWXf9kqqyZbGj+HMWa9k4rqUIg
V7K+ivlfEa1IiJpwvOjOu8Uit9Ga7RR+jgISlhPifS+G9BlxLKcEV+CSswX9UeWb
eG/okDp3K2heZkwoNX3GCkFmZTOFcv4+2J4bciq6esUYLOIHWax6Wx4MPk41qEOV
9waXqwHTTikoid43lEtmeoGO1cdjHztV7Sr0JQ/rM9kdgjC0OOa7R5+FmEZTf6CZ
r4ejUWPuo9pCHcORVa1bOL7ovh3/5JYlMfWdN5qC3oQ6OfdV/tMoc5VydfjnQEJI
CWU3whmH4Yn1UJcUoik6pVfzA50aQFVWF2cYG7hOTmkekse9YG21OPsnlEZM2MLK
/UjpKn3PPiv5ltMwsFcUj6dCEcOfjTdeOvGdj5jloN8tK3eEguy2vUMABcOkC6t6
uVTxJw9SK+cw832hBBVpzCReNoUvCJdjHfRMnY0X1349TfYM+wyAy2K7rDIarhLa
+9nZiBAtULZsiRDXQ0/sArATPNBu1lX5s9YZ8HYCBiMurLtvpDx4UwN6H4Psw92l
DdmRCJqDRUiJ8Nl81WKgUgRWHlKd3pM0zYymUcnyRwFNJMLum6qxEkvlnTyNyFjG
3pthKYzfBeOAXiF+XvaSMyC+4nsHidCRvk9HH7hOKdlS1Pk2Ttw4OcLXbEN2sXbY
t/+ifIgTbrHs1bmj1V8QO4hDKuRNk6SLzutxY0UVy5JHw8cra3owfB6oTI7ATPLJ
f4elfKlvGItOZHIP1JEwyfA4p7XUCkAJp1qNzn5Q/9/itD9cG/icJ50StrFxIIZZ
HKx6rQtsX5jzIWXtCvvzoKnEsckpVGXmnhu55CTf714m1BbmZUqwC/OIT6Ak9go6
EUn/VzEze0hPyF0qCMhXJYpDnzfgMSidUMS5owmuWs54ATZOP9hrXs8Jjp5pZopY
bekXxwDpH7Nmcrk6IiBuiKqZNB1xvr1GkSfkuGLgQ6wGfuPPT2Fbytqvyjl+nQHV
C3w4ZjaNzP3ODs2J3fooCnbXJ6oTJntJIVeHSOvRmFfDrcVwla0iJ3rOhc/7UNGP
gVS0rC7bgjBDWoqT7vKLBuGc9ccGt8zoMPIyQfF2b3ABM9UXUHQ2Pnqu3b/MV7FN
afI0KW5uR0fUHQiKErc3BAmbtsNI36QY6AKdtQFsnlRGDrC/Ae1jZ9VvpOQ0RWKO
7ZmCT5hQjdqOdH+VI4jRWygmpCjBX7fEqvVyAQGpTKanArqEoBZbE6Lu3uH3KeSR
tn/5Y85+yLj/pfvUCGB1C3DHiPnk1r44sQBX/ynOtrenZ4prOrNEvQ2gz1IGZRaU
SOsM1suB0H60MlH0P8IxrzvBrM3NofqOE0TXQhHeannQtik9MJeESwhMM9vSRj+/
i5SBuXveNWXDtb8ElLV7kpqh8KDV5ln5bwP1gmhVar5zOYU5eRDWjD/07IKuwJ/2
fH3RvoNbO1e155WC5iXTRBLwUNPCeKXwxwmspOd1CfAgDxgScVuPlW8LKTj541N2
xIrl/t5xCERscr0xXMsheDTOIQmeoLjf8EwjoteH3E0ClCSzfRiFa8LIYMZG8tiI
UOjbK8yzhHZ2C4IXBUnR5uXutC2W6asCi5anHmJMyTXUGF/4PFd2xXyBWk3FOcXR
44gRDNZANyOzHUe8sMFlfrHYdjxUsmSivFuLyzaSzsr7Q2CQ6V4SE1gtgkAoteJC
kSE+hLnZeLqWzn/q/coQl8qUCppFSY2AhVH6Hyzp4zrikj0JZ+JavgS6zRjISwdr
++MyBBGC4M7H7KsDIOhMTLuyGcU6FMfjbhddKI40lkjAZfA3g1daxy0+82HvI3AA
slmzpJFL2IJ7SApEqZaR1WS0EVLgLozAHMJd62w+RpObgkkxY8hPc+gjnjgfq4t5
DczMtLYnSRss7qLrxboYC7023lh6yFmXpVZK6/KWPpRuVrilWz7IYJVCMFFIcrAN
NckW4SKSqs4Frqg/rz6fPmktaR/L+Jk11kVu1GBBSxI+4Ph7b2PeqnuBZqyFfLEH
1E7suOM0KbDewrWNByyqUxTe2qbj7n+VQlXxlp6DwCgV1kTofopHOWOIASFMtSA1
IwLoEa8U2q4V1xhP1CEWWVTQafuTb/yN0KaYPgcktDO77QHaRUAE0FPTgk8xbxZ8
SQmikwTCgNCsNepzTasXyg+pITjCK+kSbRIVM8sgQenUBhCvt3nMI8aICiU5ftKb
LvTE1wTrFQUkFnM4/d/0hYTyf9QKyzLCM6n1ys6aJhYhLv9p6fmPA0ge4QPjR0Ay
OpCHJCVJ3VJEsL7ncwpv7upm/QBCEgkeyn0c4AWU1ocP/EiBBNzKcyq3k+bb0iUk
iDTAayTpafv5JtZp9zPIma3e+Bxa6c/ulgxXVvkmO9VK74wvgTNMVQamnD2KPPvd
s8qz5HSkTeZXwNQLQZ04ZNc/UR4diPlQQ4kB+yr3V4Ic125uvCXyFAGNKO9FjLR6
3vVyxBWaLpNO5VaviPOCq+BvJh/VwdXa9OJXfEGpP21iybBEC65/ekeozoTgPL3B
ZMI0pVrfZyAd+zV7TVz+d2KIf7rtLrsgoOdEI3JhOJeOu2yeFo/1ex4hbZIZyiVd
ixwr8mRU/S2Tfz6hbJRcRzGxCV+wpMAkzJ+kbAt8lWddgq+evEV+Rl2b27Gpubbz
hQTYusMRdmsJkz1SdzgqoPTznNz6wrcfMV19wRrmrJHLVTzjvvrpkSP+UgAGSuty
PBfslWi6H5Qx31gIxDS9FK6m8tg2KZX30G0+258a+BmWZv++ScsjQwHAh971BSjn
6odti7xCwCJDUT57EbD4TcRBX/vs+41OwHw4CXweujyxHwOEhdgDpFaC/zDxPgT4
vVHOk7Ypgaz5n2WfXq83FSCBcyadFYfylmSTj1HK415LLO9r8W4VITsEFT0L4QPs
mWrRVLwIYTEl+ImVWpo8t0InLapYl+CJ7qquSt4ObXxAE4LXF2SSd2unHVNPr3aH
x8bC6RUqekqOb/zIt1+PFH6t/tehrISheFINo7lEwkjAz2llUzRNbyTLwLvh5Ffz
JQSwNfQoW7SWkZKpJzh2D2MqjX1eE/hwc4EpiFonX8k+pHi8H01sfw7UDQzP3RsF
r3S4LHMiccCqq1cqr+uh0vD8yRpDYTEIndlHUfEkgfTZRUPMNCMB26GUL+g8ot85
oMuBCdsl4COSLjuQ5R9fKG1XR2zUSih9DMubqICmdqaq5K9L4O79u9tGDjt2ncPA
+Kycyex+uKpaujBbl4OZmPvEPPYjSTlcSydNxr/r+XgyzTEyi9CPwNBUt7g4TNyb
XICsUKakSo5Creng08RnA2ghM8mopL6Cy0WBit6INvlVr0z4JFKvSWyOwaMC24X2
JoCClHYT8cb+7fz7XwbpAslyqXSoeTarqwIV+FoSjr9eAczcLIYHQhxt/vS1/6rV
39AYHyuTCFoQzZ+gCqQfdDS8EpkoXakkQXmTcojhfwL8Bufy1Q4K4yDk+xI+/glc
Os0eoPQ5jsDWEV+sowiAZJfXKMrLDr9IpeZmsYk8fuZ1W5TMPwbIufVLOpotGXDk
54KMyhRvVYXjsgCKZtPPJfUj6t4dEJyeqc/xsPMJ//1ZTEs+JbLHTKqOUgpzXZJV
lagCmZvSXRbPx0udEqff/jRIThAXhPJsMHV4GN8JxX7gmN88jzEX/EVfDlT/jppB
gdnpbchvfpUh3hpx5J46k9LpX9jm4xzShLnWhy4z6rqKYgLSK3HSm+frb5H9s2DD
IZ1ciI1/Ww782EAijNPZiwSK9mADzxbXUDSp/5OSU5Wd9gPpSTHGVe0bYY9xbldt
6ZpIgvX2CMGwJKfmfFhhEBHb2RkhXBPDerVBIB1qJLYysMIeVk6g8AmgdCCyQeV5
4XIXA9ezPmdcKXicK84e+aBOqNX2lWILhX1dJZkAeRrY0djW/V9nxKYtSn55qlvB
IsVOwNrHaNhrnXAYKx5eimPZuFp+3T6k2EXdnx7mIj1GSsz4QFOmFvaFn61UaAYH
h/REWrzXaazsKWUdWjpEUNanlN/o/fTAuQOR+9sjJjRka14UpxorhGt2dT4ovXbe
DstoGFIQWuMkPwdJAs/7F78DEV24aI4C14buT6jLr4rQudjCckDOZmhwBzwibXJl
3pFTReW67nJvFpvEVoxC7JQpiXDAKXjvahKI+N3ZgQaUCMdXlYjeQbqtDGJ6m7Kl
/b/KRcUCJ0u4cgCob/e9sLJ8NP9rBuXMANA+J4OB+4LE+4oDvvZRaDPse09Le/FW
WVqvTkjFGINv7TMSyid4Yb90pmROJTRNkfTvLBqvj7QgvD5ZWrxiU6mW31ccDo6I
zZ6BFEZQGwqUoJJ2WL/AqycV33IxBCkrOodcPxq43RMBtcqOcpN6oDW+1PAxvFVh
YV7WEA8kZnlbdKlQ0wcA4bDP/xyygc3po0aFrmIfQ0Eo5pkPKzSopU2IEZNHqMjj
8pQ+xsddslge+pjQNwZ1LVSWMkoPh4m2eUC0mzwDldNIATUrL7o/F1gtLIMrGNcm
345QnYIs6VuKQdpNGfxR5Vygekr6QpAC//y+m3buhGM+dkwDzUaj87bSa86o6IJi
kHxiFnQUdSl9n3TpbC0LGHmBkjtLSPXN7uwOFqSibwNwUuJJtjrrp82NcORpd+G6
9UOJEiumZ6QpkV81ZBhRrAD2Na1aCCKx/LPxSzV1NeFvoUy2w6ZQtD9a96TGuSdu
Gh7JzQdjlrJiutDTzSt2I0/r/Bbs+SiyE/ldY1rrwT5MxY0M6PksW3cDsGNZFBoc
ZUOPouJHpCdW9sts3jhjjljINzYmbrqPQ9PNq8jCy/GsZGmLoy2gCvwf+//DMCyo
17o1dJ2ZDS2EGUJU1UpTHpiYh/H/5dVwdXORT9pQ22XfN5PUIikHyoFv3UhBLqmc
f/ZC5Xq+vC2r4Il0RxhOtyDwZycLNGUgf2hVIwuFGy8lp8i3utPPAYMGyb6Ky1if
/CasMAeUijwNUe67FTSt61v+XAGhGPDOxrEuS95R5txNYhCWuULlfuB1qMQuJa0/
RxDJtMCLeQWsNPvpLuV75JU6ErltnYSg4Zm6QvkWu8Bp+sx3fUSPAmt0Up9xKXog
DhLjkxfsLMHLGHXL3beQqTGLWxzJ+lXDuKU4rK2GtlEZ0tptggIqv4WTkQ+vgg0x
VsK4clodn+rACkFSNVlZgvPD7jXob2ItsJBMJmGJibF/cejvF3fSx2T5cj+tRqQo
n3vF1wYDmJMkFpYmVJ5wnXaS1ZvAxHPBIvauptYgsYHLBqEif0F0wHK5rG8DHZWf
JtNOPJC4WEOwDhoizqKuo+28GFETkDpvA+/EJGJgsh5GJPkmc/rteQbdG9gT9r6O
B1JhsXAlzUmROLuiQZaeupOou0h6L7I7NKcAWq5Ktp72VbKQ5zmh6fL8E1ywe2oi
VqP8r6NHj115ga19s6mjTGn48v+OwO7FE5mNBI6v8jOZAIl8tTrZGa5kCZO9SFDM
rx0MFNaBZMY3WHtNa59uJjmc0CQ81h8bKp1tWIZ/ea4ZvKpgXrLo8xtSjukLgtv/
osF+8FBsISWaCYclV9e4jvk2RC0D6KFzNwTTr6+UB/K3njgEqnJu+O7jUGS4XEoT
UyyfORgnO55YvJ3CF3rJaWvPZ4Ochq+z39VtMN/cr+j7X+UqO3kNE4PCH9C6QrkH
KA4ISDoegC9iqZy/bhaGpfgYszW8pWXPZs4fTXla77wKjvhxa+4E+Wu7x+QBCgCc
chZs43xd1Be6cuN7g9LWXjNXFMunCbNVtbGvllt/yZgDQTzN1ZySYTMH0xF5Yah2
SdTTZm5ocEwuCXpDfWJFwjnSSM7LpXGkN33CNZjACe6aLJ76eFW/WutZ5Zwnpz0G
3RHlh62B39luIVWkAZX5or9lqgDozlfSmmyYDEmKqX1W62Gr1B/gnjTLo6/UIyKF
AwG8G1jQctkto80qi7Z9UoZ0J4UZpqn3iPOqZgOChAoXEgE04RqIw2pClpCtC73v
jTLLU/tjZwfserwicinZdSSzvn8kGrgy+Fa8dmk24BQODtkscjfa6KUe7FY+Qbpz
F2G2XGa9XCPrSVSjfplZrtJo3QQFn2OKnW4mbDjkpkPmF0C6LCcdpOtsZxP9VBXN
YAHiwBwIjxnYQV0tEL7px3mCv0li1pQSqmU1b+vReDQnDkwNvXYGne1R7WJ17/6C
loLpznW5O90EmzRI3PJ9mM3a2JNVPFgPz1/Gh56uqAMFZ8jiHUHyw4L+GIXy87mU
LYB8Pow10K/e5O75XzG61nKg+V0ebWfIdnyX2LcOMVjnqqKIbydhcfuiXWSWcLYM
+glXcTGXfN4Jt3iuzdF3r+EfBDC9LA4DxM1Tc7ehGGrhDnl7RUC6q5JU8xZkUmJJ
Okc/xeBZYrNp0P6q1693ThpBbvfxJ2zIdBr+jLK3SMruiLBN+DEhsvhgkzFyJUhu
cV1DBlovi7VQ1SJkuQO6uJKT95u/eSX6/Cb9vzEztD/8KOTaH8+Nz+uu3avxmGS3
EgSMM/XRyw8Bn8sSQV5rk/S2utFo4/b70gYq3PJWNEAwOyS4Zs5d4Q60TqNUp11o
KAJwkhTC+v3eyMQLYBbB+Cu47Yiwkm0P2ffm+JG4QqLTzcxNEo91Q1bWmULnZANi
68yH+e+aawdz3ssEZXK20apOAN8suzYxIrq7CpipYq0P10JyXeNTaxbts6cQ15jH
eRhFVw4oF6QiOUw5jIBJn1VoTXJItXaM7uvypFu9nNMDH/veXHaYt6PCTtchYuy7
Zsj5sYkniHbidBofwx7VhffgPXDV1GKytzzhnVRz9uza8P3zmlPrGkejuHD9bYEs
pcc1v/sDugJVQZErgbUpgPdG35rw4Cfy+tSLHhCVZnrFimgYJbllZTopoU3oHHqZ
8B/1jTO9Ed6ez481AIRFtErDK+/cp3dkQ4v21knqr27ctkL/zyQDjPEXYXwLZD+2
g9fCtdYx45dx3VJKeE8MIMJHNQ9COPCQdaNN4nDYxuxI/mZ/rlQrw+G3Rcz4GKFj
OmLt38zyZCzLL9Q4pA6EXKLPNGCGbg2LpH5vU2V5NY6DGGV/7rLG6h+hF2+EdXMl
Z3iWzs7BpYZMNCtEZ0+5UotaZ8HKb80+uj7pp2XBiliqyG6s6h9I1zKNiHqy++Qx
x7yovJs1w8P98EJ5EDFr7YwOueFtJY6dbZfASnrQrFdkp354f3QgO/tNVPpH7BKb
fABEWCSZ3eSIrAol8KNXx0ZAYKCUVpmz7xPvCTSp5QA+MDy+/gPkmSzizyO6bMiJ
Vvb+wOTJXDk8FIA802nFEdLVsAGEPrJgeO1kD3cHtnVNG9tEtwCQPwZ4W125a8Yx
qmsQVd9M6xADQ6vUVOUljJCUHBT9BOKh++L58Q8QtN1JYsorT7VTBTtnd3dCuR63
Az/BLhtlvTVscTMfjwRiqxtLq9ygrD19vaoDMQXCJeBoAYTfH30THQFpUlJaK5zb
xyNkepP9Pamv18hdZTxbC1BGDrYglViiE1v8vZBi7dOjdW6N+3GuELn5h3Gb9u7v
OD42kU1dQw+D0dJBBUjXUrYIFMeeyDNxICsYtGc4riaw6Dg6kVDZa+vdXzXQa54z
BGFOyQy8r14hdA28gckhnb5m114Il4jUu23oeDCIAqetfMhlZxhDu498zlPSjY2a
oxuFZKikaZaua+0w++6fICysuVg+45zjFl9Wr/6Ftmz1sfvpeP5Wa+iuUwiRctlR
m8QriMUntmm91PWTrRvVCB5G1bHU6HmhuSlmDrn+UuDzRhsAm4pqInCrt25D2Tvr
L1qRufNDbxeyABMrAno1wToTsbzfhapQUJc5oFf1W95zEw976NvIbC2b7HqRR66h
45iAWChA8vHG/Y8H5CHdcEazAlM1nMghFJy+DB5qxj5/UHBOzJd9NJMrBYI+87nV
tZx9KrxPfKQuFYFZlH3fJDGbV2hn2Yc2LRAKLFiLMJ9IeepYEu6nG0PGXveLI1Ja
Ge/OUPbnmBJbfaVW0DFq12b3KKW0oq6nrqoTV7AP6XUV4mjjLTPN658ODJh+nKwH
AslB9Asd/UWeENQ+oAMfkI/wFN3E0i+jEq0SaVZP1HARepYx/uiIHjuJNzmWI/Oy
Gab5mIxzOeek0eSWBBRyAkgJcZQPUjtyAavgX1arTDYhafmYtqm5glwCbJGoPQX7
Q1kvSEn78n7ztDkqhc8OMuOQUd+9c9pi+2pwmQOw/2PRO7ZLdjda5yT0kJKPs/NV
zCKe9+alc+eJ8qwgxVn4yoKtrg+pbW/9ABP99lOxei+gLfnIC8JCukipp6Nqm7Uq
5cSxLiR98UfQk8M7RBg49h39EpWmIoBpEq8XVxqSalPgusLafmH5BvOyX4qBTlKE
plaaQw/qSN07jUe+aGYqdb/DvBte8fcZ2frWjTheROdQL4p1yByhXFpkUPE89z0Y
I/u1VBMuv6uitqwg5KywynG/j/bZCmVw6fhHpb2lMP7KcsSkRvOEo+wSGpe9ufXS
c1nMDLnBYYoPTwo9IvfSN6gswEh3zItytd64E3cVDEVjZS7DIxi+W/qU/Yzr4nfe
rSgr5BSFZIj22iMp9HLZnwSTdcpmKDt3FDHz5BJ96FC3Dn7D/iza3Zdeo5QhGadP
Wq9Fc30fZ/M6ILW5GUsUnyLnuT0wUrlS2aF+QgaDpe5qUrLo7tVfcn45rPKyDK3J
UZl96FM/BOX/5lDCjTcJNN4Tk3m33QvWx4LCVf8OhMPTUHGMmZEEioQxx8WYRJIQ
6wbruzNRh6i81b6/Vla0wObkOhjeCroXDsy9+HyO/mDU/XVQRNnkgER4Mzwftmp2
NEOVP7eVMsRgNCtvFjF2m/xxww+csFZF7X/+Mj4JGq2O87iY6z+s0EcjQu4EYEFa
gfy+5jITbdOSf1ZJ0hu0R+YjKjkaiuftk0eDGRcaftN2+sErfU3VOKpqfcfzxSlH
ol2u+IyiAMnSfWbP26ngItShs/ANZhe10V8QP+hp75W0PfnV/SF9oLtw+6DUKT/2
DsL8jH0k3RIiuYuxvnW9P98SkPU2jhDmTU5qtey6TC+RGa/4M0Zev6Rsy7+DN7Lr
bwZSI8c2JW8Haoth73BqSeZdIXfKKhqOUqzEIYdCJ8c699H7CKgUKlxh32SLi4OO
CRt8AqmGyHw8hKYpefyLyVCNEiFoi/dijTrfwOZwARcsa1gSW6qPuiN3XOqjZiHQ
O1D1q0SSpAKfDflb0OoRop5Rc99dzkfT6F4X+KSLwj0KvOqwmhXgc+C2hZ61IpUo
s2qjilMPsUcta0e2MZhIA8x7S+gQLk7u/IVoDw1cPJYpfRtVC0oyeLofeIOE0e7J
BHiH7ngmUaM/EdMLNT4U6tQN1pPSU24wVvdKB2kRNd5lcu4e8c6GeMjLQpplvLmF
ab0TDx4fqKxFdMkx+gdUj98ySOpnewkeWG6WEQeMGzYUgJJ2JfPzIDE2plI/Vrp5
Kx4usYOMKia5pyn/McyeR3etMa6plPYy0NootzgNwbrx3WuEDwvxIfyshwGYe/7Z
y/PPe523ZfjLWfT/u7VJDiJFgQXNk/03/fqcmTserq6RTd4lKvCC5KmGNM+H/rY+
bcXtzjRPqgpVyew0o+pYtn4jUcBjYPd0iWBLDVRduNFIqhAabuMDu03s0cY0sTWY
XuEeyUiRjGcvWckeC0JJDBGN1vI54gqg7Nm3xBvdFhTdKJrC3S/IADaUFC4Fue8d
aqysBqYbeTe1oxwtYZg4squsIKnKp7R/p3d04AGRKdWSMgBhlgj8BrR2KPkubEaF
RAs6RsqiYIi+BdcAczZCEeMTZkgnFk18AFl2c1QNetbAtYEXVFc83uVCe7oXhsfE
oU4T/kl5PeXYdw9svV8KTf8zmJg3P1nZQ2Rg120fkp0GPiZEyEcHepEdlpSKXaZ/
kq9HRmsu6SICivVIycKICrR0AbDVS9JkGwqwoiWSEOS3DIDlHmFuoPAvcLiFDZxw
FcY1Kiolvctleaw1w6jfzndRSEQ6Gd1pzYGphfp+rBubc5HNGkTSUe1nV5A7WGkm
2YQDI1DIhZPK6D8HRSD3ligo5T1oneTlSC2MAhKcoAhv9dT08ZC46+CMJkTxUb9P
c+im9Yu3yl6wA4bEKO6gKtXyGUF0a/BC7bo6M43BElJHfIIEbH10a/dWQB1uzRu+
DOC19UgX2IwJzUtDfuUgBmoILj1oz3D9/H+llvn/h5ElUdiutMFjeCOqY6cznkA/
Os7NxTiT+sXJAklEN8RsOOIW78qV9L6w7wRcM2WsuDqHsrsCTOY4H8K4LtkDlpCV
wxm+mEaxF7DzlLSdlDhXoOU2dBQ1KdabQz9qdnQinC71rEGPdOzT4qPub2aKkFMp
+m/JxbO7J1Fa7qBoMe6Le11oNlWIyXzbAu+uD6xuZvOgq6BWm+4zPgicnN/UC4eK
w8cG0sjYhielAsE4iZ9S7Oz8Jsxe+ID9MI5bRuDmXe+B4sNoYPrAi7tay+HbZOiR
0UlWcekT39lGkPhWNih1G9e1LfF7Y9M6prPSxuakFmVhOyJ2Wp1zv30pUA2ouFO7
RgPkUJBXD+Ey07pzAbQ1zpp4T1q/EGDIYq4dmGVVYXrx5ZelVbTxCMeMLcC9TGcX
Ame0vS7A9qAsyntc5LQTm5OOpKPq82tpMvYUJK9qSfdXatbFaNn5/seZB0Pna7xs
xXx86VAZnyfu1OIW4TO4E/rvwuGYI5eYFL5ZstSYpkrzY1p+/B+uE+PLsgXDvGea
48bhFRmcTJO+R5Nv+s23ZENPbZlqiDuVvZ/XVA81BgeItSYYs3hxoVpJ1ruTIS0q
Y66j7VF7nkIAfwvFR56/xIj5rIuEDFxKitz7steUVvUH7wMT96S+o9U9b1gEO9qc
LO6hRRXc1oPIyVPaX8akx+gumzlDQ6zMK3Kc6wa48PbDx0nmon8N8DGbyKT7A7TF
lAaP27hqB8D+O9fRqkXuLn4x7j+BKNe3bFKS5QDGw01u+X3a2WIRruo8eIEEyi04
cKvVkGnw6xDPDyfhCJ3rbfosTym5nznlR4W4RZVNM1AwIFWUe0/0cVdaG0QiE3Ky
ACCBpqLDRf4apeujBY7N3twkHCPJUCsRNlH7IoH1Q7ZfZ/KaNz9a2ihxPQxMHft7
ydBDkygC1DAq1zLVeVyBjERo6vz6fT+/sJkO75ruQmyPa8Bm57rHlghfCKTma20A
KT6HnAWkWe2V7l0tZCZNJNWygH9L0Ofy2D87oRmWXqwXcoLtSklqaNy9/EsBef/a
WBldkcUYSyIbtiPsJYuKqbzignSaHs67IZtcU50EJnjnmfEe1WbjPMkSO+lkUm3j
BTIJDgn+AcxPd9lJ5VnPkRKxsaIiZjatxXKCP4DtKMxUVGLtIol2F1ntCwUAOOUm
MtNB0e56Q/qq9eVdv5sPjmoCkcKrZwhL/jpGKSxiqaYuP0satM0NrnppxFYEuuY+
RnSjp2ewrJfbskw7GkkKxSAV2Gp7PTythtpsuFk2GzdJE9ngw/5QBKgA0cbuPj1u
UPDaf24ndr6ouASdS91GBw==
`pragma protect end_protected
