// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
svFqf9jgA06CZ9/Wcu6dKe9ookDz1tSuvkR/LI3OFKmo6MPEtHQLOrUxsFuo943F
L1rbXTQFtBvVGbvGbY5ieNei/Y3Zf5xH9lgNcFREggs219xIKk7+ZC5XuYqgGoFE
kwII/u0vqxUCG8EjvpC9CGgX652nsUj+Xf2TcYel7Hg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30160)
zcPnaWNTYlaZ9I8/dxl/zfPz/c+K7wz4TS1aSmqkIwXmqN2NYQ9Nks8E6PER4f6a
y7U3sLcD6bBbVmXa/D2mVFi6vn1Y54wMwhtI60R7bFMEFvEFIoGSlQRK9+VFIZC6
nVpGLIufvRiwjXkXUPk1bvE69WWrAPUKaIIwuZ5Oly5Ck94w6b2XsLrBKUxg0HFg
VQEJUi7dCwSJb49GCxPIbuxS6yNnEU6LjusS1EUdWB3hYsl1pyjwCWQcgRPy6a6e
kP44vmoDdNlTZGuEpkKeqfTPJnsg7DLWsGKP6rW4MDFepd+xIj9TokNS2YIilxLR
vJyEYRAcKLTGqTPj3PuJyGJmgqxFrxaCZ+rcFIJzsP28n8X6l5i9Di2x/iIxiPvp
IgGqp4B6CjpAVyk6c2NHQgt1GSyjtUpr+yrPVSo2BMaYB9KQmn83FA+U7J1v+Aaf
YR/+RbfhXzDP9ldtfmPC8PGKM7xj8YobnxanQluovybeCDT1+3P+ipe9u7yNG75H
UksH7QdLoh2JZck8gwCpHphGESqdQJVWyRzQS7jG7wmoBFfDeEYuNPOuZbkNct2M
RJkr5m/2y5HGtcsaeSEwa8xF42f7liNs7WYoo9Aqv77yV8ZBUPbRipqlcJStzbi6
XaMlF2AeySwFpLGYhZFVLRI4NPvRSfNVeR/epcNCV9VA80fg63LWvYz32kG3Ezja
r8yk2bzjArL7WWdDQAdIsQuPO6xbrvyR0krig5hRwIHS80zhu9jiMbe81MQRGo19
7WZ0FcVMtWKlLntxV7NYfI0suke06/o23I+NPHcXCx0/8LT7EtY0vJuW+wQmYRs7
SxftrWmqo8BiQQIkM9QKzv9ZxBMK/AbWnAZFmkbqjIOK1/cgnsXlX9NdusHRadfo
lL4MlCZj+igSr4ueiagK0mNqTMtVesmSuc6T7Fj1KE69z0TuNz+kPZ9PKQezLPwM
XDzfYX3cw7qln8XSWHjF7h6STzPj+AAQdQfzbHBS3GskJ4RlQ89Ve14dbZlfuAmy
yxP4k/esgC1+Q99Co1k5H7dv3fhdAeEEx/SeUVJ0iee0M/bl6nc96m2P2j2tPdM+
lVkJPk/Y0ReWmpMLO2tNJJGvTt2tAa92F0WIin5G37w5rEgWl2bhVt6FSza4VXyz
/Jrg9LxRxDjiEjGDqLYOovBpkGNXmDum1/HRICDGH9CgR3GGXfeic1lr8iM1xKlU
STup3/N9CsQtxso3n/58mcRK7J/vyIJRMbqKV1xiHkVAekb0t0dnsgPuxbkw2ton
9xdtRSj6L1xxFlzGLUS+u4M6O1QOYJPV4TyEbkQdPwpmC7Zv5psXC4PlQe1gn/4O
+j4F20A544XEPrYB/XKf6BGD1iOsXPGJra7gz4RKxuE15HvXEKudM0vpTm2tJcbO
Ul16/TZT4KVjarJ0LbmsWG+Zo6+z9/Vs29Y52RwAjZQHR9QWxGT3Fq1C/wHaqe1r
Era82nDOAK3luVVGLxZ6hBcfdWAwHpEeL564+IrqLmGcSbbuoaeHXAe4MEAfsnnF
Ji4a0fM+mbRddRq9ULmJbkIAjCLZcuflyu6lJYAaRiuX0cnqmW88aAtqKbCYV2Qm
dCMnN7qIdxLtqhSiG2yvFKlQ2F4w5q2rNOFpXi8yh4LXpxphiiVl5FRSOj1CNo1A
tm9Z96zWZUAIkNnfXBHS6DV3XpwJMjfptQE+vS3Epen/KzPnSwL6REDeDszmOY1c
fGVq6s5QZ7xriTkjjmgaFxA4EKV2XW6X5JojNfTTM25yb3ex7kls8vIg3C2BDMUK
68E+s3MXZTRTWOz3OzCz/2yL1YwEiSINVWNOz/80p0lPIWgTVwdlXgjdjY7kfofS
fWddXhNjE2AILyZulZWsdsfPJLA2HZAtFZ9pmXGgtt4wUV3LPfI/abwZdo57uifG
tVURQVHO5n0lajxa918/brcP6x55AbVN8mCAcFc5KGE5/1ov6/bAbGniUg4QkZNj
iia3rarO5aHQwqCeqrNjPiucC4Hk0m8nfteIuvf6jbCggVN7NJCpDwGbfatp+Kj2
9QdIq9VhyZ3X2pqZEOh5OTKbXur/clISQZlPuQM1tMrFIQH+OWx41gTTuOcIcv2a
0+yOZ9akhbs36wnvaXKz1LdQYrk+aR330k+hBbkdM+iqMibY8uG/ZnxqjerWztGS
lohfRv8ykEu7Kl38qM4FC8Sqsp5yHTawMLNhH4HCRMCJPGAbMwy/ZP1AH01lAST6
hCtnSHhJ++NAyQxlx6cBs/hjwNdARhxIoxOijdidJuXTJv6n6L/O1zCdC+mIMDgb
ySTtnAV4PHwIYZjcT5+xlGXIVrkIsfO6B3h8rCrNeeiJDSrd7ox0o/OwcE42yCvF
rUPmplnRdMiWO3XUxZ6kigx5b0v5rqDm4jLod+hMJjQOHKG7h51lh5LS2rCFQtGL
c/SzEGlzjfo5c+vErMWSl22rA8eQpBYPmYnSagL4TeV3dYPFVFvMns4kn+jMlMjr
0FZuRjnA50Xq8geUJbjGY738n4xkr6KkgxRI23UKGDDmeY9PMjTRojIDuaw2aPLR
AIrsom9OE9K0ChJ+7C2zqUVULXWGPYoyN95Sa6laMM91Pqee+kTYtQUvf7UDqReI
qtiAnDV3/5lfuj9SvW+yd0qBk95nr4HoxSR8k9DzizgpkNWyPF1NzS/crFbFZzU2
YCTiiVKk45lks4K4wqMidfYdJXsxH81mcCWIuHCnwOg3DwO+jZlmjSjyRKIOEyba
rfp+T20pHX41+46mIQcXcPJEjYVI0JI0I0qhkukF/bbzM4aKJ6b7OyMm6VE8PBJH
Rz0nfr4muOhvReBenhqeE/id+/sXu/qzoGfUTLzuulFdzcNxxC4x4d2z8MtA6dS7
IdrMOcS8Iy4Z1doFHn6cvhI8Hu1rG4G6uFesptJdawpmvSW/pW44yoAPikwn2hoz
EL+XZjCVRIBC5MslgsFRPV+kmJbPlH1r3uMHOTQLymBZzKEqH9KeVb2Mp4KeuTb8
sYkkZECZgJQV9DWXw6KHD/RrKx/enLeMKO6B3M5QESYi4pC8eUhMGaXyH7yb+mcP
ZPh5S7mQLY4ZT6rL1l+gzG6mzT8khRQt40tGWu3r34RyOi1TmSe5pdxK374XATXX
vb+L7gho/y4YaG5nBsdbbNd3guWz3R+lB62cnkLZPmuo1CyQH6eS3Au3DyyQWu9P
Qhk6JVXDh3C5/RIDvviAQdvaUXApLK0/059m0kxdLTIVBDgJJndTwqD2DUcKGy6X
bsYUxp69AZQELrehoiaeanowi961yst0yLcD1Kj03zNROSjvkznF8ligblFuUCjk
QlmvX/a8B4Uo5y93eiuJN47qqVWR08h7R28ybr6lIQZ9zF4rikHVP4q96ZQBZ0FQ
ip0dU+IjUUxbxJ5KTsGtaDJo5bYNg8M+hUOiK062sGaPlruE6S0i42MAZtdM0+F7
/PMDCcHZxgGTiAPYhBlVKFQt6i3hMIB8QMaTe/irzYqIZqIRHq7Y12NO7/GeGeuv
FixXgm3P2IE5RlwPY/9oKtoRHphzqI/wer6NDPYOBjhKttxu2ZrZPAbHveX2sR7b
gruLqe1j2R2buf1NfHNC8OHCOwxSp6izAcSao07x0Z98dm60QBNDr1Y3aWYYJi4R
I0NF/pskbhumpbIIOtRdBsJZgHTcUAL37QTLyRFGdteuVExQCjVH3ouijOJXEeXD
J0DcyKr6qT2Fp5PJUFj8bzAQFUQAVUHEBPNAh5o2r03UAdZFfdS5ma/IsoxF6p0K
eNoa7Ii+vu9F43vhLn5pui0y8zlfjMH2zRJghaeW4kcrPuIHtJRBLEDA5GRIPip0
9ElfW3lQTbkQHC0E9SEUZ2Nu6sSfM0f+0sVgk1nrG5UPttE9hTtvO8hvPeIhQ9Bg
YEK9ZOkaOJmMy36GzkYA2LOG4PLAkYTuCh9O1baz/NcOPBa7VO9dU3VwTTBjrTub
nKyvixUiwRzDL3fhgZT009mCWL6lYxdreF0cyLR25HGXVBFZXonp+CfhSjPFVnx5
C4fGBmIYuixrniBPp7tSfOAfU2pw3UVhIs+5bBJm4ZsNViW4FKslr96MuSoPbK+F
dC3JsseO/S1j00o/BV3tna7j+exjZXZhT5VXDDshCz8Bkdk4uo0FtJmBfrKzl/vd
1dPZepYsxAuFgm0T9abASYNP3cBYaGK4OgWJJ9cC+/NTIcVmnO84qJZoLpVqeIkF
d4KzDtVfyLAxPU7ZnTwhhFpvahtgxBRczoATzWRrbzkvhFqFn+RL0x3blqeF8jbG
YgZzNyJO0VfEIR7vGUaskBXp9aYeZLamG3UBG5rgqf/1DdWDkhnoKhnqjFx4x6kd
U3+fLBGABhz7YOlug6N8UptFPUYlAlQStnDzdpfs+RqWqHFoDmX24DmRnGkIiYZe
wtMRxJPf3wyYHBS/lHvbVBVR+XugW2t7BRYeoYGgCqQoMmvcafPUTqR1jRAMAwS1
q6SRf/DR/UjcwK/sXidcatu8BZSgFoaFOf69sZJMdGy5XSlyOOIt3osA1FUAo8g+
3pvYvN/XNotqwMXZxHUhGqihEE7Nc8KQ8zxcFrpqbI3NSK5arHM8iSj2neVjV5Kq
U7kgLp7e57AJG+Tn4CtrqB5F1wbj3tz5r6dkFCHkrQhihHD627D+04x3GkGSGr1L
5q2RTvniijwS20cmA//afEmCg6DCKYt8HpybLa9BSRQvfAgSqy0UUO0t3ZgKQc2+
sWEQU0luMAQOrjPLS0aI5ziveJKcN19v9Xbp2n7w3e8DiGYDbslh6FqRQpTrnK+o
R+14hwpv1IRZCri+aw931Y8gTRase+ZBaG9olvc92UmZUVipPW4kRLilPIci8ZH+
hBgee+TZIGMob1rAWPPe+Np3IYTF/x6AvLNKJcrTO3ZQ61lhm1V/MQgT++TK/mBe
wHDxixavv/w0i0g0UBf/aDjBuXgIo/g2ahVwWBYKZR4CBNZrrCmOTNBgT45MVHeY
stcZQLvOSIaviq/oi1If2qatO+7pNGsuzpBBUFnrxQ4QzOLR+VuRYDE0sDpVcBNN
tlY5aoXg4Id3qPSDyqrzcfcdSjqCsrbPCGjSPkdmeKzFLUSr27ewkSQ/jatbzyyJ
vXaJAO4ITwzGOItxP5LpqxueoJyOHmqPkXC7OKQa9G0NDitgbZw4PSbDT+bXwKog
H71zsr4mDrnPYzm6lFMQE16Nm/ixAJFLh5HvytDYG2EK+5mx9h9ZlBC8c1/m4Klm
8BdP6htoUaX+TFOaQHHwJ/MoZADT8btFocUP6RGGHYZjJPcbTRFtFOw0EAflYS5+
psDgNfRWwHi3ewDg0vM5KhvrrT5krKJmoZ8nn3eo7Kd7AsJ4s2WDqbXGdLA5cL38
HpN36F+pBkKV3ZHyHQROhMMV9QflEUg9IqQM+aQC4yehIoAY1kpTWRESZaEcfFMW
2mfpw/GXJfOh980wbo80gtkFBZgttAsxKvYMquEoyssqyqen2wPXz0MbOv3aQedL
r153OdxdhHkqBJ2ueFyZFMffEXYiSe7Wduqymvks1TBX3eTJGwWajYznhHIF1Vkd
W1qJ7jlPAS1n/ByITCH+o1uJGIl70LJ/hmAtZRFoNF1IxEDJn4BaU2SOSaD3yoVU
pTvaNweNB4lAAZH5wN0aCNHsO7qwDq5aRn3FPyjERV8RNbDJnK/SURPfCahwfKfA
Ci+9AYU5bRM7nimeqrZjy8KUknScEIweNbfYvLvB7gVNg8T7EAwnKZpf1qH1uf2d
JLBflw1tf/9VCMQ8sasCCWPcIu+XF5JP3raIUGvZUp7mSTSRJJjmEYd0F70toV30
fqwleAmQiajvRg+11zy9NUPQjtDx1J6rQBlNRRPIKladcpZiCZvq5SFGV8Tdl44S
2w94s29xLTuUVbVgkxv28h30LCslZCuGY7PwGqVEXO13JPNTE910dIz/mcm8434a
0NBl2WWUs+Q3CgnVEZDiua3QCpFPmFywlW7IhkY39URI6w6sAFTIzBPIigL/EtVA
x7kkgAzV3HBrHdNvPMNEFerxNu80+UIqMvMknPePEzHadCvUqMqqPs6j+j/SqnvJ
B63WG6DIr8+ETQumQy4rrIbmJC56S8q5d+Ep1LTyCh6okArAG/xiTiNdSXM7SOQZ
3pcH0yh5BRHL35s0I7l2i8SC/sr6DBPq4JFTEs23pqyxv75vgfuVa1eEwsD86/vL
50vmE5pvGBEYenmLYLP01HAs9U7xLGr157GsfLkC5D7Rw9XYto9NCzvOxpkkYnDY
hR3zdUAM3qNLI/3uEFp0wOqGrD6c/x/aWVRB7Gl+L5nfKU1DtD6kkuodSvTyIKCY
w0emvEYMC9U3IoG8XwKj+ZzAd+Dee2/uWPhTrUOn3oNE8S0g/+RphqctT7tJMNhK
Dt/IIRqMQq/DzJSQ1q3H8k0CdiZG5MhzE0p9I3cuG4Q+TOnpTBPEqE96owiFl4mN
GzpVrhyw5WX5kO10e0+nhX/f2ev517m9ZMW5uLnSLYXqvhDCc4I1wvicTzJlV7oY
swg48u6vb8Pz9tpACejF1STQDaxZ4wOIwJCNxc7Ovw6GhE4dzk1QqUOSjveWYnEA
zJZZurOE2pUcskDluac9xZeSDgJhG6w7dlVtWYGwXpek5StAXeGHHQutI92i4D1J
ygIeQ49WyBTfhGHtmEzh+lBEcKe5bavnvv6admSoAIJu7RLMRhxp3sMH2V/P0N0F
vnbexUX+4PpygnmQsIaaPPUpxyyPHkDsGMWD1oqBnJmovjr0Ympx36UNcdi1dUad
q51x4+pVlqjqXbqYa282U+LS2OIfMRClQI2sQMEK/F53jWA9/+8DotOfp0pYRxl5
QazkdxUToWwZr5SLUbOBIXrsLAnUEWSEw7YRnk0QGi24ZPn/Ll8V/ICWiB8poaQN
atDlmvL3LE0SmeJUwnkximkMvNaDuyOo4jOwJprhLbZ1i4miQHjsy6UJmZwnwY9/
XQg/OD1t5YLYnrbKn+lj5PM3uXJh47PdcwxHzNbb8WP9cMeFLWkuKYLtLCyUwdH+
SwDiBicZhDHxsLfUY8NrDUr/A0shBNlPsK4Wbne4cN1GGtoHnOjf6aZ9sAJUTROm
233OBhaVssQZAKaeTOC2L4DE/UICU/nvALB1aFnp96I4uiKlaawXHQhdITNWowJO
E7/7RxqkxbIW5TvkKPfB+kENH3Kgh8cwyTParfF2ntbmuCX4W+iT60+6iWIRK4BS
81a50yWuZXlg0O6ItbJMdtfGLIINNIQz3/9/wC4WvsjNb+f/Idg3hnH05Qji6f22
9XUljATeedVMG/1CGd+OzREPoBpLVMbk9kJBdPM2LxW94jUuSaJ5eCBszO7yMnFm
wzUXCj4oNjtFE+Iq4dSSj8pXUIVo/XBqYBB6z+r2YzOLFqXBMUu0Tdt3x3rw6x8e
+pvAS/5oliVNHYU2Gg9mnBu2MHX9o64n6QHZ2sPwadq8yb/xWHJMbbaYlH4I6x6j
bTO6ijq3WcsS0Nrqwx36Pk8X0kEOhBsyTx0eRHiT15FTx138eP5MIaw2YDqA6oXI
m4lP3L53o9SeZLJ6vIAFf7dzmQiMwlZwATU5E/Id0bEd9Bwa2hmRgEGA+yWI4WLW
BlUp71VoQc1hyghnRwGz5mZ9YX8pCJXK6OZj55c6LvDsvHwcTL0KSxLoUrFAderb
XnfRr5jvAfXh5bUaWpW3xegCxq8cVy3tj/etlClmqmMfn0PlVzhWdQIhWnAKBbgv
BWi4s8fh5xBlYGL5KaxajdwjxjP09C71VB0KCaRRexcXxD+VnbtcQHnWQ+FtXLPl
/Z2vE+t/+tDq2HQppIb5XvD4ZdQvHbebt7xWZkzgp0uSK13tAv8apNvbaD3GlQcY
fG+lK9d/0t7C2dvTT32ZWcI9HjqEe08uZCkc6kMipln3IwwQMdAxSzYVbhIYeTC+
Z5HRsjIugVsW5POu9pWSbf71tKUvqYhNFLJgZ4xfLNzvQZNt96F2Ot/tXOHXC/nc
MFBImU5chnTYpvUEUpcbX9dNFD1sxb5UKahPM/2ZkmVAytF2BZBPcbpBdWZs6QYx
f8xeBaPbig/RT+cmKIewHdcTjRYADBw2OaSZ5lraB/YukXKxCvjrLxG04QjDJu0D
dGh/qAQTSZrVhel5gbxlCHObSiEy7ApmL3RkU2yai73AMMmio0jTQH3Uf3X9KEsf
lZ90Ji8T8t58ktBds9yaliZUmbM4c7eMQ1GptcmqWC7EgJh5UTUMJ7ZvYfgjCaO7
ef0vHdZhLptgw8KvOEVh4QIoLrb5ZrUtG1ncPo4FcAmQzJqR+kC1brVvCvrOf1j8
/dj2/hdqN2nmVXmT7CROEtKPgkJjiUU/Dn9nNboh/fwQsA2Fs0PmO8SH3JIs/8VQ
L0pnG6eub9qCGi4U/b4ayfTcswF3gYxJstdsrQW2c+cUYOCvMOY5y8B8BzrQzWfG
ZAr8ic1pquXj6f/TMIJzlNWXSKxTPd+wYSonVOlF2gxAvLoepn2+Uav07Rj6DEwd
IzYLm6HppDAhx6GFZPTxktO7Z116xm8MzPyZSIGqIarqz75eVtkltlwcqR/Y23FJ
2vAFMmhWfhhxzYuOyOXt2hvTRRZQZ8zPKh3zE0VihZXTibu8eFpKaMX9jCgx4Ph1
TFSLSwmZhqJweA7zPdhUyUCKPAnk9Qelu8pE5ykey63gQMJp+ffg8J8bGHf3yFct
wahyxxgKKckrq+FwtwkT8R60z1IV3iG6oi0rGAhmXZfTH2Gsbx6V3Innf1Db7Wmy
GZyFb1Ke+MJ3l14Xd/+r431ylu+HGMuPRr+Uya1mEdXuj6ukCg9PQr3CBaHygHd1
LZoEX4QYYr5GDQ4tEbPIwR4yDMJ1mOHMHZu2FWfYPOgiVK3LMc20gLKBb+b3t3py
1nbWPQDnxak7DlX9W18t8GQoKCbibPmn8Jvh8R93Q+C5ht4ug5PxpArEqkyqg8Jp
V0iB8XkjeZ1RGT7BeyCqmAIi+8Zb7T20vnuAG/xrFspXtVkgW7mTohwlJYTp10ty
+4fU8CKxqmAIoUsJV5kdcmOWeUGc/qfJcxxnmKIUVt+OzeS6mYEzJSiDH2F///aj
lPo0wmG6fP7I0LmRyxQL03/8yfoWkSay7f6fCIkMiLeNoqa62LMg/BeM9sD7SsvS
b4Y/H2EBWR5DqN1SsJ27XiumlXisPt4XbrYiaBSe7WYpZ6LChoSPmifLImBPIG7A
iJ8LeWCrpNPpGuBOE8VCW8fsw2YmtZJ71V7UL0Q2yDBGABsSITYZavZcSprzPvu0
IRrUKEQRnY/s6FML0H7WiwJm4FqO5h8h3NZpjPvMZRpVfN8fAcc843os2uEumQIW
lFIWmZx2zPZRs42V1DmrGVvEiQI3GWJH+lLN/lIl6W0x/iPE8GIMnu3ljcrmGpey
ozdEJTA6I3YHU8Xq0/XU06HdOhj8xQeXWRynu8PRaF1CnrElMJLAH7ih4korbfyR
eTUiWhF7r9XH0Qh/1i/71uZzFMdzsUGVl4AP5csu+oDr3HC9Be23kLpcAQz6i0Cn
65idGi1cQ5wMQ32qHlh4/1DeFspXO2Knd71CZl3GlF9jyoKMtPvlyRHbvnvPS5kB
dllz6K6Ws/CzsMJi+NX7SIyhaCY+oKxRtUnhNLJa4uJ8FH9BABjmsyoz7amARcIT
uXVynmRlQL464CwiT4M9aNHUtu1KWJDbuLph6A/lDQ7ZTxF2nyFSmruEzGHEypSJ
2Wip6aMJM+rSdg0GmQTX3gUjQ4IfgbWiq2eeJ7adm8iHq99GsyEp8lnepvbRA3Lw
9/nizoe48uFLLP0DY1A9X8SHd9pxiOJqr5QmV+HnErbRNC4YDqRkTtmBR2R6clSX
DS9fohjqzQ7s5ThGQRioMKTa3IEtcJE3PjL4o3KFzrvNm+ya97Lgo6c2CNiOvmL9
63NjIvKl9DdbOgBt1EgnmkAc5h/XDC8xVrtdVLAuOjuPOvqnBh0/j3+favWYZObQ
6lqYW4zveE6eN99+RHiIYEJNV8cdoMEsSen8yv+WgBo0g8vTVHPWMy/S0q25D8mS
c6R9OR31lQt8u8qZwb5VH4IGiUEvoPWJFDK1Hluy87JOLSsDfdgLvzJZcEo5vfuS
V73Oq5dXz1NhpT1LHEHt9IFM7MXLS55yKcGz7IrZxAOJJ8DZYZgmbcr+FKot8kkH
/cQLjyqUmL1Dm03zAnsKpETan5t3Sdfe4bfpWEf8ajJy46yII4HCReiqE7l9gBs0
RAy4gsu3zmphQL5TpD7XVw1ReL4PEs+of4TFxD+D1DiIFmSizolkHjqn/dt5YKhg
wTYlk+3d+hFalaehKh4jidCwgkA0+0ITSu3mT84g5mLALapL84xxNH+k3RHAKnfO
GqYNV2c8+hZkBShoenXntDp2YHckdopNrKpyXjZLpL6g7+n7kRjpSA7fjR4E9TfL
Ne118smsUBe5fNklT3zYUX6qIAYJiy/BZnllEaXTafNldB9MqVm9WoCGtaesP7BK
+BUoBgzgtDK170pEBoH+lEVKGOKlSYIr6vdEe4oocxCbNVHKtVhmnukQPA/kLbOw
9iBzJ8P+OrDZS/hK/VvYM0SEe1P0SruybubdCxnoptDFQsdQC0uOPb+wJ6aGBmvE
4VUhmF12Imd4BFixtA4T22YL8ioON9CUx9SUg7EHa42vR1ToAad7i2jFOjp4RwL5
FAAvzcgsLj3hFEqp08qYZQKBKJrFF47+rIekD8ROsW/tH9vZM3V9B0IkiXv+X5mh
joD7GG76HfweOcVUhCep97MmVoUfn5AsAniAprNJkCPf9eEXgqGwbXEOtBmxvy8q
6lb1SUvSt1lsw2cftf4v8Tb9B7KhfID57Lvq5QsanifTXgFakmQUWvL/Kges6yXV
zb9jWstGKh9BYsICTFeEtPPTa338rVow1V02n/xDmi+F66KcjPS5wNTEBoMv3kdr
fBcDSVDO+Xhm1aH/MSfi2OP52i6k6/QuQspOJuQ8d3otqvJg3qtYcjkQHS28zDJl
KEcyhcKIZPMkiFw/QuqWjTXwKMUkd81p1nHAc3ZBZEV1JjYfsWU23sShfX3PTHZ1
nrRDqxcGj/ZkdID0+UrcZGXUQzBAV3Pbdf+CZnE/+1qctjJ2t8rFymqfpEs4y+lI
gtJmIPVdbyOJsSKRec/6wjOf69ptghWomQBjN/TZacmwtVOpD2nm/SLPQ97uZes+
ZIwO/K2+YJr+KsqQdiUQFEwTf8lh3HHWaaQFGBqcybP6DNQBYpT7qTJUdrNnCoTf
CRDRAGVQvp9rqlLGX8GpB1MpgorlkBfTwUPO7xfrrR4YLqRZaTFPnAxS1my6N/+B
XtAblL4UqdWbzg35nXwbZctsodxLyHIwqf7JXlUrKmLV2Ik5XAnivAODdWbhp6XY
8LBFHDew4UesRl2UtOWLfzi4RYIh5Td0fqeq8P3yHPIib/UpasUn6ufq7WVCeNLI
MdkHID3nSis0uejweAC6NPYtqUqRADk28Hug5p3Bc7641e38i4rH5kVDaj/0iShs
U+Y2saa+Ca5D5SbfxuTFrlpKDSOYcmU5QO9Tci5rBd4kQ4CpZ/2s4TCceqY3/qSv
xd8GLyPpI3sodD6wcLR83nqqRtzm0u+mA+i0CSlGh1W9092l7bfpiNLKK3T1gkG4
Xu5bsXQkZLSu8r7QkTVWHPC5nk1FAEWnkx+q9GQzLQqFStkmIX1BnoHIaruCxQ+a
IdsTQ/ayGTQ5FnoouLYxh3IZoIJxDPwIAXh7fpguiPt3dWcJCh57NDgS6SoKg/XZ
gX7RxcV60btL2RB5Sq6Wr1z8GzuQ2Sl2nGOXFMYoe2XrPBa0zn8qjK1ZAFG3FRie
vEci9axNmk2T+w5JTCg7noOQvHAFYfQVwK+GeHn7cYgZGFt5BRll9ljf+WTMP8e6
CPAYwo9QcsEQZoOmDvpdTsz6b0auBvMsWAU8fpAtCmNRilCcVfLtfFPdd6Yod/hD
N5+nCzXUJVUW+RK53dRzIy+xEXT1U5GmogtTDieajteH15cEkbsNSrf92SZSfufo
kOO5Bb67g28aHqJODD/w0Q9SmNAZS6S8f1Hti3pI5YLIoLrUa8+G2XWePzVx0S86
53Fu384jv26IOdOJRvIyyY60gM7F44HoVwzDOf7Ce/U5ZB4gdWcZ4zrX/Q3dDveO
ZQFUOAU+dxnVs6fUfEGh9/+3VlCo7FqmDb22cZ+MIYc9XCYgRVR1Cuwcp6EBpPIL
Ld5KvkYtBl4M6Ex6IEAbt10cG53m9RaW2x0cwVoYl0AtlfH696UPIPNZy70kCTOX
zeplB7a/KFmbWXkTPmVxSz2qF/5iefhH2JNP/EHAcr38/j+CP+LqLxPmt1ov6Ugm
v6i58pUTlh52GHHWUP6nbgpF44fBpil3UIA5MjX/dm0jKYh8XWSu+Sutsbwds0fW
1FpVPPlw8CtfR+lGJgfa4UV+ArptfEDuTXYYz5KwR23U9nla+aU5FjbHvHdtJl73
KbZjizj1FXVWk4B7a0EypipKjZymig75tXQIX89RAaEUnwGEcKJtTcKaDU+wSc++
jH6hvIz/inOCpI39PbN5YzGnS2x+WYVLkWGPZTo4sYIyOJ3tMIaFQDMe7UHhj932
l2d7g73jI76A6FDI52pxIvmoINuySEd4Czi6gvUUhYy1j8//59ZNuf2BodOIrYnh
6a1SNpu6A/Kr3vcJidTyucl4l7UfgKkClJ6yUWQTWkqjyWvEaO9jMZqtuaPFwlSZ
Z5FGWkeFmmjzGZvzdypnoTb9Y5JLtMDlbpgE08nYBB+iKTgW+pK+vG3VW5rgyg5j
fWerkr+QxTqhhby/JC3jBUMNfV0cQdmaBEx8X1K/w6uiGVbmEZ7xOfo0FsLOApB2
wOjEEtVr85N60r/faAJklVQNjAJy5UVhj2O/sQiMkTuvfKCaPjbBMyQb2HMyqkEn
+h7PvWMQlbTAnMlRbPBimyeZb9R5Ktjj9INpQ/rzSwze6CT2EZqaFT2DPE+LI6l1
daZM6xIg1qipyMzJSYHCRggi7UkO+HTLXnsO+8p/mxb7h4Fogq291JPBiEiee7aj
1eAjbwEYgvwARU+FdLViwQlBXFlkOaheFL7Ts3dRkGUcPWS3a3aRXLFfsyLlWASz
Kinz3tw5TQqVbL5+z2wfWo1Zu3DHPaq01dBVr/aoiV8mVFdLkT7MwMQU0UqUktBa
ASXhJE1Ogsxze67UQbZ42Bwq3zU2lR9Fo87A6h91VSys5rPcSilZSrByxZ5J1wP6
miqd1/PVsYP3LatoY3HaBm8oCBUmFzhaoBbAULb8Rk44sjeWSeyN1CWpnTKyk4AU
qLOwAjaaGuqTFkPOOHzVwDPAVstJWkwSDjXGQas0/Ee1BI/zCoKlpzekIyC0acUF
sx+nRGqcqWSR1n9T0QRhKGBqSqUhDSLSFilLgbme8vV1gtV9A+5bWeL+/R4u4Y6m
HEUTNT6b3vNEiq/Ib5D5Yfg36odXNwVWMfp0FVxoUety1joHpFVtJ2UGfLbyI9UC
NbWt1rZEyzGM2wQt6b1JW/pdG63P8lmU66Wg6e5BZvxo6Hee1I7A/YujzmTs448L
VNraJl4lhD8XAnDO/4+/emr03HiMvZ3Vp/fIohmbise0FgM2XSNKJj4toC2jL6O1
dtjO9ZFC5DE7c+WVEPF7/Bz2qXANxaQlRjfBtjHpqE1EX+/ucsTx692bb2pYnRgB
eQn37G+NV/x+13J+3USnrOsBrOBchSNIW+r3aMdqzp1PwRcobnoZNFBmr5YKqHH3
uWpB6mbWZhkBswZ29L9SCcYVQc4LBRnJnYTbrwIQ3gdJIIG0xdcnXc5CajT0uYZK
H9HZ+2uJr6jL3BjoocN8MmwgcsKF6dtQdjPqNmTbk/lmzNq7wpq/g3p0eYSgJRNi
JTU3jX++xCep6gMzPK4c4LUo84Xux0JrDPAzueqtVhrdixZ08ud2/zDHYOhoSW9C
UAL1as4wkq0ikBdkQxf2FnSHhttQRJ38Y+yq4XnpWtkPQJTrpwLHqnyLt5/jVLFN
bsOzB5IPnriL3MVymCTRcaxXp0s55s8vDiVseBCL9j6RNTkMi1J/QQ2mTfD9Qnni
/bt0c5T5aPutLdYTUE5JY1aFjOLCzMUf7wr93kGleQyDggqdMi6AHmhbpe9G47ah
T58BWZ/0cCJvTD+d17nSsVv/MD7tg+beJfaCqxTcyNfvvO2+2DLQh42gCU00IybZ
0GOTcS6jOHUBth3Phv+5cxWuYEioMH2nfobQ5tzZICzh/o5WxqZcsvkobmvFMI6M
MsjR3+KiVqFAhAnJxEa5VygvJeQQ+l5Ar5w2YPXufwuA4bJXbStflIpFQvRcRNQX
uzxkecqCWsQMyYyfjvf6MSZHyoKyrXMs5F6+EcQ0XZUhH4M+TtHj9Xgjvkltb7o4
rJGrP2EsAwq8feBcfAWVkZMIy6Rvo4tLcVOn0WVmp6E6rwTclC4AY/gYKqjgYOEb
/k8/to2DfPSyYbvW2ggaaVqj/QbMkTnQaD2bxcqjDPrE04zkhMyFbmZJmL7/wNR8
NqQVdDdNryfV5sSpk7MU+7hiXDKiGtdytyTdHTPAa76xnLQ8RwMMEl18Wk2y8dg8
FmFbhTnzVd2hXGYJaMUWtAmP2JJUKiMe8xGsdMTkU4vC6a30rE+eDjZEklLDbe3W
izMsgQG8LQxWJkrq6zHNVfQoVQdynyPnH780bkIcuiBKURuu9oopO5lsVHvJYV9A
gG3tREGo+WpFNE1o0wGhHt9Cw72/FPDMyISiMlf4egdC9YHYckS+tjSOWOaG+uUj
2X9qFoS9VWxpfE7JrKg4U4l3V/QLU/gg+RVU2/21+xIwUBARrUS+u28v4tF3S+2f
ckiQFjUzEYPHnxYjKchdOE2Eol6N5KUTQL9yOhsHd2rA7vVG+reJ/pQYXvPj208l
WCc+LHIYWNvL8y6D0OOKiPztHZ1Lps5sPheNxPLWEDzfCzaddqcbMljjxZEv1XHj
IBRMRr98U5hAigp9S4oQF4KmO5/zAN8nfWFmFnyWh8sYeTMnlo0Nvz/nVbF8FtXy
JTp8GI6YfsN/KPW+4OV9R+s1PmYSPt5+GcHNUjdkK0n6phpCVKAi53BQqOQMVKJp
TCA0exuUuGklA2YcRY8NpAKFlf+Lu2KMgtABCtMrVGs3drvgyqxJhgpdM3yUJhbv
pVNlMpFigrI3A7BKjMUo7+aGYeGZ55CyewxjkcKGdFaJqv8CuSiBgNixxoIYyFH+
xB/eFZ2KTIzbdavURbA9CIs2aUZPVAAtnVd9v/iXAA3OGBBBivHMnji0ImY+ONr/
U6H82EKgbQjfkihv7qx4JImdXdvKC4dhH5l3ZxstzayUTBhdSOSvwyXPaOTXCfoY
QbRTSybXFcrdyNeP5/BnWH+3zq6gQhxxBHFhIWgktpPABwBhB8PjdbQ7GgRA7yF2
xQmha/WQloCHyEfYwv/Ch29BFqTB6R1f/+esMRBIPSPK9wSsuNIJadvwagbk7Ca6
+kXXETFj9YGlli5cZamPho3PrKrHPXqFOg59sTxohacAuDLByARlaYj2ntkQBwEo
+ankhcUp2kjHnRitnSw36KQnt4MB5VHDt15N2HU2HJ9g9Do2Ri43ks7gRC8DT92E
UzH+MY21c7XRAwoe2kQj3BUA9wmcdq3rfWOtBm8Yh4qQzsCfzwGa6ea1+v9gbrUf
7bdy9cd7B1HJg4aAK8HfO5dQFDw6DMik7zgWz+gbHlrTnmV8z9hCfZ3qNPXhU6ut
1SCpnRw/hpfyt7DtxRdDQv2HkgQnyow/QYlYqOhrnOyAwkX57u1FQpdUq7U1s5ks
+4ThoyyjGgitYMEaP7bp3jWR4fIOyAJJdjpDdcfYPXsxUbhoRSutnh/GKB8ryMh/
Jv+GZafDpWhp5Ps3HDQtgB7hSI7tqqysuMrGUykCGUG1KIqDeR8SKWgjcMvodYUA
aZ4LIU1CoUEGtEP3BUdVQxQK4JoyENVOf+jAhaOG2C/r977dNd7mWLJ/21MzIM6o
p9usAraB3ewdpSB7HRExnKO5OXb3rK1O0rq3xrUt0FTNbLlyoW8jKKnlzk04dEO3
QFFKqIjnVsBvVpKVG+/pp3vyyw4/7xsR7EsHN0Vx8UTH/5K3VMa77cdxuscJiGr3
vLNGS4l5tH4I1ZgVVDk0vFTtWTyGcLRdXziKjF4rT+29hBBSdkAwpbVNA6c1JVtD
ZnT2LJJ8+x0HOvccFiWjINHGpWVWnQRTOrvi2HZ6HQIKaWS2FpA9bhcx5C6pqlM2
c/Q7thzClO3C0DKjiN+WzURVRG1ACQ3VTmdnCuKVAdmzfTGoxKqknS3GZ4RBV5Tx
nHLwgjKuXZz8O6poGGXzKSTxPtvy4bToK7ZJHz412FmaxosmOBHzTIOSeR/RBvT2
mxVwmoBy6yJTUgn6PXskGH0QCMEl0r6HIINnklv6Jdh4a8FTA+m38OwRC6BAU5ai
Y/AQ/5R1BCm7w/Fsys1RijPgIxoWLbnBym6LNcNzohSQB90ASjcJmADYkTye8b86
2C3HQG4A4m+7j4ZHPoAtG7fpV4CYsbR04rzMQ9kcm1qGEMuC0O14Gbmbm8k5XoaZ
oc7kxQtMVUYkVoH7IWWOo3kIzz4euro5vgqNWjcxfbOeOs69Pe/rqYb6ijOhbCZJ
Jq1vvtXKWyViAPTy4GoMoy8dRoOgtDGqj+I1fu8z22OJlDJPH+n36LlM8LFzfPI1
yt8DWyFnaB0qbItvqX9Zwes4wg3X7qMe6scXG3o5XwDYSeA0Qc+YYFtXsSmqf9Q8
qg/gZJdUVeTn2XNJw8lTY6iOXlN4A0X9YR0L/rv3zAXs1ixnE4D3gw1F2WOrIp73
C4d2fZG4q+zhpeWAppykawejcSZT20UjcBjUBEQed6bsW8h6bndv3UC//AofIc+w
XhmDDfLJ/a7GwZZiKxpCEFrfeySLGrkqno6QR6+hrPHQI9FSqEMvnXWrC2InN70+
dx7/V9AQlbg27UW98TGMU1Co8Q0un7O0Em9s4ZRafWoZb03CNsz0uZa6xoXH7Zsq
O8a+6taphg8ozLz+zQubDSOUJG6Hikxo5ANK5G8jznBcAheVzRTVriVq0w8tt8L5
amcyTkcvdsDsKCRlcU8jdY+BzkQ+WwjarfOsA7xkwqfS/lmR+vGBNcbqx5FK5l00
yySJlt5TqUTnz53hFBEp9mIpTKUNbAKf+xdhrbRHtPeJ88os76CXAXwpBW6fkl3x
+jU/9CInSBoCqmKJPlVZ+O6iS+6x92PBgMMP2EF7qP7BjBoZRLrUP9yjBpkbgl5X
IDmvuReuayYl91CaKssvHurNkCfdgdVTDsEdB/NOquaVKk/22eaFBw02In5yVhAr
rH9LpVKULCMgl3yjRYlgbrVPaaU1LGh1aadoPVf5wCihdfLx4iNex+SzUC8DHGmr
rvFxBxEBdQRZuJS2pTxNg8XDBsfSB1OF061OaGrSwHYcsEuZAthwOacX+j5azEJK
0OygQqNO/R/YNeeefTP0v6K9dbYYLr7aG+lLbTjKOPXc3beT7kYd0+qL9eXAbhdj
uTbVYDbBcDKip06YhF17WnaQsKimquwk66uoDBFNa9th41ecJAVDAXFjEQDvI7YO
JpZDw+r29pDym/r5iqBHmmvf+2XzI1jApY+8tAlS7tXuw1o9IpK4z0KvA47iEURH
1aS8YkLOhrFvNTtA44NEas7hcB9FDU4+k12zX46JPslXRz1LmQpUqGIwXNRkehPT
eZoYppQsJnr5jxLfdMmfB110npWWw5gWaCyRGUJbDj5fX2WC8/qPLT+3ugRmjbys
uyPy1zvjLspnENfT88Ttppy0/AlltdU0ORWNnFO37PseBF3xbZddbHhQm72Ibx+g
Q035b5ApNaVhROweF+1oh0jnVC4sXEx5oeGzDPefc2dNKl/dQuftRfElTNJVrD4g
oVXXSZWXuLUQHRtx/Uhtr/7ZEzAQqJl3p/FiuNlZ03lUuY9NxNVO7grtByN9cslQ
2ydUnTggEXguJ+5BdKa5gaJY7uRXCTM1JeyfEbV3ZhCW0Q9ieLdLHfh4OjDvcldJ
LqETUcuVwgW70w+1ppL9QidhDF70mKy2XTxiV8kYyEmC14mygzmNhShfljDJwZFf
B3fL+A17/2QshzVhvlxOvIcM8lknK77L0TNnPrc0WyenklL2pVjgT0H28fLiGaZv
6kkSNFyKOyUhJscV0JWUfSvHPvVf6DFcsXNZZclXKM/kU3DEac2DeMkgjhnjc6yn
ohEIXkCEQuxd1uGxVC/D4fjtvMhVBqwNlBe1ZOIAMq/DpMjztd0anuAFPM4qU/Qy
8DM5+sYe0U+iL66lkWyViAvKiUK7r2gyfETBaosSLoNRgMFoxBRsQc0qBn9i5Ob0
CC5xCxIgNFm2YDc27XjVx+QEucVXN1On0bN4AnGpWiW9t8vccGxiGxK5854AdqI5
NhrkFixwjKThfEhpDu9baU8MyKm2dlhKSWMazJkvpPR2nspsRcq5hcxngNi+WTd4
YHfk7Iio84JuWOKmkNUXR4qJ8was+k2swkLHcPp0tmr+UrsVhzGHJQnxXtE2LWqh
zOet4G7Kv0IBQhl1fCHzFEBAL8rTvTKUk+LIzkI08Yv82r10vsTTY69pR5cps44u
OlM5DQpwH4+ipIpSAMYz4UTd5HfZoHwEnXrQPIsuyRAcWviISvIRMC4BthPMfxNi
GicO5dWRLYgmc2CMFE/tadC0lZG5GZK2Zqv/7arqn5PKaCBJUOMWpfA3OEjoWlCW
6/MYwdbS5iyqYeeHq9YBVP9cKKUVPZnhwXk3Z2uDa/mu3STBKS3Bj0ax7GbMK3vw
GfI8/KwUGusHazXbb/aSuW2RlHsDo+scaETgKs3xCDwiYbNv+7sL35r09RTV9kgs
yYeAPl2MVLs/SZxmkZS0dpZtDCjtcBFlPI/pm6e23hprkb+iRGbEntHEfZowmGSX
f00YZOMVOy83i+MkE3RhycZvNYwg3EjWr0FDrculohPKk/7HeDDVckIwgmWSyzqI
UTqNifKLSUKKxWgQir/WdnvLM4j56O3aESLeFMYPwSEYHe4aljtvcjCUucvbSBJx
GakZWUQpFY9IA1Bjt5ecC6Ns8FLGNAbEE9TdK4ZjyoOlULBCDnCWkoI1n+YeM+Xt
S8ziBp+J5d5WS4qml9RrCYr8dxp6KdzFfjh0ohlt7xMn5UteX+wT8XuSNgn4Ecx4
5WHyYGH9LTeOmsui3CsZoApCFQYUNUGMKpTITb1yuM3yP85GQpMwC0tWWMMJ3QMT
Iyn1s0i7KW1wlsXplNJwLtAQc4dmk9HjdjuWY2WQh/OLW1XzPaDawDwbsIbFaVe+
c2YkWr+mVTcwwxBGrQLAWE1W1PN570PHSyyL8rZh3BDeod36dhUD5gaQayb6BWK/
4j1Nsp7WceTSQ7XMPvWoG7hqHBIST8Y4ALeqhEWhsSmv1IjijLkubL+LmbloW5/t
EW20U0nzHEDR5J48qrPRlrwF1MRlzNNk26QsI6cSfyMJ0ZhcZtxcv8CKYFrNh4q3
l7YQTDPesn8cAezdZKthAk0IiggScd76JzWvw92j3EBwOA1uxI7g4y0q9uM2czdk
zohENd2Abfh7XqsSpys8rH4gSxmTLs7GXORC2xmTp62x/2rKvuVOkw/EwQqAOJ+7
ciyqkV6cqDGaz8wTUgBe/MRPdl0pv+7wtzGCs331qS0skFEaMwhAcGISI1nHBKy8
7H3apLG/XsajyIeiYcwLUE6VW9dAVmP0UCAJgqoczEWsRHJgaBVlppKQePnVBvCO
jFUVZ9elWm0Tz/0sEUOlaklANprL5FA6eWQgjgn8lBYfJJgskES2978pi/C+IykS
1VpRZ05BYDY5Ckx5tvDQ2mSgTVr7j8AqsnNQChPB8MwWel5rMXh/TG4UdXrbr0sJ
a7aBI/3i7XSsrMjXC/v6VLeDk3hF02QBjgvNPQ93LWWjb/yeUOGdlPkUACrJrr4T
+ScrdzPeLcPaiBrC9FOzPBPwMYfQZim3XyJWcR3UidpJD8kidQQDpCRJLX7Wp+/m
Oxhga92L+LxgsS6JTOWuMk32mQ08saY6Mw6lNEafHjjTzQCJycuswIvW3tgYdIH+
gXyskJLlSbfLit5nyaBDc2uDvGtJomCOWT3p1V7TRc1R6gU3LY5N62oiTbxnkuZl
OgEB4U2Y5I21pD9dgXNzfO9LyRYlbrlJqT/hKz2CaeDk2hTwLGVD4/8Isksoy+0Y
+klVJL6KlqrjEQ2631URsNDITr73abksDE0RmdRaXMoArAyhym2QGCD3OwqjonIu
llNejAFingW13kDlPf8QPkZMwD4XEtjwztQwQx8sDwbKqnYUq2V+3mDphYY1R84+
UNeQNeawbjQk7Yo4CVjjYu1wobErkdS5ID5f0hlzMlD+b0y8wMPRWQLp7T80TrD5
p/zuzEUrzdVNMLfq1XSs3c2g13qxgX+YJAdhtYvCXO8V7vGGAOaHwdRREywd4JAw
8RQ+rrH73lXsM5KDd7/XOaYyZkiwVNe/rPAaXqgHL3gwmMVSRKlHaiaa8O5M0hWC
7Nj6ggX7ldfGr29aasVTXktk+KA8dBYcWiwjMvSbVimmQEyhKkQCz54JK/p3R3ut
D40KB0BS4B96Gy6m4DBwugtirHD8wNER3lS+ZULAH9UbSiCODB8ps2oswJ9sJAX6
vZwqjnmULgpU9BLAWGQlW4Q19WpaPqMhSoa4MW6FGFFoqoZ4Q9QBrnChFM/azZpg
76DxtuEJ0zJ0iOch5V858FC4jBtra8QRX+lTLcvbLdH9EHGRF9qjodYZOLEpcgZq
DKkq6e1f2Zhxw/XR8p2kyo0P7KEprHlVTWWZ1PZUR5NC0c7OtETAsPF51bpGnC66
GEvp3fbuYqovKUwGkeF7ayV81Qy6OkQk2cB0dgzpPzZCi35JHz/fJ/UkZXBHJLfu
Tx0GGDoQPLevQgfhZ6G6+WjyvEQEDvK+Fo684fm4IauH0GFuxrFauU2w/ZbxxNu8
s4dH034b9yqIoy/23srCNG3iH3Tjfpradq07pbV1qanM/cXlZYciycDyThUs0UEm
zGi2OILqlBEPaMwXJDeHZZrSNglnOOdXhMDuLHuAQr/ZO8miD2todjTudmgWsqq+
NdnB+ZjEH9hUdJkeNb3yVrAr0thd/2zoU8I9AlSD4ZrxNrgaekp5UoDNehcrIoaE
6z/wbLdgf19BMN+pPrjj4J9m7zAh3Pd55+Z8w5wuPGPotP0fE4MFuODlXz6o6H89
mdMavA7byl68UIg0dIfrCZ94LJmp+g40AdhpyokzlxcxMw2U24xGzuNpvoZPlatZ
36TTm4M7ZS9uQzo8W0xwQHUJKdggl/eCHUpU5VYO/3b9TfoHoqkZFHikSOxB61Dr
+x6o0WE7m8YA2Sb6G0a0lHZpSS1NMRXpsH6BNjJtHbI/+C1P2qp/uP8Ylief2ZV9
ymAvvsyszdsuAeNN7bToWzJY8H6EeNeGMm/ggCdhdOCfqpMr7olvFFL1eCDe/FmK
16dM9nsKsq3VFS7Ppqwp9w+dHivPL77lhqxEIQiBuSNWyw1q7lUNY3dCG8IIVQdB
t2z5slVXxX2uziJncrohCvgifKpAhlsncHIQIxPL/53+vnVLMI6wQF1zbLWpB1cE
vS92ocy5kQFrfRYF7ab0gMmqUI4tSm2i0ZL9XDDr85gQbsSnVUo29a7VNIVsqM6x
07tkhADwNQfAUfbtHJK8FQzxAM6oxdZpXFWm9T3+9fEE14zLyAD1LtLwEUqrmucn
14c5vmWsgWo+g8KaKGPQLXKrYC5KDFqBJqiMZXOk1LjYflqRu669q3ycyjv6utPY
qF9BqM+oLqdfuYNSH8nmij+Df+mZGT7gdmAKSa6WBa0PslzQ0d6AUWxzyN5pS9ou
KS/Ql9W9eI0HOcvJBgEJd3YBSmAAVoeDFfWgOzGHg7T8Jlkrfv6sUAWwvBqWWtqp
AAJeIyrvZKQYSoA+Ycjbr33aiD9wC/YVzFralxDJYjR5yA8ylgFhX4GvRQthkjEk
0aql8ukf49BiVsN/pVavsMeDXD/OZnPtANwZRk2+w0XA/XBHiZWaZBemCI9FbZ97
hK3wlQ75LIKtFkH1bg8jkfb96OAG7PJBtDenG0gcXmQKor/eETd5dWbcZbx92mwz
OfgDq4QCKHoUn7WAB1FMI8R4pnkCUQDQq4detGgheMkJU7U3fI4n4EG9xBufSkZi
3WvNlG16dvP95fWKwrKepjAxyeJAATYh65h06S3r48X9crWfS9ngunC+74dBQllZ
J0M1SDgAtQf9tBXCO7FOvT31cfYsRQORjTu7abDjYb1Y0Nv7pNA7VLz6PNvr8ktD
0KSlcAVh3RuTPtiClHKep87D1++Ti596DL7HxkoOgCEf2C6QTiw/zywpYjxrialD
/ySuLvFfUhGLcLgvb9iLGdr+BYubHaqZWV6JICPHPzLpMVVWEC/zfTWz3co2i+jd
3rph68n9QzDKJmAfu2GNxtQn8wLxVC7PYUL8/FULnWkX+MsJhIMX4+wYRsxVkEFu
PQiE/3pqblQlmd+79a6ZC+n/72hdtjGt0w4zJB9bowlksWZMtIgnYQ1VGinoIC4D
GSJcGijIrUb/O87xjcthnqMbyDovURTLucu4mUr2WTTX9OZh2DMuNRFRWTyzYTwt
BsVGDvMP54U1fmj4WQ1YjOlDXzQ35XTTM2l4wdao3jntT+w27PYHldrXJ+Du0z3F
fXWkzZETypmP2zjqDgBd55UnvtAWDmewUYZ4jKXol7T99bAOpmHxJP5oDedMNuAx
/6pq9LVAR8a1/dK6cZzrJ+V//IqJq/cNHqLwSIvNtWFlKxHFKE7WKNUZ3YtStalK
cydY/wmSmwLCVMsecq9Ybi8TGLFapQJbsoijAAy5dlX/6WL1d91WnfMxcswBmr1z
MpFpWaQKDr/0cBiDh7qfrBaGgA/GnPXLY2XS9GfR9cxfWDYymEdWD1VZjFu230TH
E6zn95q2W8OlErzuSK9Zw6MVoqnPXApIU1z99HXhNctveztuqeRxciBOJLVAqP+l
IjV2i0YjM/Ev4b3/MKp68LlkKagqvOmlt2msLIIhTLTq0TWXCGmg7aIz5UHpnpBg
Y47GWAw9mnMxX0EWe2Ue8K9UgCM9LNlLQDEHCqx85TwcylZU7dzLysoKoHHGaUwv
I+jJP6DnAdk1ETq86rTkrchBawC5r6JlFatyC//hd4J68Z/BMmNk8V5MEModaPNe
GjJDHfbFLCFY0tL3fpT5ecTQnXQnEMTJQ4o3oy3nhongUqYDnvRiMzEC43YTR+t+
oO6eOZcXWFedaaDyZArD9I2PZpmEQULAdDdKqvDYrZgcM1YD3LGF39n+u2RXu3g9
2/e8yqEPT2zjlAkiFFz2LXSZVoZtahZCbPBMmMIGow//OhMYpJTZjZT0H5L8U8bu
raxeq65TqzKZABbcxLIuGToZpixaYjmX9olafFl+hNJLJYkWGsMwpnjpW/d4cjhz
0jJay4iJxaNgtMqD+RIOZpyo6Df9VDUW6BFzvqS2zClA+HlCMfAihrthcXBg3TVT
IwOgg93CejaYJyLebeH9bfV9ulBE1siP7rt6UexW7bxSsKrgGDjTz6Eh6QWZihtS
FCAAKCYU9sqphJwGQfyKglqV16Q01aRAyKMh7NWYLxo4BvvoLcgtE3e0nR5uW24J
fV+Gg6unjYWTipLFUmzY5KXbjVzGk9l2zAnIO7L6fi5jzAyoaipO8e0yCEJEVD3h
WarX/Jp9LrQpmJGl3hM4k7tkEoatOuSYze9LSvrLtplhNG/BNJ1LBJ6/s9UXBFYh
dVWqTEM+Lw8QkO7PDlY1hmJvoXEs+Ow0JR9q5sCesy1OAcYQdbwhmQTHDnYa5c2a
6+BHzak6BwG7xShGaIukSpFhHkEzJXvwK5xgl2x0UF1wTzM8FNAhhYFxfosI9JIS
Wg5k/EhXsE2vqL/d9QXJBx7Uqhf3l4KmMHpPbpwKeJivnHv0eyGi2LYDTRbcu4Bx
+MXiJfGShETZH3Atze308hfFyzfr5rqsVJru0LqQEV0EKnsukBjwzkfWJuGGkrkU
t2bOPtVhHeyoIOvVs+NGbcpXQIlkJ/r6hTNumYgV3hjBlN8L9o2Yk2keEryIgVT+
qFhy/ipNfPmWpAiNEZcYGCcb4G6ClmooG7wa6UHzWzVDvrXsrWbktkPFBbne+vRK
HmKer0HYuFdYtTObVbUOAYTvelNjPQN66BG1Q5dey+3nuySgyMGU5d/l2fNs2O73
qQzskwlberpEBZmFPOd2aU9iG+k8NaosErkOHqzb3IxDHc8CtT9oa3UZzBZbHR7R
nSJFlZYJ9Eqao+K0MUVYrQUUHqqaTA3x/28zMhiKlXcNzfkNANKWqNdwL6bTYNIp
1rdht7kXUxGL0XOAmi1ZMKg3fnwdrYOzG7OxmbegI/+V3ugqiLmzGAxc4r/mnbYk
ESJmrVtv6wyZF/wj2IhYuKBFoNCm1LMD/MY0mITZFv118CHpv9KPqqWwOoGjeIXz
7K/SX2ol3ZZox/3P6ctsLCkih2gqs9UoWO8MZrxr5alEHD4cgxBqHu5slbqGWIHJ
UwHTNbvSQe36iM12Z6Bu+/jINR+o7aenXIbzonlAz915gaAcNn6jcAoL1X0alnBd
KwYxK/cy37kVKwoXNdJ6GkLKN6gdIKZh2lFvYJAodHQM8x01h5oUaRFZW2ECTUB3
4GnjrTRQ+dEPs7mJW28KqH4V3jUVf+GCwvs0cQv4jJF8948DxGD6IY6HB0mcFBaO
n1766YmOnywLXIKRYcpZXmDK9Zz5eECyxD7sUp2L6G4ckWPzgA6u4yvyM/pFG0Ak
2fEDOFHuNLYcE9ZjPQYzl0nhqf0qZtKDBXtsLDmts2Dl6tq7C9ePxgyyjvjnxOSj
4aGQeUNrurhQZwEHwrLBIGyhydO1DoIrez5XPPkvVDP7M9eW31KvlDcCoN5jc5RM
Wjy0eJvZHSS0WXmjEosUhopPKFpBnSbJDIFu4TDRhDxXmdI7l/izL/9xYxJ7z2g/
NRfZ2i+2yCb7/CcIeLDZGqU//au3wRO3ik7nNmMEKPytO9fprXfRJ1NGJC06YkeZ
TLOyKwbLGCN16S8mjnkoOyNYwVEbSnJr34jVlk4OsogMoUXwI9+K8QbC5qcepaJQ
0/tm/Q20A4mcaeV/g/UzaQwQNiUStuhja6D/n5Ig9AvCdbBdvcLHagGS+Y0HQb3z
ZO/k5sbXUOFTODYTDVYREn2/k/BKiLdbTo88a8ZqkPMGe+EEOi4BtXxyHpGO8l0d
+Xk836jm140JPh8PNAIaD6iLzWvBvY83o5pmdNQX0BbYelWAMV7zfFx8fQRwxWsc
6IHpjCvMAydKRwHF/GEArbB4mZg+auLJvW5KT/yeGw+loD5wIME47JZcAyH4mhwY
c71oljIoeiJypIUxLpWKP32DHK7SgRyewr+KXQkzRRkdi0THkatiyvMCteWAd3b1
WPQlrwnPYTVleLT8w6EOYlOBYNjOnJFinMag7i+lkoS1wfkK/dSXP8TUf5eEuroA
m7ErBxNBkGke3FkBnvvi5zwkaG+0NpNUd/IE6VWysYt5HuQJiCKT/2ubeQT0aZ5g
CVLJ7akZWF865bMn4L0n1HyKITk0zZGkuZbqypQkQBr7HwiMN+V7+4euVJAUTnST
rpo3k1teNYEP2Wt9n/HUVJy3Oh00G7PSnS20Yx1omUsZBeLMIysL4EqLcO+5H3uh
JOLhKIIJLZPj2a9xuXgPHkCONXiGk+gqpDn76FlPEpXNfaPLsW83PmxvLGM5wDNR
oyU/qmTiSFORtvcR6kWisuLZ50RHUdYw4v8m6TSNVF5omf4L1faMk9yRoEVJ8tS4
apfe/T/kuptGHFDljq0WkVTvmkoLk1P1e9OijpIq9CL4S5l6oGzlTauFb1Sm8q+m
f5PZie75ZFzUx5nrJOQxcPijNcMcLZiFX8cPuzkYuD5QrJhuxn2jskqDSBoxhGzr
3CvLR/3oOs2B5KLnv7tgx/I2izQQ0aAuqLDo0ycdfCnfNewVbrOHhUyW09OgQcBQ
UlOa9pxuECTBdtScniRcPImXxQauYDLms6w/msWo2jX/fWNOBMuE/Z6zXsElRan/
BNZ3I41r3McnjHVSr8sWsyXtJfOITIobT1YRrEsZXmFQ0ViOwW1fA4fvRmgBFitY
xKxm46+v48jKq0C6cXKhZsswu+qHBE8VaHdIf72A8vkknJJgNGXbZgHtimLFfk40
FfsYsoSq5jLKplzBw7Qk92y2IzwRYN496gdy8/pL8hniEKByeVlZB/M2AQ+ZNh8c
PkGa4+3yrC0+ClN0AfSmrr0Qx/AQ9dKksQZyo9yBNoSvYm22imCbPQ/DFY/wo7WC
VNTb4+SVWhBEnTA0q42qLPgJVttA7N8eaX56CvuMwB8D0tjErsv845IneZujiNy8
dUlnyWDlv/5PdM1qtiMRrwlBANhLsKF+bZEtXyB2D/w+CDE4ZwcdWaPXOxlunvJn
E5jUmr2luUqZx67/x6NZg7NffLAOQ/G7uIbNyfftd58uddfx60mWO85zBtM7K1ub
03kIlLwxsGyWphg3by+ez22wetQ8fwKUsemWJdRdRc3s4jKgk0RpscYDQizhUxRg
aGaBeDqTvljIdS6/9vexAXTV//ObdRsXqFBIdymi6FTy6iMwaudyUVtT3RIvISlx
YU3r4HOe79EHeHcyV4EhZk5V53WZSzSknPYw+BGxXNmZbcV+oP1p89cb8cJqDNS6
jIo7CrQXHeVZWFx9F0NqQdffeO2KBUDA1NiNHSwyW9vfBuTkYNZ5+KQwKBrek1MG
Wzjiz7gko35+UlMAkoTzA/JjPEJRL+VYu5dKG6efxw4m7jYHH8cXt7Og7aY2Zm36
lUwblLGKt8/Jj58ETFNlCIYR2DjnmocRt4DiHURDMK+D6ncpu6+J1rYHIi2bNO6E
MBF2A/Qnntz88eEZEtwlnaH2bsOoi26uOyXe5ZwCDbvwSI7iIFmOq/0DT+NOL9bQ
tyfrOTeAouFhK9puSAz2QDjXqsUoVYpYmILu4jZtJTyVpJTa3KnD1lCLDiiRzqNT
RkK4AXaokh2YqjFG8pl8w/8RGnIjyg3rDqounNz16abYi3wQRp6B89HGgivWSp6V
vl4riVJwK8JFqcoX4qMjaqmBTTIYWwgMpjL4GklXwDugIQyJWJRtHTAVRFQwWXj5
vXVcMN4laliKHyOqIUCvqRMEwfwNijeClIljMBXYTDJEvkqrEGZ9wo4eDwgtGfnB
OKq9qioYdopMt/0NEDNdvD8slWAxQaoLtpmsQ5EK7OFtN15M7f0N0EoyZaIakAnZ
rtuOw1g40rBDQyWx+WfdZF7vb90nyv4NQaVjuqr/HWliWkqgdYPwK14vdDIcQnkT
tvJ/UY0kwF/XLyVc8DyWdif6uEdwtlNJEryB9n3h80DL8q4YWYklM0IDn5xTyMqJ
30mwlznuoDCJBQ4vKG03UwK+DHwaV7jY3XDDmWFbL6OvbtSTcSarlwclZxN8V1SW
SV/37Am/vgTd0cxZO8UEE71lVkVOkQxZj1E5Ca/GG45GRvYEq3w2ic9VVOsM1Fnd
Gn8jXhi63mdJGAutXn0pXIpLfx6TZbEU1rWygUdXet1CeUX04kTmj1sAFJ+UTl7+
1BFTUoKpOzV5PfA5NP1IYOrMYKKd3ovWVpBiRrQTtp/wZQmrgnz9SctvpHRdi0L3
/XXEVvt5bYcS5aKzYL0bjtVU5QE7lwysdnc5CIolA/m2ifJCJPuzA3RF6vsQV8RS
3Q0BFQYQ19OLUEFZZUw0bSnvFfB1UdeQlLqbqeJTC9dEYlhQ46dqahxulbdl0t/B
Org2iNPTyE3PbmQGsid/2TNvBxxbjNeH8l8vGWz9I3775qm1LlQhwVwAMm+4IRQq
mQzUoFjew1a6IPlMvTn2hja6TYFtq5tKhszlLeG5JxPh0kk+ppUw95N+iet6lF0d
dvsPFzoUthjRDrXw+cusnampcgZQu1c1WQZpb5TWAQMgL/NMJXqGCeTOzS/z9IZw
EdNXoTuxfIAmelB7Ws0X6OE8nJtwZOExPQB9BxvoS84AlPTYTaZKtbrqpZO1ztq/
GlXF5UmR2E3M3Dt4Hb1mkuNK0hUp3uZQWliduLkc/5hNn4G9n5KAZBlHNeJhPueh
iOK9HtzUfo2hx6OjF7kxb39iQIThxTYHObyHCecfzUKHOuWi07WvLJKs/n0EeL0W
6j9LTPqNx9X/ZO5xg6Gf8UXQzROs0F6lSuop1p3b1juNn9I+RqSWqvcwkG9HyvlD
m7KDBJwWrGgoYthEg+pVZNHVxHERj47sC4YOXkaZ3BALgAiCNO3v2bqE7/MAzZp9
enBHY5o9A7GsXBVRmmUSa4c+hNSsu6iHZHels1abjk0D7U4XdkfVbyxXMJ71AofM
dc3OqHYVprpv9aymyKSb2yFH0cLJC1sH7IkiZWHc0wJKyE4K6/geysp+AhYPUDzn
3EyHvBer9R2h9As6KD+JH2wMKgrogt39Sk4EGGbaft5dGURoxJnPYu4tsk4ay57L
6tGu0zlUn390tudbWmDSP41DIT88k69w2i59Vu79xE3TxQXqwrmVR2ip+e1JybrI
5FPjB8avgoijSFQo6p8X66adA460vz+c20eGqpMggNZ08y/151aO6dLcLI6AIEP1
jDCNYeAZVQgNywKohd2cAawMfgJoRjbZPgOQLIz9ky6zvUWMJs8dXkLNFt60rwZ/
cP+wIscjx2MHKXQ9lvuWlFBHT/77fnECgYTL2W6QBETWDAanMRlqI0pZyf776WtS
8rQefPYvxT4pf8WiWKPFUYVLOzFVIEz7Y20FM7cIiSbSLbT8a+A1ev6Oz4t0DJOw
K4Tbw6aIu3j1AmbnSiCq4rHLrMVhNKHkcqNAT9puTWrrn3dmOiVCh2z+4R1EO65J
mukvCpxhIbJHqG8kG0mJ+3OxRrsfVBpf32wh+6HFz6ScspMR3VcqtbNTAgh6N8MK
tmn5dCHu3CiagK8/2WMp13Jc7z7NdNn3zADRgQ9AtRNw9ImvV/x9lQ8QcNY7U15r
/C0csiQwD6tZ1cIR1pFk+5hghFJnF9QSos9j4j2kUhpSlEU9pQDE2Bh7hSePPlfv
v5S3eeSUSDa5lSPTpW1IWyFLDQZhLcIyH2C8Cu0Kmj4fKDsfQnqBRBkM6VF5KIg/
PuEkMce7b7h7eJ4vcPwJlb4SqK1xeA3k7UqanFEBF89B4MU8lqyXJ7vmDUjB8wrI
z0gC0d7BTYe/9Cj6Pc9mZEFpvZq8HdhF5DRyIyRcssc/antXT33ApNiigusl7sBA
pZ0n1pBTsXUgRRtiIemmiWFJK4P4Y82bAHnlIMebr/rBCjOyLpaUpxCuUXOGg4mG
6/oWROgA3fGYWj84yU095y6DCCA8PZGW1NuYfuJIF6Zrwdp3ShZOdeV4J3cY0p+h
AvwPraiizuSnRaWPKHrhP8nPqDlxSQQoCGCqFwTLPAW7mpaNjps+Mc4+0RYG/h8e
TF/rDmNPJiHly2VlzhAcQlKzg43sA3wIPycbcGIRQy98SftQde07+jPEs/J2Erxy
93glk5GnkEbEMGOZzGME3XTFGQ0xrKyzmpWibuzqgZ0VLilwCoxTHPThyY0ELpzG
lY6NvOkl8oRY1XzJnIDz7FZvV2iRep8po7ZykwKf2H2d7Ggq+bLQ7/OIQyeLcvtK
VaTA6nLVCPfaYAKLTbg3iFElcoOK49Qjs0D3VIXU3X+TYxIYe++kNroNLrvVju47
zRExT/qJtbkDlB06P+gbjrieinC7AAZ3vlGkG+PfDIRb7h6uR3qcOzN9vG0xlcsB
E4nVqlLc0+7UOvuMLbXWoIKu+UHe12SUymycguOeJf2Urw3RkQda/mt2tMZGj50Q
g2G0EO7epGrRcGujN5wcBqeK7VADWzU8qpQjsa8vU0/iUwz7m2bWNphuuZLYvXwd
39u3IrmmA2f54DtRNrXlHqi0+qOSTzkkxiuT5ZeQlhDhgi+gGH/5rpPK7BuS4R67
NW+9j+DTqKFImLYbSSi0Li/fCyeipAu52GCVdI3YYOrhaVbsMSnkCpmEUtJTABHi
sH7nS9fuq27d21xm2vUnmCvZjnGFHCNNRNKqMc3u0lib1LGLhiKl/Rste6vpUuUK
fz+EkXBWORfHAq2fudZfBtE5eW2c8pi8nJxACDFwNhJcprI08TM1rM44dn9zFS7O
jcqeXiS5XnrwylUtx3c1iqgiM0Y6qTWfT46zOLCIioHWwz8Vtb0sPH7cvTOkeanj
xGCk9psl/T4cz9nMa7Nh8AARsSEJHIExcAoTIF18nICP1NjmFBn3CM+7zfT7zBlo
X3GBYIHiXXUDx8pU/ZUq9bQmkw30yaQPH2IYV+Ldg46yeXF30ZIpem/RWUSxaBvx
aw2a/zTlRlyn1pZBHcSXNvSVjPydjYpMTmEadrszVVKUvAifFwMXbfo1t56UKZbs
iRnxkPpfRfQzuZ5MP1RaTrv5t9ZaHm+YqqfpCVauB0U5QBuEmWNlY1qf9Y6Ey/pz
xYZ24hWnRnOBhSaT/6aY4Svb+5eH6md3/dBEWjlEIf8MID49LyvX+Ozrupkioh2h
hepNajZ7kn5kyudkBu4WXD8OjFu9IS5yxDo5gzwfV1veqc5Ix7YaLfjYBaOHcJEi
foxJWKJVfbohHK7AuPsbWqbaSBOhXyTfoMcFtNamPJ5tXFjYyofEh9N0zHgnMg2p
5t28KnlYjgNVgEdRbbMrVekOcBI+lOO8y7mubRQNR53FnLTjW233C60PLJrSkna/
JrqczLVagUUUSA/tDugq4XiaYnZvF0Y3PsCbWcSC2gb82rLlQlc2zHN3Bz//Sfva
/WKfS2l01BxBs93F7SiJIqvMRkvKRXZ//jrljg9B59EkBbHuw/YY/2czV7sH7lqf
dnOMDkvQY9NxuZ6nRuDU0kC4Xj1G5+dKYpb9yHFLBSVFV+PrlZ4vFccv4Bq1RtIE
1DaRlBa9ty1SrAa0NjYPtg75SqRW+LzG5I67cvKMOVQ2XMknTmHlO+pwa6i7PQHH
lcqiFOIsGqsTwlPQRhsaCpDwOOAkZzWwNLc7G4hPUEgW1Hrtf602iK9tFz83ezhh
DZRvoWMlY087B0vNKYfil4y4iX34OElTiqUi1yBJMV5VLos5FBFNTWDtwfM9zqYc
NcleGDzTDni0mu5ee2afN6Coi7iDrx0w/6rQUUgU94GXW6JzKqLs5adBvJOuK2hA
XGyxfZ/WShT0spHjyWoq+9N2CTKoba2zilh2nNuEkidxJ9+NeaZtroOlAUfXILUw
wRWPuH+qDMvGdVpu7RCEs9RTbGaBAXv7QJkukzkoyzJr6NU++ocJriZB4Pa9Coiy
1vexKnnRkr3Y8nq4jOvJGYkbge3sqVP3u1g0EHvaE5cGjG7ixJ4x21Hu7ufO+Jh0
2UbWDPX+MOc7DWszZmlQeWtRtd2o0Qv35hdaRr2re8IDE8QEPXeCRp7jtzevVPxM
HJwdoIBvD7d98pcZDt7X0F11ap3S2jINPk5uuw+nzYL6KIvyHRP/YsUwNCHtS9zQ
kaoOr7FV6sKYSrSw0js2v8YS6LmzQtt0w7HlbGWTpwef2dgwC4KAIongzXW04ZOT
F7eWJ9fVbGnOmlZ+fl5Pj+wv+ICppOtyDrlfF2Ud2sz9YUJsmL3ytNuRvb3ScPD3
LmUl6SmcEHlzHzNK21hcPDC4ApDWlOp9miq/3Dq4k0aTxReleUdJW1y6tvhswzsR
s+Ie0iFoSMTuARUk7qssrFhG74N3+Pd/YmtcA56SFA8abJ4MdDEgWX8GKZhqhj4d
pP2By2UJJS3ec/U8MXfjRn5v1evrFKMNg/FJRZW3BT4lF9tLac/S80QEg/0+Tjn+
WEuSfh7FQiCT65nm6F165a3WLfoq1C9A1Qf/OvSslsoxSr4KjTtJnkhnlpcIOQSV
9hnPVQNFPVQ9GXd4HQJzdhlzsnCIo8aTbpbBPxiCM91f1GXypxd0SIUkmGnfq0E4
kyHnQDqpk+Az2sgX6jXM4LTzvqYVbJ0SE/vD87GLHepXeutwY3UmCHFnGaxncQPB
PecfsS7PQ3tyOW4j/CwlJe/brt/eH+wdn1whNYtEDaZJHQEP9Z7+G6MlI1f0U3Ym
zkcozqqGGAXvG63oYIHLGHW1lJNWSe1wxMFkXZwML4pebFMBgDFy/wODnrCx/zL+
hNngXAZhuY/zTaLpeVasm5uvXPl/hm0JzhFAjwBjbh/YobGqNtSRwWVpw1w6bjBG
p87r1Jj20WaVY9r682IeHUCzQrPPx89Mu0v1kN5Rj87kxi6H4CcPjeT1hoBUA/6k
rd70KIcwGN1kOGKr1hlcJQQZDj2diryliYK1kjAJudXgaYUYxG1/CDB7AwRNsiXD
QrKLdX+vcSA/GhmhxHNJdxVQSYoO5Tmy6nSkrPcV2f689Gn3IG5D1ZEchinqxt/q
MFbSxTTzxdPEV7edh3wJkvjwMlDGr/LspGv7MOGeAqQOG5mUpIQyaxL8jYo17js3
YdECBm/q+tCecUrvbi0iTiQ2zMlMJ/Go7YvRZsEd2lXDes+OSKAeos06BxNv1J/8
sJYsin2kPp8862lQsR8l2bLraN9iHDWfnoZpuJKlBPQfYiuTgsIKPqVZHpZuVFip
B7A9EptOiB2ul8wsnuzboRWHjql0HkhsIx4rG4Sgs2bKaAHfbizgjsw2os/jsMA/
OMi37SISjG3BFrWDCwWjB1yXYxaAfQBBrbpxxV7TqOcF9IYIms2Bzl+TSH1SC1JZ
6DdJkXPMyQEGYnJn5z3KjuCjW9s8b1sOhQ4OMevUZkk0oAsTiKGE97416VtDiI+5
/iTOkcWE6D6lLC8p92G7LURRxU6I2TUwXL4EFRl5ORz9Z8DfykMaNj6nbqsbgZpe
jWFYnWpuq9q/0oU2t7J2GuE96I3TvtVDrJsvMh2OTTTAhuwNxAq+udtQw2PeXGcx
jLnqnabLdFI0fOon3h6spqxqFaxCN8qGLO7UuDGAx1CthDrXYA4GMfTpn0KQaF9q
Bc58E/LZPcYb7ed3WEBEKh0Z21v2bL7C23ZBZY4T1EK20JercnxepDKBeNwNIL5O
3p3e94BlL9RO/6aFlOBWPJSuUhVBh1r6uX8JGzebFNRv7tWPrZEtcq3OvrOQ9Tbc
k/FXI0ZSBzcmMSSoMTKzOubxDUoVUvhnQFCFmpiD+nQQstMYrD1olKIT3saouSM1
ZPegztsdne/qMM3az93YUOx5t6IAMe+uNtk/NKpYw/zk9xq3osBKoWzcJ2snIbm2
iuYbaAPbja4nx+rpOBvV6yWQlSrJCbV+RlSRTyqnWSPBgiE1DIMkkjl2HDiFJjvn
vQhaemUW17kKJgWJJ5ulMkGdWjOUFEdVqose1iyG7oGjeNd3mWDf4dTKmzYXq1pM
GaM9Pd5vGHbqZjqbftbLje2oGf2D5r3dFYTl+LEgfuUaumqjnZkvzdXNtOtbtRQi
Ugx6nss5q/aC12KYnQVB+YUX4NUCIaoGmFz8DpZqId9c0U0wNOUXUuM18NIxnXmL
GU6CNqafBarBrHumhaPph/F+tNMj0XfpcjxRvb4ZzOLcCQsT2zh+pIPWhTtz1BLt
rn/g9sHVuZMlduCgrcQqhj+zM+si/VPW1W+Luj0/YM5zO64Fv0/SvGBVO6GrV3aT
DRmD82G+epf5+LplBqL32r+NCp//hicGPeXhj0d3oIpSH55kPN94ERorjG0saG/h
9JyCe2nwk5fM17K4YoZOjh+/uCces6wnijUboaLGa639Gd7emxSNIF0eyhgyo+hi
VWQx4o6wKUs285rjL3okM5Dgwv1pPP4pViMGQtUuDLZcq7NxyIqSRNdPbdMJfBbb
zOQSJfZxLKq5aflMugQa4N/9bAWXCA6hUlmG3qdc409jRLHWeXNzRTi+IPqsfzPU
GIMAbQAt6PJNmQ/1aqCj6KKGCN0D0NAiSfAVMza8JeTDiMGKlyjEdYMciQNrAgGA
PBSvR0An/tBs6GpSxH++8p7eoMZAfYoPIWVgaeSr1QzjJDYq5/enpdw+NP6TLChg
ig9sHAnL7JZ8HJQnc3gedBiivMUqGWC4i9BhWUDtaUkNkozbrM1Hc7rlF55INghB
0ij94fabIzwP58/j10/jLrsin2DEJZutmARGFDmtzS+vTkacjh7CwLtQr09jsaBi
SR8vTUglkqtG6pGyb2UhnHcKzMUwKfbPVhEhGz12w3fn0cFP6KO2uFlKIf1K7DXy
Spx9M/STyN8IOGNjzjEnkNxAzYKaQzjyp2wZ/HJeE2AZJu2Ml7rSOfEkwKQDG9xj
b64V8BPBRe65fQsLcvRCVdUu1h9cTzAfeh63mW5ivm3g3+UohDfPkZkNuleGIjNL
2TnW6O1s8f3nRK9cuJN6ArCpSEqsGajMtj8t69j5D3I2HO3w6zxCEqw4qGAipzpR
OZmtSCCk3UYYHJseLZ6Pjn/gCdv8K5hGGDNEtYbrJBBqG2c6v+Z4Aw6HTVTK5QsQ
pHnD8wr4i3jPwLe+M2hMFJK4K0SFf8GMAMa1c3AK1xPO9Ym+9k1azXMaypoZ/MJJ
SGq7b3rGvpapaAus1C7irUuIMd7R7m4+VQDxYChXugGsOYT6hKbR/ARYnsr+a194
KSJxBJGJndrHQa96dcniKkkC6dpxxdL4CvnDjMtEVxKmaKLbYlyugqYFbjEgbFdX
bX4PSNnFMvypF6Ty3mgQQBpv+ipt3W0UrM1gLVtFNH5xrAgOHOryfT1xO5Or7orL
yiWrnwpuxk6EZhzHqtPcswg4nvn7qv+I5TbgFK/awM64Ff9hFEFIhBKof+N2Qy/X
0EDNQ/HJk9PCmdNULLQREKkWFhIt/kJMord9rAmXkJu968bdHKXLCIn1rKSIv2HU
jwTwj+/sTX5bwQ8ZUNgO8HbGUxfGPHgZSOliax9GEPUEaJXPgCDbF6XxsUJNemSQ
cXDTXnrextgC0/Edp2pooUfueGWXUpidhh8e2LQteHnV03BMc1sNYh+A40msY08q
QCIV0Db5ZWVkYjneBIdrvQnIUdSghWHnsedv0tvhHw8GQOsXZ8iV/UNS+XJP/wvU
QLMCizxXIWvGMnRSpC9s6X5AV4Rtd9Np8JeE2GM4y69enHHpv45+RVEL5/sO2deM
jPv5/9OKFmQoivG023WPv7KyrA0dHWqHwOppg+DMBrmyUBbWDEVXsKp7Ax/qonpg
v9HFECztnJoXJ3E7guAAgeB6U+D86c5zZR5MEN63cp8o/JtYb3SfTqpnNCmcXlT0
1pNhHq3NEjPpmEcZjKLWVz/Sjmm6bK1wTSfslJPJbIfy1ZL6sHwdHUmoLxSrfAIF
8nyKoizJBHrgyq9PunIrF8IyFbqv6PXHrlUVmN1SvDVbmdTVqV+8Xz/yW8yBIEss
mkIcqV8AStLv+ZfD7nt88V/1k5crZQdQex5uizKW3m3ajDqBTEMGmazRiDtPuLPp
LDDbBXEIO+hYH7tKLDBgJS/6x+Re4lRzAmrqQnJnXHCJyiXfSKUUYnRZilYqgKGT
uQiaRW9dpT9anWDDqm1IbgP7rOiaWD54Uzcig98s0vg90tV/hNyCdP0oPCSIEfI8
/QYkU3qBnjOGIgW3vzwmHbT56gF6LBp5XKWmflmmqou+ifpYZs+6BDWTVmLaGKzX
MRoESqE0F3/YRudF+yDHSD82/pybyGS82oMmUvTci7Sb4AeT+hvkxh6IdlSFjPzp
9MJnnBT03W5YPcGdgqkXQrTm9eLA6qUg2ZQyHNQTi/gKCXV+2Ju4cP7cf7fSIZ2j
kHncbw2zPS/wt7Lf0+6tQyWm6NCMMK3v786+XJFp2q2jz0lxCIL+vRTdIQKKQAqE
P7sJWB0fwQAQigem1GQNsNkrznjNpI+IEcvmF0DAte4xHQxAdSKNUQL4weNXN/Lt
Df1lSEVZaSNFPQcb04RtGeVmA7YeF65LeVk0Co5md1+GJksbJ3pO/P2uUeZzMINg
OEpiGZERNjLRGfG2BijMnKThYAz//3c4TiFvlYxzAyTdjCcZymQXCEie6qff/36Y
38c3RRP1jVjE70Hj9ZByV4oZyU/QyOCPjKD+4TuWSBeWDAAMBUDhggSBwpw9TNtX
2II86q0k8HQrHxfM8s5Fxdz96109OX49pds0Lb4XJFBxPbV6XZYScomgT++kNOlm
V4pnY5XCsTf+/hx8stWwyteHsGQ6moFOKc0SpdjJgx/Uk4RfegcvmC0tVJdaHYv4
9p2QN2Sz5l+OOZ/yBzP99y0MUtFhzZ/niKXddxOlv7FJmiVIkOMWXifZ6YnN0OpZ
gjUenZTzBjqPZxYqs2jcRCGzGK13wdcOtC3zB6W71cs3eO805I4kM4GatgWXHnNM
Od6gySY44MhOE+3H20bjmsEZojSx7pvzKcILSGoWIAcYh5DOds4kpaoGnTTRAINX
CEiJgQKuItOQ2VaiLYEwhX+Q0g92FmT2AKCNQXTOoRE+Yyr8dLRYLnfuX+7QfQ5a
29bQoreg1W+64mjbzUtRvEbUswOHT7Pb+cVS3kU9qQ4CTbIfnWRbpnRNeoB2vHfJ
EAuiXIWfPnw7MYh3PPywzoxMA6tKDHr2VJRxU/lNdAmEteGYmDe1Hgxu0Py5+aTy
B4pHVfkYypw1bNwmfexOr4daA5mF0tgTng8yoMaOn0YAfXfEsUn7IimJezK8RgEe
1Adq8wlXR4F4mM+3xGWlxnnO+xrvGdkSI+iRu08UjVB00NAhH9LGUmKPPX2epBfb
PBPvnepd8awS6Xw639PsTDLdw0aDtJQphfGK7UHFq7bigPc4g1s+IwItt/5aK5Dd
hrQq88kqytCmIi/hO6a8YtjAjyIs3U36BW75ScKTXKbeix0RM0whdgQ3ckEe7egM
30g1S9iW2hje1OsR9uN6iLox4PEdqA4A2Xw22F2H4n2KuLAlULyyfeHMrwgtZ3Mf
iOUSGqRwuTCjKQVtbWm8YHRJzgdJzWQsEKHf9Xe6fe+K9VdiikZixeWWOBcw3Zv2
l82YP1gtYAYXnTMIa12qY7dB7ixALWtfgYNep1XUQBQkwynG9LoDaJLlc2wOKP0d
5Yp3Bcgp5OOqt21LgOAziqJLwyp6Vaavv4kh/WXd8zoBSp6ynkCkLrBA+B3SQ/pm
COJM+bLmZDtSTjfMuNYW69oQAZdARmhNgeFX3uQf80havSasVEEiVlEEm7S6qWK5
fJ/9cgqQeHE2q+W8uPZ9RAmMTo5Bo0611WqTVHwWk/cKugVQx2LCyAibPg5QXWoC
ZNiLh9AsxAhTnGEfwNVqGFHnd9kpXn48aT1GgZsO4REizpLWZuEe4Q13GnNIzFJK
5zeIXAiXMqSf0/xjo9mzEMnQezfnRAfQzy4qPExCp/p4pH+mZBW4JYTaNT8ImgCK
jtffTAZgtzClevi+z0vzZJvHKwX+zUb2NOxf2q+Qocz2fGlH8x+BxNiFT30qU5ba
Wfh+HhJylmewwKcwJsfRo/PLJMkOdKrLvD7gtorhCO4XIJry3PMzoU5oOcGpGoEs
S9r3R/PRhMHx7qeP9jMJhmK046A94lhccnnZDCeo7pnm2ED5zJBBmaxQmyE23g/F
kuVF0z5TsHigIoLxp6bYAk4bejmQg+rTGPzgesfBELYzm3A4IOwRziQHnuJBvqJ0
3Aa3kESQW3er2RBrnf2WPE+SUmXHM5RzAOFQNpRh0mTIqxt1OLkxwMEHzedbarMy
moyslR9CEfKGiSs/RU97BYFcLbqJB8DVae42QvqZo0eygvUxRO38bi81TmbM72BE
njIkfkjQx63cvxaaEG9VhIBBLUV/5EWasQ1m7ZJDTjNxVybN0bA1EdK+tg7ACBX8
7En4ln5yGyuCn/gpd7lADVIPuKUxaCLNZQx9F80PR0kyE/hb3U4fByqEXIwxXNgc
CI8zRmL16ln+SD0bFOyMdeYX7bdvQLIFCOqoEmjhUUpSt9n6v3121Duft80GVaXQ
pYkgk9oVFnSsXI9bPSM1bZm63Uc0q26SItUawZtrIgIyFtq6p7B1Ih7b3dzCv3ZB
ztPNQa8wfVo+wUmwX+ZRCGhFaEmz7ECY6v0cLoxtbrckANX4JIpF57znueTKpmH9
nTLL8DKtKODWb+BipZ1VqmbGbXNvRQjIDPyKL7YlE4aPCMsrLH0qpisgCCg7/l0R
V0uzGxItxmlzWu6y1xreheyW8kiujEwqo/l1VRrwI/vANBeFOVru9lnIbdHIN6AO
E2gzl5a3Gvxag60tqsY8jdrwCarnz939mNSdeKKYGAEwy8wbq6D2MuIPVLwSVW0J
2aP3rP6AouxbQQugJhAUI2huHmDgIVzkQ/GyYHgJ0Rc/cNkBfHh+NBlDKponz29u
AztDWueKBKT+i6prgivw4aTozKgW8fu518Y08a68uWl54rAlsiT8Oysy0G7+bRUT
o8goRDilsU0IZzJmQEvTFmTJU8Lj5iQnVAL3J0T7YBENDOITIYWlyUbPYhk3m3Be
3Fogz/dDIOEE3VXt2QGkfRQzruPxnItxZHAu2PLsRb9JMEcv5c35pIqsrl5cIl/C
tJMmwLqdaSEX3wGQUsuSSurlebObLOiFh5pj7HxTmYDe4xum/4HTRLj+wY568eLJ
6IkSwrwTW0MAPZIYqUNZr2jUpsQJqYtgblwuOic0kHJNfT9GOFcP8afc4Zo42/EY
KQeLNtz5ZzXFDZcqoQMPxPGPgCfFwVpkgUDjhlJrTUx7LoDk6foj++xEgGb/KmVo
upHA85nnW64D6hSnKPI4mWGxOaJhAqCuRarOlR0gjBEZGOV3GOXdiltv5J54vSds
cxB4O1Hb702A7NowM0AiofD/KxHA18+LyFDJGl5ibUbWEDQKEiSCXdLtCsDI1ru4
Yoo3Z5lF8/oRWMZWU+FkV/QQ16yMKY9cpk0G8gBEJBqkrXVKNfXJqkgO+3oRJQpI
/wHxLqEX3rosKTQoglyqHMjlYrgZW2HkCAgVqLbeLJ82ojgG++4zdpOubYitgtA6
rw7JODLIpetC/RIg1+qNQwV+0AkH7VEugdGVkXW2qVSL3+g/+UGpn+2+zJothNIA
or0rBBw59sye3cQBvbZCg4G6zmlnqJ2l/qOqkjLiWidnJCD2mdn0BrPG2LfBkv7Q
qtppBSyK+HgkeuJrxg7WUsxDuFkYd2kV+hUTDjDGk2Ij/UgUWTKTwfEaB2k4N0Il
bnFpoNXBL79gB4/YaEl3U3gwATqsnvLw5fMPlkWYWuQX2d+2DxZ9U13zpNT4LTLy
vpxpkbPPJ56xjrnil+DU0tfAApFWDmC9lHMTc6ucs+s8nVbi27FnuVOg7tqGBZlh
bj+AmzLiM/b0Y1+ucqyeDE6VXc0so4gQDKiASl4uMo9rCE6rjOtJnAoKeMX3Mha7
TeWbYv2SJ9jbJEQm/qHtb/Gp/h/KDO6uVFs5X9OA+OdJUnHpw/LDEBIgvOtqb+fd
s5GMBOV2N+daBtUmdo4VfmNOhaLX8FhnEN8E8JEpUV/lYXCsmTBgyo4NOgOdQcb1
hkRkvVZ/NwDkjuUNrZppCWwyQoJ9KMVhuTnrFiCL0gLWXLJeGJ+mB8TTr3BkbkVm
0mXyIKbv4ptBtS50fem6KmHFQ4PM8gknA73u74+0G+UUkNH5TbB65596YUvN960v
jlgsazwsHHwTDkLq4yEN48xtGp2pI5mOrpanxDNrvEgDbWXKBGlJ9NBFLgRg2ISr
uAYPzFCOZ53fRZb+O5b5+7w9/VnA1kRkvsMuYMII94MDUYxoEJcFIK4cfO085jUK
EHr9IjDab9shOgPywJi75Cb2CFd2gyZIy7w65Xo+u/SKlEO+FIza6rX5+cwjz0Cm
VSG744Z+Fx/SPMHtGWvG6gkyFnSkXm8cCaPYgHGu28s7wQ7C0eFBSPPcSv0usl6N
2rHO3v5yJMU1JiiGCJe6NEetBvHuIBbWpYWOD2coSdfpXL2PhpRhRHxuxE8WPuIn
BjFTTJlWak9ToiDw+xG0ofEpbGMn0V09yrLFC0k55rRA7IEwJwW0+yM5dDa0x90r
8Hs41ez3c5L2m/jUvR+Jz9eT5FXZL56JGxpTR3ttqJykQAJdVSJ3Bmf8njaNyH/D
D7GRlJiurNVVlAY/3pqeMbV7VFzv117Hv947x2vNCDLFL+N0MlLFnIAJkUGebtam
zjAhiYiH5wnYdIOh9Vn3FNq/fDhd3KEwXtl/b8wyLqil9HQhL38iyz5Mwzxzi8rK
9NDD30Y/DdRlBZv8K90kWw==
`pragma protect end_protected
