// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:46 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eRyf38HsExW+krm+ubQXDgm3OLanRMUFtM6LpvcKn/9AwbWTgsDrO2LoEu6yzLo5
676giEfDylmltkTsKQeQcihikXjWJ+4mmPaP217dM0pxBkdU1ABZy9Ij3jtOnbEE
oTQ+K86e0/WXwXcoXs0cEIYQFzDBCD7ZVvuiny+eZZo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18384)
ntNUisU5iuMspXK2uRqxtX+qTeUC0gtaiHrKpfTKwUKCmJLLoryx694OOmlOo/ZG
TlJ3MI1N2lZBFoLg/w99vtbthvW73C0xHiQOmjIhdxu5bHt+lNlWNy0AM3J03D2A
C85r0H/ShgwcZ+HZTOky+DCWc/wmKyN0gYJ0agjZu9kI1Lu52NWQgfSN8uTjFmdI
pNEmgGlE7hwCacs+PLWIsrlPhjl5/uEmqZLbZ6xmJxjR9rE+ttmAYLm3JpiSq9we
StZK72gJGYtiZa0ldWM4i2wJz/aTQV8AvsVdEFALpf5Xc2UvpXaQILFVJfvV4/nT
paOXLeLZHfRHGfObXxgO5jLgm0uq33OsXO8TzWJB3ElPa9zWFVMZzCmQO6ZRFHHb
fEClZiFQ3ALme9vHK+84/ro9XrQIudu7kDTjDg5E/eHaJgoS5xpA8FowqOCN6Zwo
Nmc32K20QKBQQQSILs3GTLOSBdT/4O5HOuJ8iN3EkaXOh/hO6HXFk3JlSNFDP/XG
FBjyv15XrAjo+fQ7rHh7P6DDOirMMkN+wJgOqdhEK+GyNm9lYbmKEoVcBlHSTiPq
NDSgtoIructmyuGfpekHcza8K+meCM2zaQShIEjDMWKKI4I7vOKUg29AJ8k+REth
SRC9QnQCZXbyy/aqKrySEF+GhE4GeKGDla5y6BQhAS3OJTpYXf7vJedjNac7ttBj
0eA4fkExpRprSEJE4oieJ+Y07Uwrr413d9hLfR2ZWLipbnBK3Bx4slP4QU35mPHi
DGMTGsGEZfmJF06a0iArBCJ/rEmb2FzwlTaWADcSX6VHXg2N8i59EbM95pffeyPN
BE+snO9CroG6Dra3pVJuM/ntReNKoXn38S4Uxh66LR6Mx9vfbfB6A8SBzWIy7bwu
bV3Xi+9UEyBjUQBb0CVN8SAt6upUJ2W4G7bx/Wl8fonegA6pREVaDqZNYGpsqmYy
bjO70xkJ3RF9kuoifwO81+q5O3/SD38epmcVkjeLy+GacBaso7qczNYTPFkCkmAc
b0pt/qjkrba3JFtv53wVgIwF31dkb1MC4b3OyuIpGnm+AwPuIz0/XQypc58bcx7j
AkUEgUwrqUte4gMzLuTFDk8abhQrJY+2N4SWapIO8HE5TGblDi8mLRII0825EFYB
eNs5Hglfdu6HoYsS8HsDhMCubKon5hBRFMtIUo+DqTpC963HDu22QTIs4zvkOELz
eoYtAsyjGhTitSdFfIx0b4dkkkqVDzjAOKfUvo1i4dXezxP/885bwQgO79cA87dW
IlNc357vNVX/EVIcbNgLWmfXjFd9/7NIk2f6H1QBj/tZz2OalNE7enEb8L21B7lZ
0GvSiSvfyi28Zycgev8NTLw9iNeSoserD9AqW6tVtRz/LogzT//fbtjBY5CsPCd9
YVj3DWNycQC0buj0l4lGM9lQnTSS6E85e9LMFdEgyXdGpKxvP0BLpCn9vzVkr+KC
UykkyN9AIW9A+elC8XY2OUfsTMFzOPx79r0dW+5IKbCWW6U1qvF34YTOTUiPGzgt
VzuKiyPbx5ohLiTtUeaESVFvNvxA/NVfYWnPM4GGlOJFGGU4SjG+zL8tQgJU3ymI
cU8Ij+MJvJm0kLNziRei5VWuo5ffw8Z3OoQIFdhpogZ0bIFSDlTlZqZyfqtWCdFR
aB/qAfNiJ4lRtvYCI7Mh8WYkf1h2KMUGiHOOPJ/xHfw8/SSA75+wKiSIp59EpKT/
n4p/+wW4lqunCGEA1rWcMmFWMEqygRAoF4xlxYC9Am2JGrgO/53YXlxBe0RQJml8
gj7jk/117ppvpDwyiyTaw3ZMNq3i0t7WDBkeKtkgz9O/UGf+TKHlWFgBNVu91my4
1m0bg1PmdiFeWjyHT3nfksnbmz94Y1mAM0Qv3Uf1sbiiSbLtxEi4tB5XetqQuDS+
vC/8C8gut1S0vp6cI+iuSvpfiVv9dYEnzq5Q1NB4KK4D50CfB3EKm9eKn0r4vd9E
KISFTHscIcV+wApeHrPBcx9O//UdRG4s7eZckjzmMJ9WJY94rVDYPLUdbVARHsYY
0/yPUeEY5AgN4+NdBv2AgY7yBqoZz/PoqVWyMr9InrOhtCeb11aNN2HQn6c+cWhu
LlFRsyPHKzK1lbN3cEe+2TtR7a2LUokHJPfCcK3QGTeKJYzx1OMsZGON/+BmmTTF
yNtcm4zwiKxEpvsPaT38kviwDiM/vEfHERahafiiq+a5WaTb56Vj/4Oirk6aKnFv
ypbCVX7YYoLcjzHvlg7jcgOikqnhddbxTP+g6YpEPUOYz1EJMw/qMWRtBfrUm4YJ
ap832wuOWWwiSAz6CQbjKUbeSk6q3j3H7seKwfZqX/SBPHlXEif8aiiOGq4CwXx1
ZQUHgcofm+NI+FVD6og9a4Ac3cr5OVvuwdzZfc/JrkS6PubEOLiLGWi8m34ArWAs
JpPRYsA9hxqbEGJ+/Z7HqUaZIyIGrgy6kwLUuZCiwzNNAYBWteZD1mizuZyStAyL
3hUXgVniFHRIG6MkvEYrbu9hGppeX70oXjLXA3nZIsH6A6yps0GYHDqjK3dLbR69
mKdLHdxVIDmjhIIGHrmcMOkIfuTm8knByEvMu+vUE5PZxSdecg6kjq+DUBJgS5Ju
TNFLAd7L4dWvsY98E8+nMlve+QKnVrbDtptuzako3aNbazhmmtK6F5RPSkJzqGuZ
pTzrBSo7cqWLulvndpYwpMsFEbiZwL0bzhJQ0dpxeAdkxjGUWFP+WbQF8+fCeOzB
aNqEfegU2h2i2KhVX2dq8mUVodY2h6ngs+4WXep1TS13VOLMuvKO9d2spt/DpYHM
cL7Q/AF4Ow1QaJAkYNRRZ9SOJ5VSYM9mDBcayQF1P8GlIxcAydpPC+JMT/vDclyw
PI1em6COww7bQ+ACFgF/8URhgmY913bp8rK7Ezp9qfcp/UHJAGYVAL2MHg6qURV6
kihlVhfJWzWy9ElKlMiahERdBhSSioTZn19pQyFJXnVjMIxrnAowUMuXZuxRjFIC
hgWKJccJawezGkJTNc/gdgEbz6EOKCfTlCvzfTFLSm6D65dzCKzHItNVbJc4gQA+
KLKPY/btoqR+CC8SiZzbGZzZO64UOYnaHaIKiELeTr2NzmWvptNWvw5o+92ZhKhL
ZxsY7YCm+9PmekcDPm6BEoj7eNyNsRpDZ0Xc4YNqmLpcrKENJytbuuQWBhAgQgx7
sR9avRMGdKa+id72FHAEV/qYHCJdKuLcukK73h3EoFQsNnO6FOMXkeiMwYJ1N7nG
K0cjcjFcVGtPpc/MLtPlezTTYntVxw/DVJCPjVyqDC0lwQHXqOskopxW5ooD42Q2
jN8Pk7SRkVVWL4U4W9cG/jJa5H9GSC9c6P4DyvlrDCCZ9gBFjO59LfurVFRpGB68
gslSGVwsKK898Tgvch7vknNwfRdM4SqFwKQpdPUYM5lzkWjtPl8ps1UDTU0X8VPF
rnNCXgo7Npra6H/inwVvi4sO59pNpHHQj98M5MP1pmuldChSLYrbg/xCA2ndZKUF
catzGczPfu15NmQaMZZ1wW5tjNSZ7GvHYcgLGwNN6wCLsry9EyRq1d2SR3Dmt5d5
9SIQJDfQXv1hbmdaD9DfztjdhHE/W2K9LcwbwCvjLHl1oXdYy0KWORhxFEwvaad7
7ZUC4aflcOBaBb7pZ8JRxTqpsCJsGJhyR9tw+OmjXdYOL9gwEsKgDDH7SxmGUobp
rylzxzzkPYa3IjnMBNQ/hsHj9+PjLfOceWowCY0QNiXKn4yGOWZB5APLZv+slE3U
T7+0tBr/WRGaurGXHtgTmX9Ef5C3/RKwBGbibgvmS+1lYV6QiySUPgXMYOuO79H3
OhocdLbxQoPzsTNvvxxmuHNPoqkmWQBiG8IpCWUIElwcXaTbpaK40jzHn8yFW9rz
+59rr9lwEwhceHgAmyNe9Fjy2gmud9DF3lgKFxczu0VALl3G/z818o2bV4Phg3L1
/zUYPJega7hvAMYFhVjlyndyZdvCsavZkW2ZPFcx3LXrlJgiSt0t95pQT/V7OzjE
X3d3qlhVuwXV+OW/1XRzvWL65BEPJ7jSSKcTsblJv3l5sjZtvkQh+oHGHzCTs/cA
8rPhaJX9O0M5XpKVdnXES05toO3PQaCSkMmlJOg0CpmGsi2t0cq+4FSALEIxC+99
/8nVv26+FTFbESIbfxJgit/wJVsMn55Dg4E87h5F0cr4tdFWmGr208Fl8gSMHzHB
9TMRzzmbEHB0dz+8U7l4SJSswADVCJSWOiKIqPp/6Mak2+VAkgrOlySYvi24+Ybi
ER2K0r7O0b6+WbOGuURaKt/yzG47fqjYKPqYqsphmk07PHaeAtppoSyZk2Zh1AEI
oBW+JR77wlBAmrKIhP4nNShZjtmlLdHXZWaWPivKt6Ul9eYEtyT6mf9YsglrdIVF
ZJotvNuU4EuZiud4CEhxl2BVR8KAN8QnbM+XbXSp2faMcMnClhJwRoQ0+syl2yqY
31/zs7C/1mwCHdMJkqqL0iG3ToAVjwbRdSLAyIuhmgzS41Jw3A47M+lkL1ZCF2/S
bC5bHdhecHQbie+NTfwfLeAwwj3EmzTvl0em1UDxdzbd2ro0wWIeOBmTzO9dGZ3x
/tiEjiCl9jw9mybczbDd4FVdq70/fYnzVpNWWtQiEyWg2sBXIOfaCeZ9je2X/V4T
+VtAYEGUPIsfVgqbkscQ+ZwYOH7/0b4iTEgdC0BFoenYhjxNqnHNctkmd+je1BxS
DLN1g3lqCvibQspc6dC4DWxEUen9sZwvF2KHYHn50/7kP0eCkrJkYzvReU9muBkg
8BynrI8K71yWcd74m2DEFS5g8P+F6BqdP0J7F5r8PeB57SPoprga7K76nZmd6xSc
ZyIxwTAoTaWVwIjPBIkNYNKT+aREpseIQCylQDMvo5d8JOOaKbC2zyAuzrhb1pk8
jyIGufrxeihXUg3/ExsucF4DzobfMZFM4geBoLAPiHlNYBRu5laoxe4WTEXNYQK/
qILYMRVCPY+6TYvqiLyihYU40jt/J0NkeHNRaDjP+RNhTBdbyhZpAvPmDqV2zy7C
SoSFIJNTD0hEef5YYg5yiTbpphSFlXdWJW+Us8sTtQ3K59KmPttxToPL0VcXTDso
gFOy+jMb3qlC/GOMqhFZ262Ymv55arZUsCANmge7D66JcaljVmK8Le9KmI6KlXRl
QHnieoJBahjSyp8s5EdQLWb0g2qimHKcAz4JTQEAWqophuvnBPAEyBuf62s4sxBj
ZGfRaxY0tdpCzl/J1phOwPvr0g8M/ygFpmGskPWUXHPbdnxQDSQRMUghgvw3gtum
DAjFC0uaOivFEogOOZHS7zZU0cxg7w8p/O8H9YBDGPEqV3cCXq1azNVaP4FjO8A0
idRzjhEhS+nqaUiB3W4QQCs7hHGEpyvsUALGA2ML34YkrjmxLDkUhi8a1EVUI9mP
dlorkzOAdtlqMI7j1z99Xzr9h1K61fbwYiVYopTPdcV6k0GF9pgRKZE23GOq4JfX
zmXMyLghDQCgKLGTCoP3z9SKGCV4gvC3I0CDvMzfxMCsyD3DONOKuBdqpJpseCH4
MzsvxxAq7J37AeqLzn+dXEnf8GECXoosWNPPmXvKHuVw66iHuIIaCa3VtZ5zuJ0V
TWBIRtl9V8RSE4OchhW6qcytonbb5wvH2mtUpoZE8wqvatbKS+TDVl8HV7aCqUTc
PiF0FJrKK1EUicujmnRMTcWq+K1IxUOgbgd6TsoSvB4DZslTfzB1UkNyPdkLFp+m
fUD7zt+66yIpB+TFf85qQ9YmGoAJhMq+qPNNnNMTG6/rGPqugO+ucv8xXBUjRg7C
c2YgTTy12kWaOnOhF44g55efjOyANRNZyka7gXpPpYe0GTrScMQ3CSI9cRFafMXa
C9Fxz+eFKq16xG0RPSicZuXfeqCZm66vDzdfpgBjucdGBrD+H0yms7MMaayXiUGe
GXeex/KqHcVhNE591e67f898f8aT3I/ua/F2ldPInC0rAYQ9I4JtvQy/YRy6mZnx
zrF8AX/RKwXeAPhANwyJawXazZRijfCngRK+0eOCjNDOdtob63DR0CLUqlOChEB8
dNiAu6NgOr6nALClumWrdG6iQ8LaWQ9SOKBNOt4rnWlVDo1acIhX2WGX5CtJXLr+
lGc3G+CGdev7qupx0m0PYhS5tPi4gh/29KpfnN+Y9bLTZQfcX7/FM8EZPwSXlZPB
5gDMTRSvnJFhtapfOgF6BSh2ckCK8rvRGT6bqNGlaSwJzUtcImCifA8jSPv5hizK
npq5VaHpOSyFfc1QBsmWUmBnFfNhpITTw31mT1Q3DtU8TbVBcANPSTfKe239Ed6k
d+Qlh/elZ5B/jd5t9/5hVjt4O4GJ0zg+ztlL5DmXSbRXuXtCjgQ5AhnFzPF49P32
IQkEqcEqnI3tm4aai4Dk8xjPHNnqKOCUhNcSgzF8zJfyfk086k5AxjKIH9gnSP2s
M2jHY7lAxahb634cYXpMDAtL9BeiiDPF28Rn8uOI3lt19W0vcbXJWrZ3AXcCy1Aw
cAxV1m6ZBWVc1Qq97a5u8yP0mDJD1Pkcd3Sw4Bi0cnOHVfYkWK6vTFJnErSnZNY8
GFGBc6qqWy5lIdUp6rkSlDmKFg2XugticRVvvq7GO+2Ni97IfdbzTwgw5PyYZhMS
6P5MJNJLkyms+EUXYXR8afjNHyCsBCEwAaoSG7ZEHcJAZjBBJnHJXWRWouJtxnVs
f52+3iQMfAwRUF0cmjQQ+n5BcWRXTXrP18qKs1UHWSKM1atfGw6XC2ULNtlEcOFo
7qNx2oyOaoT8I3qaYrHtYozbUJ9AqNZ6FqszlHwd3T3Uv+vcYN641suCvTCVa0hp
Ox3NR8UhHJCkJbX+XFiBUy+D04FBL3EKhoJXkQZplNYMIw2EB7KvwjCwfkpS/1VY
iKUmeuyK0QpkPJdQ/irFo/uIr8Oq9TiivCiqs1smPnkTMppP3bVWs3dJU5yftBGW
Y/wGOyd5k1asD45budpL1M+WaM2kdcnG41ia3DzcqYwVKtUz49c8gori+AzdbbQu
X5TccqUIDSNteGaI/Sv0C38N3pKQ4qxO8jvx/k5P8NEewYq0vU+tNf+DZYO4nCtv
xLBlVmoMfrzWjthUEwu3onUZYclPKbBdpnNO+vjIesTvbnlf/tXG4fKerB2zhAPU
XixMSUjf9ZjIgpnQjizR4EM0dsTWCiBLR4TypjkPmld36p4qN8/bKyIrAdl7h/Y8
CyIRcs3ayBwKl432kBQ54SlGmD5LqaFXe1OJPduYdFzwu+dfLik0PxCOxO22qU18
eFL/EuBjvoTcgJ5CaVQSaBrIhdNwVICmtGG8MvRjd7or5HP9GupcHfEfgjqz4KuF
/wj3pf94vnG5FAgIY+EhLrJmojiJrwHRtEXzAf/8NzaYzLdjrm3sQN4Ky1zUmQI3
tmEEJiCxxjDqMU2nsL4SZf9Zl/43ZVBXsh76KQHPkJ0Gz6uwBbcawbacJaXKz0tC
zKdamqKo4NVX3WIokVQj19oK2P3//9IaIiGyh6AFPwZTq2obplwWtqhziZgYD1cd
H/aboHDbWCes+roh3UTGA4Yp3DA4U0J3CkCh5Zs1xkhp7TmLnyrDytdRLsDFiIPr
vHQ3g75KvmddNapFNRSQp7Xfznjm4uyGx9R9BgsN6Zpk7M2cqnqig5T10bmv0Fdj
1T4LrZFD5uCRnyrv9pXIgVl6qz0lsg6B7l8J7d1NtDmSSRZ0xxRIrvpcHPw196nu
AO26TGINgKkcqAJGLgh2qdMP8SjCSvoh2wkYvYe03DZ1qCFTIXfiWHiLsKNdkynS
lzNmOveRwXYYpN7rC186lQGrKTTxvG5TNhlVmwWajFGUiXtCFfJqwjW3N5y+bZpO
QhxM4ee7Q1yT/8upbfy7PAI7WYwKK+ReOg6egnCd+xRRRE1wW5sDq7EwjjNPq494
e/IhiZRsZvcXW/iVM3RRCuLTvVLhWuDI81jftSxLCoR82IFfvPHPCt0ifR4ULLXS
IutAV7VvCgVp1Px49ahbG8Q/3VgiHQ8ocObATkWtn3fTT40UraqeIfnc7kPUD7l2
KNHri25fLY6abJFB4IV3XnkLGOrllspLnfFybTNVBqs4Fh2UmtdhuATF3TBQJ0Og
P0D/YIVhsYCcvsoLz+nRo9fPd1/40CTWu0+HIsbGaX+KExkUUUAMjJdwh12NF++C
56pNwiDWcG4ILpAAyxyHEqb/EdRETFYDakd5hj3bLrDRD5OqW1ZPmC2Zzry5PvjQ
ORfD0OpbtLNmus1YBe/R5KWn9jJgqIodx4gFA/Z+uLqgohC9k9elKEIYJKfJSqZG
l8KQZ1n4heGQp90iUTyCBdpO8lGJAcuRT4z/evwpF1MvAS/qOsali+G1fd4c2p1w
9YbEZdASvS6yb4ZR2LLof0gELdvfN3o4eGbckmCEUJIIwpH2UPmckg2YU00HV3kp
lJ2/VYaeEdGI1QUHlSDpYeQ4E6R0hO7JN9rgzCzTz20wl+ZfOUtm8eC4+PP+bI5H
c+Ex6dTY5wlArA5XM12KDWGIff4So7KxF6PYz+8B9UaCBzxA/BvEfNrF6q1mm6F8
DTZwXRsDxFYP4YdtunJ8f5w5G3ymkbY+82V9oo1eUnxMZ/eir/4MlxiAgUvBuZ0X
+TFuiw2FpC9aHGvzSc+ZC0FtSwiWvtgDpaOqo/cwSE/0QBBb1mkCZyZPjUDvLxpv
ML8dLyIedhb2ROuTWhAkiJ69tO17wbPWn9THBBmURmd8/9tiC9E+ZAQ1d97Phs1P
VlOpsrGirLox7GvOs9v1+g1EBbToEkpAKorA+z0aOsxr//px1Q+Ysomtr8BwXGWx
Bzu6Fcy5Urn0v4r3OxAb2DNlTeyWo6qH9ZH8ElH4vNVyg+0oJv1j7H8oG8v5o9RM
X4dYPxeagx/RwxtZbnEOPGkSUTSNgQFpoZUIf+lJxl4AlsUbjfJDZ8NJc5vjubGG
el7JnZYErm6hd3gyfQaWDuuQeocSAfGvFs35ZCFlDUFHDja1XCY8dInuRehNpHG+
NNrZiotxmndIUpNNUIiuMMXU0E/KK+7QzWq+2E1XpdWzbzU3pBaavQM7Wk6vpktE
PbX1E1OPZhVg15H/vAJJCXUhFDu2T61VWLSNEB38CbbRn05m7b4Y++FCOYfUrAmi
DRf+P8JFUBKHEDapoKHMRqWZVb3nHL8xku0zrPfL6dKx5UGxsilSD2fLt9/Zbphb
OrLKLGF9QX6R1o3nEPUF34DqG2/c7qb04yWVjYwdyy2Vy8Asc5NczonG0IDsON0H
yxSbg3j/CEM+DueJ3Rl4KhoGqneiTUZxVJpj5xZqXxdb6lHJCrAkLw97lT4a9esj
Lm4GxgJ9CcU9gGfueRVHPfYBv58USnwb21fKfPjXubeXVaGUSTmBXnqeZC4FAOzL
lVV4+/ioZ+7XThXr1wSV9RDwYp0soeWhKDqa7iQLjaEGA1C1/AicdRo8pBKSRIYi
0gAUq2kh3aMLZncgKiM4eC2PNJ3RrdopuVlzzBVsokDa9gUSZsR6a1tsHlZP0rT9
Xsg8NrwtRxPBD+7Lzko6Km4xbBQLID3B5aOGLq4ogQbDgm8lMfcIOYI/bE1SEegc
bEB1h9RNatq6pLoE1zW4B70tXYaFU0t6gjq/60agu5JZbqU/+/xO1jUjq6I6tIgD
z2MoGAWK7ImoRwrk5tBdEoYtbCdM1+TBVvX3MHyHgYHYscJDAa2g55lk8qyOKWia
VV+K8L8mcCt/elCyJ8hLnuBAOkl9pBnbpwl1o/1secKIUbyJf7lQD2RNa7jw9ZHW
GZP+VmVkEF28Au5TL4U0v+c3k3aEOxD5xM4avzt4TJ1WstWsAPg2+MEIRenPIymf
JB1P9JdQ3/LapOkiYVOr0+FSHYyjx27cb526dL7RYbBL6nZOMm3zvJnKgVoSc72p
ZL628I3hWsgQ72xj5wbyC8iVOiuQbKMgV3hEKFbpzqDyKOcTnfZyEq7JkpNvzZOI
13+ErYnnKjd93SVUtZfFE7jImt9UP/niZ8vGF9+JgTnfgeiUIYxbi/owHmPM7HrO
SVS/XwLBydPlALhMUxJQoRqmG24hPfpTwebZr557zRHM3Tiyo8nt2aTc8Fhkg20C
EldZrLGpSUx6AeUMBMxiDJYOf/vJFxOOIFAADbTXAMiwx5v+ssa1AT5iRDgRuX+y
7U3ClkaQ2gujWUphddT6JfPf0KX/m3aqUPyuLV4xM3fY+aWlb+s92cYDbDxoGzBd
i1y0lOiey9xPlzg6LDJTBIXX4nrVAEh+vO/XmEvHn27HUVWiPLjTzAO2zlEkgrWG
DJIM/g6t+prSmOproEnk+HgRDdZw1eJAfYHtEoTq+JGkbLPZqQDQf5e2ntHWiKKA
oX6w69etLWORlCFtiOHahjf4H3xTXjvbOJx8OMr+wmmz+CW5x7eJbPOze/npWxKU
G/vrhquNDWsr1YNKfTactmWiQbtdw6mfvq5pAQDmX91wxGijjE/if4EKhhUcv+TX
wXoNOydbhLQ//73lkh70Y0LkkW7oPN8tL/FGDQyzWA+TPu+fLsMwLFGg681MhOEz
HP0pkbYC/wwpRJ20eh10Pl6Z2kIDpFO+m37RXRWSJjxjyk0525ViXKy/kwiPzhje
aNK01N4preMtArpcOxqfakW7F3lxQ9ZTCS0U8PsQNPXFxy8lGFSp8QK0NsUe8+D+
iL3aiuKZF9k5qUW22s9BF33umXoSwbpAEe1A2v/3emFqCI6eyebf+tzjE8Z4pqXz
R+3+B1O4tKnWpc8E6wCrS3S70759QwDX8/UBpsD7AY656aXTC45vLCxDoZU9J53W
s8VXUYEJV/su7lHBimwO3CBtIsfkcYEAq65A2YZE77anj2CS4x19j4MCzwt1naUZ
7SS/as5MCKb14fybsu2X/arSNHlOWaOUmeBWutmErWYaAaY1fRl1F+ddKEFbTiQF
1WSEEhciVMaX4E7QAH1hrgPizILYMczbZ8G/t8ftrvyjfJZRxt5nQ/d1mc0smohU
+WGdNPkZs08u5ST7DOcpytvNvz9eqXFhs123+HNyKg/ecvI1Gpzp+VD+qlU84J3P
U+qLK32nU2iWPKPCAccJ6Xn0ShLdjrBX9vHN74A8khqsvXa/dOjLCxFDij1jk4W8
/Yi0tcQ3nEkUdGBweUgOjqtzSZuVvNIl5cCikVxuCVDNI7lJPtEPLX+YUVJ5Rp66
1SY1qRzThLCmJGktfyWoXNnJpvFuZAtH4t7+iWJa8N527LYRn6gDNIwqT3vjndPm
dhg742DJEfoM971674bqAiNIaUPL25DfmUP8pA1+1UN3C7rR1TZsG9/bkuXHwK83
rwmYrU/ZE8hlwvwm7sDqLIg/WZtjPhkmLSOGTM4+HnlA4WZA79f0uHNrI/WLsPXX
7LHH3gkMOxgKp3GsOCPOsBEgSBkAWXVafIHWS8+/HEJ3cgjLmgxSNIX5zHwxeqG0
Wu5OyTKvqGLHkOSuql4TvYVfjZVW5svt6yl9N6aEHxpS5dxi6DIxgvxvKKQPVG/W
6/WrUKTDZDs7hq281W8oOMk/LAzSZ0gyHvRBNlXvb5PELmFyXVlpkJYrSVe1iLVe
jTicyVVir2G9Ak6SuqRaE6YkEcbGiKEAEcn7kMbvLkt9Frp5UOo5xebM73Ybspqt
ONjHoo8oy2GdkJVjsKc+zVzcUgJAiFuD/bn2nC96GC2+KhSooHuThDAzr7FZVvou
bduyDLDO/CX/7Th1YpUgSFW4jIdiXBmVO60DEwrXsdgSj7JvOS+5hIZ6F+GJ9tqo
yCgvZ9HuonaxKuOOOVbqobfbdvplM93zEmyBP1OpLl8LpiEY1pmOYsf6/RUq1jmk
fRdldoSWpbfk0xwwpZPXNiZdrbBFR5SD5OrjqGU27TZKah6BOgcUK7ODB5CWXkEs
HVGrSq2M5cZ2vizgfRoVnLPcUhoMpCcfc87R1wiO7Sl0ILck317UrpRPqLnShLUV
8s8b5yaFUGbYthEfdSaIvk2tGPEj1gy1yAtt/2owIWlLO/m6KG6KK4/m+mZk+KsJ
44RJ/Q13yRo57blVfk28+bbHwE3Jiedzx9DFs45+BCIvSCVi1Q7Ss4rbsIWQl9h1
0PYHrZ4z/LOPoouQqeFPRSMocGyezssimLm3QB8pc8rE5gYdfQ3nDygCNlklXvh9
kTaP+DnSXDOmBFxe/n5pAou3d/GeAQdG62G1JQpu+lt547Hjfie6iAo1dawB0Q3l
APdO9s3bKOCFsaeiI4LAwzskEHbxz95EonhvKPmFHBfEfpN9MffhkAS9nxn9r2R0
kabd4BJlXzeiEq4mCxFj4OzHVelpIzI+/qGRaVg1pKneE8MGzqeqEfTKpCZknhtY
DXHdFKyqj2MOuakZlWVaivl4TuefDRdhw2t13ZRNcDFy5hCKzuQ9Qlynk1PzbUJY
MzyCXYztpzUw71pCij557r3mK8k6u10G17IvfWEm4nL50x/lN+Royc4rOTBBC4vD
iHvkEJggNowq/v+z9wjarAoIQ2aoS4wB+/megn91Y5iUKLif5TjsvSejJuFb8ef0
jic2XtVrofXjsClt94EsmGTHwmiN8cB3Na9VChfOiPw8YAvnrPoGqpYx/7ptW27S
Ua/+Ud1ddC2Zf7vPd3DADTeoA52UW5X/r4OIUFyFcP4B4qZmNuLbhWlxO9pA/ztc
sr6mJuRmMZzSS5Qkhga516Hp02vsvlHcf+iDE02RdeU90SWv9utj6xdo/5sUDnnT
Xh8SkMbrhrfO2XvSKWa9Qkfdf2ei4ZPYgIRQF9zbLIuHuOgDoXSnqS77faSlm8DG
gP0svtnIkgArE6FD0emfn2cUDCcCiRRcrS+dTE4mPtcw7SxW2k8qOPu3vADwppOI
c/fFtwLXlRnCrF1A6u+IHeanCV/NU72pWZsq6lAeUvPKxT7mwiQF19C074rVWOIp
7+1D1hwbBT4fjnjSd/T1kS3CjpWYUQzT32q2WzKLOW5LOe2asFx85tBx1CCsovMn
ak6gQuZB43V/w4goxPlaDu7hJAklhpMkAxXzHQrhBiimzyudQHn9ndzU9U69FgLE
/BCFH7fhfJeFnZEfl3J5yxcciQ2ceboLG+lYyC2xw3IPafBdq260D2kNWINMUSXc
ehzsmzom3VKf4o6oujT4fiZVMxrSbFJQh9kT6Tr5iqljC0ieVZT5boPKDL1eiH0Y
etq6zxmdDiEdmJxGiSxr36ciEbg2UjJTwKtnqEiF/pfcfCnPJ35qBImrRr0Kw7NF
oSn/i78VcDMtD6lYauiSRdLCDNixTgfPxBOCjE/+pmHRDfRzzdCyHRz+UkyOJgnz
PBYRQJsePdorIQCpxf/1YY9s+/XDNAtFtcZ4G0ezxrgHx+11ZQ4DwjlwvwnmTxHh
XLKEprfJpEoiB90Ousgr7iojYIGs3x5rP0dwtpE1q7XWIvGuKmHWoL6QZEZ1vC41
7M/NwSIL25qe8wo0B6fPudDGu3Fi7G1pAkawDp5DbB6KIVdUSkq3/wqqH7xyYdR4
P4L1b+Au4vwtlA3Myw6SYI06enUiDWDORcVipOHzXY5p1VOc4g+U5ZNdWSjsVPXT
NuVLQkm3URZd7gif/TANYAZw/nXQswUy08KjC55pms6LiWb399YbYByi39yyFr/p
PhMqorKSqs8ZQbs2sGrmcih71EtZWobNpIXV1iOihu/O5qbllkdVj+BfAFW3JRhg
+zSu0EiWm45fgEb2T4+v+5VpRgR63DvlZGVnoVTX8Hx/Vm9BjVge6rxlrzP4nL+V
u95NPdvIotILtIUjC/ASOaR6QTF7u5i4UJ7obCgs+/fuqLPa4XacGqIyvYsvxu8x
h3vwRcssiTZXvCKlkQl/2JJpIay7hnd6uS4AyZfbE1h/qjWXekUNQa5ULYPHg8U4
gNmfYjsTKAYqNEo8o7ZXtkAQ6et+4aqYgDVaxWrSvAujvt1HePkKg0mOZGHF5MQy
o5ihPd3CFGknx86NXK6jMf2FP+UEuSfMq7kfhKeIRn4BOSbV0bo3F8mcHolk3Tde
l1tW0H9JUWieJC+9Gdou+o99C2UdCDI2fMiBHBfKDMQ7mF2aPd7ONWeakPaoMSUx
PJQ3FXODoIMuXx2YFZeufXXzugvP4v9CS13a5kGPHeP6kOYsrjewQ/Hd0jAMz/Hi
InW4q2f6jLmVv0sOlt2QCLDNCE0FopETJoIVDADEfmH3TvthynP7GSa3JmtZZv6I
XYNMMqYTLhrV8nQ8AxjN1bBjv6WACh+kJj812lWPcEcnTUk8JjMUY/96J03FjIIt
H6w0rAHMI6iGm37UFWvaOjqx57DfAsBXGeh8JiPtST0w/vrKorExHbFMPXxFUFa2
D8/TuhUfv4z8AIGaSzw59sw2eOaUBCXtmk6Jqk9BbWgWJHNl5rDK9T9SqWjtllMo
I4NBVOXgDZvJqEGRUmxdtLTR9KQAlBB6oZUA0kc/zl0lgKZ5alZhjsKda2OABliz
MUQ8n1KuUksiauqeWz1qjSCDNuiPYlSyAZotqZvA0jOpKMmfGrr+0uMPBRUtTtWL
VeEBwmLwiK6kU0911wN2GqmYletS/dda7+DQFr8MyqUztM4o54CZ41dXGtHKg+Ij
Q1sR0k6X29sf29ZgWIbow1ze+dftqUVrkBntRoAjYcnJ/g8EbfVK7IRvUdBMDTlP
BY1BaxKOV+VIBFJsSRshgWNf/uwrTdyRtVu8uQ/gEyxrL/lx8UqPbrI57pEvXJh/
Fb+2f7qypsht6L6ttZfzmjqAdXXS7vC0ZHJdGydNKLs1WKnZqGElk8uSgGLI0MPA
EQqUmGoi5zpDRD0rEfRh+pF1P2etZjMz62D9zzH5Q98iNmW/t5ReqMlwezOgLJtt
17J+bPegy/dTCWHSNlV1IKSGjnlTcnhI6gAalgpBDb9PSQ4+5E1x0xg1TB2Aub1U
p5d8R3riRnBp98behSzBeuOokJWXijq/qjDZB18swANrF8L7ccb/7NzPoxw/3W6a
BKvUNIV7Hp4t5nz6hMK6tSrO6o0edzbsSDo5YQXJV3ZfM+aiSLTLYcKOmfSBuI8T
j/dmsCLe4oCp5DnB5PgIhuvKGD9ILsTA2UfkSuXBIDjBt1X7nwnnWQv7foDFUJPB
9A2dY8kJFWzAea8gRxP1XhXIVr1UlDnOKMSh6Vu2cyGjqbsid/k0txQP2LgPzZHD
ONVdx4x4Pstsnn+H6JmWRJSw2bq3PbdzQF5a02vdSTyOq/BViEE5fT+cEBhH1dzN
BbpFTK2NVAhPY3fZK1lsmJCSM6iDnWYnHpL4qC4aEfqnS0jLW48ViaOkfqAYecVb
ZNLeCnqgtaUaTljYHbP8WVOHbvrrbzucuL6hTmXpvpbzOhJCXZtkU0abU9G28YqN
jE8RlI5trI/vzRbqu3KOO/tG0TNRQJ6I1WHzdsPvR808RBOiQeC6re5uv/4uXxX6
xUxYPxSOKn8tErmpzKWgSr9E6YekA7WSmJsVQd7h1+H4Zf1nCXgyKd7p23s5k2Zf
B5YbykZefXx47ZiljVIUkLuXe4r5bk+0OrPil2Z6SGMya1/600C5d7al6KGwSjKR
SPIpUYU0yoA/3Vvbcbt3VXlPd8I5ufvFl/0MsA5s6VzWORNYQsQXk9mJ3FvPT57o
W6jh1KUE+8Ad0KxdaGBaO3hH19vla9eRltxEwPrLfATET/cJ8K88+pWS6k2zJJPh
a8r9J9XerDVe9DOILUMRHrUe+HSbuMa3Btw4ojpZPbdiodBObOKVkq7HIzBMmJqi
IhldfulM8nf3NM2ZbqnGtwlnBzjwT3Qg5OAn0+JxZ1n8qfewv0hmjlQb5J+Lnd6N
w4XODj7PHZ+G8GCWmvR9OqC1Zy/dSt9Ksu7pGij8kkf+afQm9J39QT5Q4jmdNaXF
E1NIwvEwrRG7/6eIdQb/fMKb0QzBkZryVcPBF5sgQmvgtCBkFPLQrTEuoxKb60i/
/MM5r3DiipcW2UuudVTYTRr6VYPOPvJFPpB+ux5IGARsCs7uAShCuV10llK2HyU5
u25q8iv/Gh66jwoUM9B4eHoS7mv8KpAYt5KTYfocTylxF8LnSDo0tY00EEtkZE0T
sdF4jf+Hx1weEaDbLIXm/TbAeGuc57AyDrJZD27huPfB/OgjsVfs7O8fY7tZNUjx
/HXJsVXOPKr+DlCHpiPvamygOATBfisyGDc4ZDsDKkfoRvI7QKAkkGTwugvXLnij
XVVzM1GxrcKVhIAOt5cdvhWDi2f4/VOzY2o4h79dc+AzGgFQqcepgQyT18nF2e9s
W/UAuB7SdNGoFUJK3wGmPwRRGhU3RPgbKptQ5yVnJKmrsVL/B53xJTq60Y6DDXVG
O0nJSwiM6Pw6yj3QVxpalcnJjKokOwJ40Fhk+K8ESGnTcD++MOaHTDuSVF+QvkGz
/90xqH0fi2656GgfXn+wD8rOp4M8/lf2DME9rWcWO0bWOM68FCD0+jIO6yKRy7+Q
F9YTi5dxxV7+Pk1N9ITZ7k1ex9Q83DAdKZcex5cl8fLFqr/DSDexR4NK53BCeq8j
6K9UNz6nI3uev4BmQPjJtNgzM/n2YWs4Tz4+No44ipSuRsUiyJ6iffWWscWj/8Zi
LHLfMtWcbO/ZYOrU5dlbYj1fKuRuIRs+0yR2TXq1JO7bvRIJai2a0gQ4xutJe1XS
gIhVaeVFODzDj6Sp+MH/zgJ7tP2BbaEtbMShc7RpCv/8O0DOnl7jTOzd7G/1HjeN
xdZMZBxUl7S6C4y0+CwKijvZEnh3a+45aE2hPaigl3mSyuvu8P8Bj/qlbQPtmB3V
redg7zeLGuO7anOELM5/Hg33jjoVlx0UN8C7UYvf4qSHiPZbncM5zivd+VYsMe23
A1YNfYfw+uUlP+Rwb1A2Z2tCZiLouUQmvk5cav8yok8u9EwjZBYNvOLGFscPXo3q
XMpoGmpYC4NrExkcLC6pO+qcpa8iimuayGkm3Au5dZgGFPoqq1AUrNORm4Tu//d9
k3KzcO6nGvYkiUc1IF01AJVgECNqMidh+40dKqMxcroA628ngxmZkwixkRNFZXnA
3KYTZufxqGrPSJiODROje9eCeHztn8rDZS3U2k8mN0WXhGB+yKu5mmod/W5Z85Ml
OpjlRUVP/2eUd57HAKmnR1aY0fqWafiCGosYtfABDw4HyKviPn4BA7nYoYcBrBzB
LpsHVsiKlzdCtICAEBa8k3A8gD7Ug4GoCdl5YrzmmSqS1n4AY0Wb0ZTmWYnGyoBt
XtNGow+uLJB2GG8t/EVe04evuqaGZCZc56CWeiME77uqLyPVSYBdAQanZSERKldx
uYvV8kdepMoCBhxROETjr43jar5QWn+48SAHbgaaP/x2XhMdwY9AN/Pbh8fYZzA/
sOgoYnWjQR/x0gVfjMDOs2NfZx8ujIRlqZVWfTq+1LpfN5aCOSBgHo/jad5cukrM
UpiXca/QvB+/izqfkqI3w6io94LTvnXA0I94GqgK5G7S+DUl1+dlFdOJKzsEdHig
7b1rPyGpnttBTtRobeakDXMD/6YtHceG+ZSsy9qwiuKtKD3yQoBa+N0hphEmJSTY
B9/7Aiu3e4+rkpNztNTPWcgd/hDzylKJlTneDiyjDqUvuF1IegKoN9GKgdfI4k8S
cTjPP8ljuedzjGT7U397Yc1EctLxygczKZTSHHUvjh6EwrCaGLqgsKbu4hLmsgG6
oqRNxeCenz10g4CTj4flU/fE3DMVbdtaoLdpKJzfI2aqq5pgaToXQrGCG3zFkra6
ND7Wce3ZIxnBTGonS5stFollcEnJU73v7EeqFcYNY8kADR6VWBanIsuDUSNiW841
AqT+OaztjvUMqi0TxLxbfKn4+1KLoocKLA4dBy/UWgW6HL/YLWB6FcVkyohp7OT6
A0RCBgRbedCf2ADvWHwrQYYr492udtC5u5vQUqupu4jtIi2UTGAZ5U1M9U+FeY2a
h31SZFgoHweXfO4RAYZqS1KWWzySusVr9gmFcBIYa9WtOngBcx6PCrNKwEICcrsy
4ptD5bFHtYG8i588h3ik8+3jFXhEDml+nq9xqYQjyem8BDNI3U2SNYgfRdzidfjC
5jvL9E4Tg89krmbICTSjcVHztCPhGTBnTM+wU4dZfr/1hxk3VU6gcxO97fQA7K2C
CGp80ulpCYfp0tbm0VMJ/N110z+necjNJxOI0xRHng0/RFWeoH24X2HyDqshF7g8
PzTDLuFC5bdhqADDOSWrtcyV2pj0dGUBxp0KQseNHvT2kJi56UH5H/5sdG1hFuXf
CTpI3iKwRuvOIqU1fSfznly73WvXbvJmjiO8QIKS42eQjPLYMlO0qbQ+GbbaKy12
U05b5BtN2phg/dWUD8TEl506jpP+1bgIci7wsxh+rurjrm9WSsr3TOKkWDKrsgsw
2utuOK/B8+4FwQA8rlQzwtyiAAq46FLvlKdNjxZOCdDa6f0RlEwWM7n5CRCJx/sm
oGjohonf4QzT84ysQCh3kqLP8nTqFkFqDAxaVSP+yD7I187sMIrIcj47STBop4/N
QdFu2CV+lzm74lwaCTEBK4byU2xxUJPj+s5MIZTM3ZzbRSQVs2R47a590oxmWZSg
yuJ+DjOn+cEWq6WLCHS0Wwyd4CQSz66axIoioYRZkE7cWoOGSfsmKzzScfOqvUkD
NpypNX/FIbfZDm/N2gXmQuqdC5V4Ba2cKoEQGAxFMbCiVAmcsrauxKAyb61OC5ZO
LXRogN9povJNsYgC0O6641knmGwutFCr6xEvoJqH4qTPdFVvf5N0Ru9vwoQ1bRiO
d6mSPb9Y5dcuLKL4EZZFag6pa68YDGopKr/zL5zZjvtDC9Ewe3ibul//KTjL3N8K
uDEFAgGNzk1IRriaD2KgtU3LPC/OD0QpIt9VERvXvv7Ykk+VmNofXmqeM1mhVJq+
MNSwPySQRDVIVnWqMuPlrLiBxL1IwfW+NrkiGLCO0JbUAxPWttGYN4HxG0pPHRZM
YQjDIg6LLdneGlPjI4BNWempXs1l3kMmjpcnbZIQ5o0qsgOtuiPILrZH/pPbe7Wn
eaMFnBkEyLzFB2M9uAQGkedu4fdtUBMJr8FqJ2cD+nMpDnJvJq4Mm2cHtHn5fQ+B
xjzrh5kZztQMoIRVm6hidoIg6goAhTSJkMvWPMfKbtAR4CLG5EhMGFCAanqkcAgB
sFIVWPG0GCypJJF91u+30kIlcUhOnzHOzYUdtgbPSOxfCkaoRqDyActiK9Lzfh7w
CSa+Q8z3936vQ5f2DwOBm8zIWAXytZMd5q5/Ob5c1RRrLlcjOBXFgh6tAxNBR2Ab
e9K/1yuVWOXU+ITw0bjAu8vFiI13SsmTPWr55vJY5Y5ftJJZBkvSh+tktpQSmN9K
oXjlyO39nXGGDJ5gf0mL7J/QaZhREJ7gNFPi7ALTpCY/uixFnlN0S58WNG7IoR2l
YvoGquDtEScWeCJLv6n5P81I5l9DRsGdRJ0Ttg8JkDOKX5KCIj6AUgAf/M2ds+N4
uzdexjbrvgKb5vXkUGf6pDx2g734vC8Vlbk7kWEVnTa/DAQzRFeYdwrfDb4ST4Wp
b/mWm9lvJDAaq94901Az2GhMmm6mYHw3l6g4Itoe6/VxKu+zP4VidGDDYDswQfbn
C7wp+T0b+FyJ4i3qOoUzq8BN1rU7HMXJDLVMXtPsu1dq5gEYjcqRT7aBKwzTNaTm
IX64/RZzgI8YsGsSaH7UVr2pf5Bl6XoKhWqgOeo8Euo4smJrjroqm+QgyzFemvVi
lS72s0lxLAkk/3lZQckO0OJyhvmGUe7sYSJcjTO8hFFhjssknoGjXHdCAD1q4hdp
0pSr2wJiDGSsHhL6HsDAThdf9m3k9nKCoPSRNERf5egOwStMXW+sE/Pu16bSG+36
1ug02SLJAq9Ngw7VXY0VCWO87YvSk5QmqlVGoFmmdB1qDSW9S5iu9x6NxGyWrGvH
EhLXbl6Ow66b2UHuAdICJ56njCNgv/9JouykK+DzIBEzijzHqYPkqVvjXCjySQZl
FodoQNtckAqXzth3hyFvfYn89KDc58vRPjUbTITHWaQz4tipWQikiew9rx6un/1h
6Nx5szeJQnpcE1MJO7DahKeMem5UI3c4RCLzUROGkoUJACitZqze0ewjC18U+31/
VDX+3l0D7hUsUziiL9Hi2cBfS3Ha4j1iatoi8yKFG9REOslt5jufnYcDBX+dxwk5
/whyFaH2MSVAOgnhYGznT4Lz4BZPYGQuQ8NOaiTzrs2EOkwGh4pxoabNNpWtWSlQ
AJ11IkeLCwHaUX1r4FhLnPySlxc2F+qI6zvcE0pdbQo4MbfVmvuFTD1hnW7K0mL0
V3booSCkAjICuiYAt6RJdXsdtJTC2UyOgIZkS+IYskgJlx/MCGdI7TElJlZjtIhb
OwwPi+c5Ru2w6SILFV0aQh9TX9+6aXKzSxDczrHSqt33dCMs/zq+oOLBFLZWvevJ
4bhrMfJCREwZ4dIW9kKlFLFSRKWYozCtRLv/o3T2QraxO7LduPytNRERvEjuIJ5S
yQj4WSR8XwMn5shXDJ2+u109wo1upKUvEaYg6Q5ch61Fxu2GopXRG55fYwc4y1hT
BOtOka2Y1e3cDwCWTw5VNJtNfXncscdAb9vj49xZCCeMmLcIOatz5T8/kwOErbKe
L+LkNgHQdOSCiOqAScSsjRXqPwzMfqgPQ8O/u4z6VR6kq4MiV4YYmOmL3V0FLwEn
Sut7NwyE3aXe67IxBnbQnr2VP66L5pCUaN1mEo0lT2Z4nNPcef27XIRPMCPY0cce
oiMUOoa5SAwuyocGksReoP6eybdKbarYWQb+wQI4Xv/PvHmgE900Qh8d7A/6104N
M7ozvsBhHb3U/xsjEjpanYZIjOIce4auc5sy9Hy9L+z7KelaMALglG3d8mr5Y6iE
nkeR/OSt5cQq0b4K7GpmrVU41eb9AconO/4SiVsFnG4eyJlQbDw4nFDpyGqL7K+p
LlpRQEyGrR3aoy8yDK7ATrKwYrMBN9Fl4xikAOPQPrv6qfXxnjVgo20v2wTGrEm8
UOX2ThTE77ZBPHOYzNiNZFG+nbGY9/+wyEhKaDuqmCpBy7TIwmVxnQtq1PnhPdHX
4geCPCErzIBnUxwjFO0D1YUxPKdGp1DkIV5z3Q5MnsuBmlhy6gZcgM1Tol0a79lq
HktKqc2HI/g3Gj4YXCF6fkdP5M3hQ8pwcvNj2uk3P0lkIXBhTSL/p+0Ljtstm4c4
ZLKocGDWrTSDstPA5KRLlCPNBLR0S1YdqYmgaiD2POfxVlAZQLIaoZueuLoP4/z1
tm1h47BFTLvdDKVpWIKHutdZH1oUqn/Opa9m2yatQL8SL+HoeW9o802dt3+zhpb+
IWLMKShZm3g+8nu6jcyrwj8EPYVyj8dW0mIpoNXDNm1XuoOPsgEbaSWCoXFXaiYF
Av+qI1JMH89Qea9eW273j+2OsKUwVGPxRwsDn+RGoQ74zjvduO24NKCJVMd50s1k
ZXH9pzRRaunuu3uRPHkBwHD8mjj/VX3wSw6V2+2NDb34Ub4ilC76/6WlKWwtJJFy
kjhQuF3PMYRtxVo3OWBIzkZfy7WoJVCS/MwhLJMtgaZ8tzipk25+PUq+KPay9YOt
eRNRAE/3Sk7ocwGrgJhuGurLWo6/Tf53HZ4TwdkZQm9konGj4RH+EodqfL31W7L1
5oerWN1bIwO8ev0uAnhPXcRNKfzNq0sfPK9ZqdXHWOWAi926MiDTBvXEQrllcO/6
HogVLZqP7zqMfqc4eStyzhEzFldJdS08PqqrgwFvrffCUKGRNmN7mJCcJQTOK05V
rAyIVrvvfYR5geTxPznbYy/kL9a/9DSulxM6A1VznF5xb8fM6586nk9zfX5IPPSQ
Mn1vvDOxchwH6J0lQQ8jcPvz9cmQ6YfbsZs4bd1xdiAmYaOGIpWjqiU56NEZCZVB
W7JEVDkcinMLVpUzDhSkbM7/tp+c98dolCZIaZqC1YKYY1qqMy0FWjAZpl83ugvz
OO6eEtL4YEpXOYGZQJO241OeyUQ1dbtWdZAflhtdIZgmKp4CD8IBsJ6hmpsMptuQ
r7jjCozZTUrhxXwPK8Cj8DjM5oguqljejCpYdMJzlhnnoTOAoVU5AYLaseee9IPl
YG/pljO53SANppB6CqXlyl8+tGFmDLEBDA4NkVddO/q6i5yG1KKVTOKUgEwmz5Wn
UlTyPoPGOBBgN8WjFv4gs18y6m+oZ636BgyeidCb2kUQ7cWlYjlMObiuDqN+ov1i
INcpfuE36Yfp3xQG2WpjGqi7vGc6AdLo3qXiZf4+dNCY1nbnc05lErIxHOx1TKMa
zjo45iHH3rMZDMzWiHePBshUwE9HIZDqbfDNPLHnBuNL/XKiFl3+xB+H9LCBqS1e
lJcrQAW/dAKgGDn5muX/svuRsu9NPn1wJTKCcoNS/oLYse5wA1+ffHitJl4/yXcG
rGbUrLPejS8wgU/7F+5vWBEwvFi/4TKW1AzpaJBEP/LhI6xdw94gSfsll3XE5HRd
WyfLxSGEgqGZxyraCEX8Uz2CeC6Lh17c7RGyzbyv7EkAKBu+ke13zNhDfe2cpQGm
2FKn9Ab7WPC82kfrnk1igYGaccb6O6ZFFBuW8bmNDhpPihjlYJdsDQr+yGwVT6Qv
848FNLI9oPkUMs1yxP/uhc1/8DSyBKlzgI8MH1EmkhPE1EpgDz/SxCwnAsKn2QHs
RKjBi/3OGIlL3JHHdKQFT0U6Dc41ClEPY42YLMswrOG6QxJG1n6yxk8rNrPK3aKg
Mf1ETq39M2oUgQftvx1o6v77MMGVZsGfkTSR9oQ+BOC1Mo13o8j/rQoW9P8GFpND
/cAX+YF9vRgjabPa/l9GAkf2dd8cwSFVdBpDS7lmfvYE8H1ttmvZoPcqikFg3z1B
Op3HI3Uyjod7AkOwflUa6B3DHcWemXaY786ydiGHyqkUfTdOt1nufG6n672y89oo
FCgYIUVRvPUzr5tOaDM+FLACwB91kz6dnN3Xu7gjvGoAD5ASgdh+z4OMrgGUSmrN
NFEttLAKCpgdiJ36bYkisqqoVBE0omAu/vjGwQ9O511OPlyCBAeOFRdUdC/o5Nbg
P8E6lBwgGAoGIIWRopAivI65k4LEQfiF02shaS0orD1+HgDt6YfEf14RzEsaDZ6P
cWA2TyVTNKKN5OaYyCeXRSkSkhHFMdJgm1VqmkxY7Vw2LbzGpVhEOdR24W0WJ2DI
YtdOJX/1/p3e3AeOMOiK6ku/qYwllUtD4yRTYN6aeb0vs8EAt1NUfJkW94IXQ7Y/
NGVCs7SU2qwXDfew/oHTi0ltn8/E9ODrGGo3s5985qsqCvVswNUFNg+S5X8J6fIO
JWOkpGKBVwmDDVi5Wep0TMjK36UzGJ5Yqzov4SMYfc6Ai3iWL/e7Axxd4/hzPkR2
7mqN9k7gpxtSYp6sIq9cMWEdOYzL9a62C69G7y/QJRlbNgIJG4/1HjdJLFzcvWVR
ZTote+vYvLGJRJyJGKaPQxtHUtNxzVkl7AqA6o6AHV5Wv6BebVKhwso9ds8cqJ8j
PuukPZe3RANTUyjwqiDQjYKKdA+022iFzUhZdXgusYy6FN/kJ9iMfW3nrYCYtGKD
E7An1Tmx38+Tlzvo0lsXmMe2xSs6jfocULtiAJVrbGQfvAbwcTPRJxxTbIk3+brk
YUd8n0lW4zF7S6JKrIOKRch1G8h0X1XJGfTE15gVMvz3nQ0UBofm9edbhWXx7oC6
M1m6n0coJaCSjGzIMs38ANiuJDkl7UiaG8NPrDN79RxlR+KvPjgjNYpRDL0ypvzI
vemdMC7rIiY9P4L9QKk3aX6Knci92tZjyqTr59hXjGqXsjQ15uCkhlrNhXuGjMES
qbO9dzGRiCxe3AmJCBiaEFFBP4Z2OIcoh/lDTsuAHwN7OqLoTh0x1TVVe6p+72qw
rjKZd3p+0PLv9a5pNfZ1oj4zWCydfhVKmPhMxha9E4cLO01/wvJb5iBGf9gYfSkf
XmymFBZAx8mJ0SVvNrEsAvTPuOuMZKfU/t4GGqVU/T/OIYYWr3KbGflHofzAt3tr
IJ/uGFA4pOOEadHL9Asltr2p7ZJamMd2Z3a6mtnfqnOzL9rRIKotnpJ8hinQPmHF
EhvSEo574xg7zGd2gx6ubtDOFbcC2uyxns8VJekTW/p29+8wCYLdFHfSUKQj4Kly
OhbthH0Nv5L1cECXHFqKJTxfzPZY5IyrBp57PneTkls5P6+NwqSiLuH/dppo2tIr
dyYQgCkxOMqgAjsOMjVxOoGBvRvYh6wrlyZyKMNtjB6N55I6y3xLFv8B6ghyNYWb
xI4MwXff2zb9lWQTeuli4+cGDE34JqZytNEwxrjukNUqFwjEJ0L0Mm5rqXZYaPjM
1t6PObYJlimXb+d6pFKZjIQAjBvbYEV6rgwLUA6gi9oISZfE/WTHmJ+tp5Etdetv
sWeLPtajntkAu05zS0LPF3hr49BGlvEaK4pPSW108fLq6F6pBDMdiMrMhkm0oz8W
t47PgN3LjOR6FM6/DAcAW4pOnP2i3B8itQnrdd66lfM9dSZruS2QHt7+XMaGy9/A
`pragma protect end_protected
