// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Qv3emCGXVIF3b46NsaOpUk6X1D2pcFtkyOpTzDCFOidPA23Mfi0tggy0p9pQfGyB
dxHsGLiDccQupYJf3Ki7skJT2HpkQc4Y2YjuJpregBsT3IhL9ZlzXfqdtVnKZTDV
5cprW6Jkxz2qOXb8yPq4MWy2J8j5TYnBwD6Kyy0EvEQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7536)
TKqlSkzjirXhEudTBbS+Lh1d43ZIPX29zi9sqHlUNqOaoqMYnvqdPY0KBYgSoBCK
VXEEXbRn/VKOgx3OyrE+0l5FRwvoERvM41kfIvtO8vsboAt3yf2WVwOpBCeSMv9L
bBY7LnmbQEVh3FdIqGGuTurr2c3CbiGMZU1jkJdFuCuYe4C/uvJCx2tixouyoE6/
+5xEfHwUPgL9xt8sGm/gcHkUebQOUZ4xm1+eOAguaprB3OPvFs7bmhd9LEQ4xI/T
j9+TpcczhDXxIOuvd8UEyGYgIlfxUPcCThc+xqfx4QV07FhDQKj5rt8mHB/ZiAig
1oOrsApeIbk1Wg0Zvgf8hEwT+VyJZnUf9Q3qhVleNdMNMwrzU1yM/ABZt6ciAAln
gdvN4J7Bb5o9o61W0lsJn5QA034fjaqwg8vgDJDvwOzRFOqfqwV96vKSi2fsG+sj
0/kWB43l6S9NDmvgNEIS6OP5Rw0neZVnzEqspZRwin75gYsWz91ybVMyLHWwk7DV
kjWi2QLnsfAQ9sYyM+GL8tlQv1BcKpcsUpFUUE1t1K2a/48kpJaRHVaoAdl21ph7
YJALCQJ82zx1f503gmjej2b9nzo2M6uyAV4u0EuaMOL0GEW1DFwP1k3RCnRqq2/W
dDd0400nRTcofI3F1fK2gWSy5Ds3E0mnW03bxbKsQJNa3Ar8niaWZglOAPf+dzDL
cu8J0xTyarbqqZTbF07eoVEe8ghyN1v/ACpz+cpRrT1E21H4UwyvuX5CB+w8AsHt
0IdM8U6ptgxd3RXFWqMw7BkHALLDMMW2sv9reqU26e0iORGDi5lg4AdoEYCoJyqw
S2fPwksK+rFomkNcXyUXTmzNoubjtcIm/3LvzKivAJW+PTasaoayOcBhOQc44osB
JJXpnIsT2bXC1Rm5za5Oexpgpj6RlU4uA5opLw3pxlxw9BnO5/lOkshyPwe8r9Ac
eJ+UCbu29X7ccHOmvtSJznHOekF2raBaJo4j9muaqZcKUqi2DNDxBXz1HU4ALyqc
Ypvts5gziy5shSHcZ9KRXxSWHUjdmLuJljyDWYtU1b3Wntq0RrgMnP45nGS74cdQ
SmXjQUAYYOw42eUoFvGwxU0dx5+oMm+HBYqu4UmxCror7ni6wOh5NNJULdh4cfPK
0sVS0vTGE1eKCYMaDpwKPUqIXnQnQR9fIRJO7hh60/IZ0TU5O6aribBkkHv1hRZD
wtp5t+aVQtOoPbDKcTLQ8M7J3Q813Bp4mosbB6aMoji7CbDwEAm8JvRvJoiMmZgP
AWEeDlL3bSgH5kgzTVwoHTCncPm+LIfAyJFo0tca5uXCp/E3vLPeQOq3d3DSdtr8
mHGsuup2QZygCxlqGMUA6cg8Wz1NBI9NhtAIkFAV7qoC97pgioepBjnle4rKA6OP
kPntZsl+8SjKfQXWWQSAKNv26R0JwxN+J3Qom33MhYmw9PivSnH+j3f901+cshOp
EqEVhbGD5oJurAz58HVjs+0mMOllwwilhSrDHT6e3d2OqIucmNd6QZ7iEz89R0Oi
8BPGRY2siLSS/4MDhbPUxhrWMv8bBrQWgJsxmd0vGhMrtUsDU2F7u7cEeNerebvX
X9wWAwP1CkX1UcRWF0/fdQNIB+ox1+aEuEFY8KfkXJynM3GI2I0gDmoGxe3ANMtE
kGj+0xvCwPKP0s4o5nF7W5QnrIwl2XclmatVm/wb53I6tSmf8CsztuyQr2KclPo6
jueTScluvppAMZUpN5lyusNnWp0tHWak4hMl7TNf6bygWWEQB08WYITrZxbYL2nD
SDDve/XHy6E8X6DD2fLXXSQe+/tVevV9HVAl9jO1k9daBszvEds47Br6iuwr2931
8wTAmgc2j5HQbwsb/W0nTZk8k/SZxoPfNE7rodSbj8LFdIPMx98H7WM4f4XnHko2
fvZpcN8soSV5hx7StwL0v4zVIfTmWksS3fbN9fxypK8ZJt+jAc3ceVcSy2o1g53n
a9ZIFtUGy5hmS9vDRBHIuQyDqU425JybICbK5zs/vmyJ1+h19DQy7uBHji60K08P
rf33mqs4U5+4XG9Yhq4sTU5pfr1DYHUu2TsDXf6bOMxXimQE5LXftQIfDHfaUQBq
bFYMWp7lRylqL5M7ALmk9BabiLdxjt+/DQpanp0WvmivqfwOd2jnDAOK74Zrscqg
vhh7a25EiJE/XTJ3qOBqiPtwXtPA2octLMFzvI6LQqRcjKvCK+MUT0cdS9XJ0JUQ
duz3ExAvvJdD9HV5eJLsYKzDT4CSJA2j6S3UY4pV4VPXziv2nltxOZ4WJtYkkfdV
zvVO0RfAzi+EhFoZLVa9mGAqXzu2L+ADEWAHd5shC6oqAePDT04iKCY9QSssQWAG
LcNE6QM3wRV/RUTEM1xkIx7S8QnK7SS0iPJGX2d0UB7BYCP9n99BXbItrL2JzjPZ
GmpxDqXUUgvnryyeivPpPY3R/46hdmvVx724XDrmOIS4hlOcjdhIamhrjtkXCnXT
gS8SBgK1cUVkiXnDUl3v7VMfjkr7NCg0VoqV2CCw6GT5p8a9Vah4q0R2FZfB9lEN
V51Ew4wiXLD7t5UiC9gev8Ja2c39uJheTt0bdGyg8BmqOc8MxCBLaWIMP8E2bq2L
uqz9OPkRVGYrZIkKXteCClxs7Es0B63XLPaxKETAITJWha63EOYQfq0Rgq6ua69J
X0KjZD+fr0UwNWMjSW37vrhzE+bLjgLkI6bm5Q02+oIQ53XLYPrrPUZCuZkx/unJ
EfpVK1SOMeE9svuypnhXpFBrn5p5qfjnrJJfGvGqenweRNhJBKJC8tDOCAzSNBRb
CbWBHP/fpNMk3preLyIR9qNWC6J+lKptYV7Dh7mFSxoLUsKPG+1UUa389RM9Mkc2
7289h7qwAPUAJLbY319K7glHFQ9KmIfQ1ltU2+dkVzL28Vk+Pcq/GvRJRCLSVBTr
SJGHEzyzAGKgp6eNLZqj5n9qmfhvQWyeLzuIvlHUAL6/rx2BZMms7zklmquxFj35
DLnRpgtEJ93iRulxtL68E8F9HslFuYQ0TbdDvMYVHHt0dHrwr7DKQXFtm+vXP550
PkiN1h2t/pcWwDzX0R/NUBf65kMWy7UT78MG1LsvQmdFjtlVri/D+2Lyv71JWF2i
F6R4prDmL8pcJUtLh2YSuGDjDNb6TDFAr3bCBVphmoVoA7OVoOQh1Aiw7FpvWs03
Mb/JFsifJh1bi6kILqqRAAG5truACVWyRxLvUYl/WebvmuvZnxl8G5B01+RrV6Nr
dY/IzaOm/4CF8q+2eZkLUjs7G0zG00RlQsdsvCyRiLfL9e+KbqSPFVNR9hkI0NT5
dKlski6YByIaBC3PSHSoG5PxLofhykpuhHcNqrwhquQ0mKzrp9Wk4cbg1GjkZSW9
htdzZtVq23wOc8zm0NEesGYYOQ28QyMR7WZ3yV4C/hvu007xyMa+ywN+yJRfyqIs
3O67NfaTy+Mn1GIs2ywL8KNkH0iP7JzA2Miw9H1unQu7aCVJdYcOHrpKiCyF6m+x
xTzRAfFVZsgjZYUCF6848wc1gOVs0KGdaZ8sHsK1ffFFNmiv855uEEsSboNCULYc
y5iZlDYLUOcN0XAaA5o5dh+bgBR9HEL0P1TAD4HeF/wEScobffVDZsfqMOTTnWmc
1mZ9Hb/a6GekZFdCRZWdiLdAEjMnt4gyuWfyW5UW9qlxwx2KVZZToBBpsU2apZ6R
+O0hFvCmuLaOuqx4/TmRLYzd3s1jG//obgYieGdPvkKNEhpF7Dmnky9x0UZVMn6j
Prj5fLyivhNgNcjd5jbB2vjYYPeczAZMcUpr6Eo6ktUqWomqC+w8jbCgks/T7BhI
P04ihD20WEt4nrtQ0OTLlD+E055Ke3iiGMEF7HhaGYteTI1YulVLHjHS4kzkUfkb
PzVAPbz+TP7I9ktHmxsyKC+BlkCoh9EQ7jkECd64Ol4WfhGb3lJ+195rEp5yIUp1
BWLVgfToQ/S8TBTz90mTWc9G//nvr5RAbobpJ41l6PWGIPyKcFedkAA75Pkxhy2q
8Z6MfpEwUe5AD5Qtl9yx1orkW7gGjRinoaLz+jJS4ZoC6GjGrJkBdvQpmGS4t2tJ
yGw5afdSw4gLUOI5h1CdM6pXWQ1tdtL64SnzD/C9mhLviA1gZYqrbnr/X0Y3Dr0c
cNvnl4nWCPgfM7OFA8QH4xS9jOPvbyPnqzh4JMBfI7toFtHtXdczUsUEU40NXYDs
GfyUlKQIHDXpzdlH74fD3Vr31XMc7J/noUHtAoKgEVwbB0k4tNvJjorlhnOufLrO
iVBOSEaFNq5jolC5CTokXqclVMkQ782QmA2FjzrfqirEd0MXSRQDYXVwabEMNnZo
Axg6EV13uAzY3SSstORXg6B/exvizkBUYgj21F4q1CStTgcuH51E7lbxIsk3lP6p
fRYVGhITh01VX76Wo5DWWROnJZZA7PPUVweJjla7PhGttxnkDbxBTf0y0YgES61n
eJup+78wuQ6oCx8bH58vr3X+8nrMckBoC+DzOVfFJi2M6VGEU36nS4ztAP5Pii4e
YC1gst6kR00NYrVphJzRPKirQf2CnQcY9A7lO5gtj2IekkeVf+sKiRDnQe1bV05i
+atVl3ALp75va3cMWzBT8YhcliScCFJXVaFIzUYJy2EzPmAsvOvB2lZMamCuQZfD
1WoumckXxdb5rqgM5QPrfQ9O0kzy7c5qg/Fr1fkK7himLtn3PYTmdq1wSZSd3Mc5
FzOMN0AWOdhMne6xjAwnZTE9+/sUu+BZ/DTarn3/DJ18H9IqcghuqdEUsgGtuZ8F
+84jH4OBp6vEiaQjYBHXff4MK5OPxcSOebf3mrrDD2I6rVrjBkpiDVnE9D9Qabwe
jeoMcrbkbDdLbkVu3NpP2kt4kpMseRnMUsHwGsejt2WzcJhzbFsAUGIUfJ9nkNxw
8V4Os/yu0gM+BrZ/1FRQz/ftvWttfYyn1RRzPtByG3ybUeIH1yubQfxXIk8Ge/ZH
PF3RsMIP3vd1TIUKrt3FodSvwcqDIrTGNmD7xLCc5hhOdErR7jU7MSywaZcf0gdk
DaiLF7rw4hdlolO/hgRnjNMblxc2bW0MLYbPMUMz2XkBhS0/UERpj/LZGTZ3zRJb
KxsUBoWkvJQKg5KPv2uFXOh1YDgiw3DRGbroo+8J9DFtJJ3/qcbX9ZqJTJgDpTwz
oeV4vAey1NbwBP3U1ZI+94aNuE08UakcisVClhgDcn51xIVfu5gBNmqoK2UBa/Km
IRJqA+g4qEljfzB/5xvBv2g3NLWLDaNQRZTQgHqtHMkPnLceUitnDV/CZS0n6dVd
4MiyNwZWj75IYGdsxUN+0XD/dLh9NtSaqNUfhUN/H8HckITPEclhubGQrNlhah5S
UnLRdOUd3as6pYVEGdvQ6pQVJrj9dyrjzaoSjL+ignhwa8x0BiW6HGtoOnxgpL/1
w9Il8h0EplVddXw5ziMFQII2YmGM+mroJDYmOZ5hBWkUJ7K/EkXWYaGpuGizjrBn
VaYGV4zSyI6FpaQ2pZ7f+mU7PBUTE0RnJuxeaWX/HV8pZS7Ch9diVq/IRiqqPc/h
jgC5s/UiMXuCKlRHGWczj/EmUZpnzbEAZ3Y+joUIrLX5L1sGM3jyC0KdfsvWRR/W
qWGhbrbtzTXUxLDXvXCj70oy+k/NL+DBLtWtChQABCUocz6LO5cQGgsPIGUebHUA
y+TQlc+vt0mSECB/Q6g043YCxJRpotroBRMrYGNzTmnNVF74i4mFOSXmfxx0hUSb
JWo+5qjRJ6x7HMuROLoctjAaIGhtyuth4YWs2IW+z4im2QRqIYgFJoIJypqybQcH
Woxw7ttObNxesH7wcfeYuamApaZTDFvqVsyPv4Zeo4M3+HPW5AQVNCn3xN+q70D1
RdMsdGA15PO3rkMpSUruYD0o/iK+ZjVrHRFK1anipRz4Cz1An6ScDP6pBAjNutF5
fyql5ilj63fJkhs1ewreWzG8QurjSBew155I1UbU6ocP585R2A4G1oGSiaO+RmIb
vjzIiKS6+Vvh+U/wjXOHf6kpLgi/Az5OY52tEGNhphaA3CET+yLOtPxmALmifTF4
2riG/2LBI1HQrFdKOEspK6Z1rsEsWOiT8aOqUr/zr1fR6i9i7r+dFkSOSnNwGfRk
C1rIPfyXApdk0YtjBAC0yNab+5UToCuCzr11SYiVw3xK+kKjX8rLEMEFzhpfMmHs
S7L96LXie2Ey/kSygnZAXPYqylPRRjqZD8mhtpq52UB7SaQMnUGHwD0MCK8Bim/y
fFayyHd1XDcYHITrOMndvhNwnZW+JJlHAjV/CkWhRMQ4eE2LddxzhsWRs5nRqMtA
P5KA4CV/PyqFxhAOSKgplxCYQPh69okJjM6Qhtpi5xLf3PyzSUC+iU1Swbusy2T5
lxisYwzNOQINg3bMgT445/IeSDebYTzrRp9SnZjiuCzV0LSy1CTkUYWUEqxQMYKc
qONYW4wFOAg3IxVOhD2hqSrtX41l12GUDkh7E5jhthD1eWXDUB0/9pSHCS8ygLBJ
91qHFA5lgo+k0s1CS0rJKutttrLtM4h5F5wzWgeb5H98/FqWpmT7tazYkcU6V7fR
jvQ7xcws+7a+KCb7aOuRk6k3mL+AEfO/Ls4VvYaUw5r4iuMPQwHrmRv5ffAP2o4Z
+mmsL555I1FQCkCRasqbAVAiwLY8iVl78jXR8Et67tp6UDDzUCp62DjaESsi5m9A
h6hJouZZ3nVL8ru0oz80A/yQmA7H17RYqknkmE0Pa9inS19/cyxnsF/RZCl0uLDV
xtvU0blprw1MO9E9jAaZlMSn/RFzwH87WybwHLNfqts/kLkMU2e4j32snHXiB77X
IR5exYSz3woon9XBi7W7ZmhDzl/1937XVgs19VYjOqnW4Hq2hcLEGPkLhL1jd0gN
LCm3MNESisVoe1hnol+uginfqxcCrJeJZj/L/T9JpPHUcgvbUTkW7GG7OM8hsbrf
GfqZJmAmiz7+VRU9Bg3oGPeWFOUejjBh9fUnX3+VuV/Mk7JXdpL8ypUBR7qUpsTm
VPPlG5IHaD9Myu+n34/OPkaHghFXRfnTEQpV/pABz8AIDxu5lKH3+sG6jTZuVy35
S8JFJp1ovJ+GiEwTyD3wTA8tm+KaxiAk26fwzzt8gNVWc66Aa6m166NY3tv8OKj6
NOq1eDhEtHdTBxBqccrzWagP4eghslfjwzwhGs5s+EugU/EFjJQYvPkaz3N2CyfW
sPO6bvD7d8ts+KRb4WCSs6XEQqHAx9hngPIMrwpN1XWPRcClfzSoZa8zXDK847zp
pc6vnDb7IKrcKGhqc0irarYC84SsoeT/5ws/5hDpanY9BJalDu1GGMO52hkVgnDj
G5z7Gwm5UQF44Li93/JFX/4iTF6fLrTdTaaq3Ye5SQzb+vj47mOBYv1im1M8TKdw
inCmxaOTT+mju06PA3B27ueW8kRyLiTpuXHKeJRY/nzD1KRQqtBDgNdX+Tm+lnRP
EqbZEB4X7bnbSEdCvj0/AgmovSqfrm2XfoNh43UN7CVp56MlN1mDCYazb98DC9ak
usvUWThEp10Am5n0HmPJx/QTfVhY9YPwl08ZUlNT5HTG3oA5ntEKpUNfKaPx/K3Y
4QMxfz8ZZRtpbvsIUJ9PkaxCwudeHZcAASB8Xavn70Dzmk6HSvF2VzpZGNwvJJ+r
vAbow23ao68GPFtcW1OSAIegazCe8heO2oRuO+9IbeGqyDC6E+nE6KKzn0p0Yu11
vgXgWslam/VwT+GVsiRXmcYA9MpaCipHR/m9QH0rH2vpMiJj0x7hGM93FcJ+PpvV
fuweGQ70TU1C7aH1BV5AMjG8aG+ZUoFfo+nkLz1+kbw7D6oqBhfw9++6U+wcQm5i
JlJeTBdVeMjxaQ81BXt5pb0kTGN3ho24H1LGtTa5JozFas72J/13K9AbIuDSY+hQ
KX1F6vKyymeIyl277Z+af62uBytRwck1tOb1xL5KSf7YYuMNxwXQd/a2GjlxUULO
nn4uR0djwueR8GhiAzckRvmoyeJ7+VdT1+7vWl/ffhutE57ImXMyslPXGlr+r7XH
IKFcgsUrVJUJDyS1BRPM+8TdyPwx8bgxmEBUOyhFQDkU5esIrOOeywaggoz7zrIW
XvtD8yg3zCNvnyRw/DopXwJq2v+H8x+UR3YtyauhFVRHRkkuqjtP26nooRHm+Ybc
G5mt88MYHQSKM3AqDLdH5w+hOQCZcZC7JB0XY6j9yN7Y3KQLRFB7O8S0fESLYFNm
t0T5qQnOMtpnDDO9ohwxpgWDt+9Emzp3nb3OsSumO9fSzuR93N/VIA2SrYGmIU4Q
GDogaa+aWyB/UOUdhN92PDctACkTIepuUtTmVm93H0uwBCeEu4wl300QDWrKwQ7a
mP/tEXleQDSYLS6Lz0v0Um+Q2x6pMUSviFIsWq2z6xtpDMrjrKTzBLzO/I4GJ0P6
j/WRxd9uvBf97SXvuF9IoZdM+ubIcAEbyhDON66K0efcBEtoHYdfc8OR5tcvPz2i
n/6JEJR8HRRSxCL7I/m4DVECh+V4gZ9NepsfrvlOhRryDxdW3Y5tEphsAREwVjkT
rBpD2O8JBhHlu5rEXym3VZ4nNgNULohcGTeKsNxUdQA81ySPBjoNOubXQoiZIW3U
5J050WWp9BX1QogBlnBMJnke0AKa4C95vuuDLCvNpsGHr1DH53giO37yjmhe1ZPl
XM25N+7e+A7Pp15oBpwq/z0u+F9ZNVSus8HEr7brgvw26jYqqVvlPvY1fRIjz84v
C45RsVqtYIfz6UxOVqVyTH40wBgNCOb8uprxJIOg1JbNAffmmVhO1mCRGS4EQZD7
FsGqEL/bcRZLMGJXnee9vgHAlnr1Ss655eYpjOVJOBIuuX+9qo+n9CUhb9RKeN8l
Cy6Xeng8LVWFwbm5Zi1xxAlHUrHKPxPWxiOQJrhCHBC5IEll3Pu0GMSO/yptW9nd
5R0ymSFf2GtV0cvfLP/NRBsBvZvFjCMxJ0AuckxxDRCGJ7OZycacPBbSjwKlR/0b
4CrRZ+S5KXaE2Jog6/r+MLsyKnA/rJ/PYSBsoIUInAks4ux7z5UFMCLZ3vf5HApO
S2Sc3h2ASMhyDz1FHRSGvBZsmnH9GsIN2H8KLvGtWELi8q9Qh7ikoAWkzL/xSO1t
jfX2BWPIiXwOPwL0O1XzOFcNFgLeOq2aQ6/8nytx1IQFL0jsMA80rOPihkpyVaV7
RGBPjvK4c/VYtFIkXsnLxauErPzNwaQqsBYDQ8QgiHAr44AIoq34sOpoAiqTZtS7
DPkyhusc2ByR1/enrqq09NXM667zovSNMDvRfo69QNcyIPWh9Q0Ryf4ClKYqpwoS
ECnZjSS7fcNgfBrKUToNP0u7L/Vyh/UDDxHDWhnmYom9IQeE2WLmiGuwpU1/2txq
f4TSHob25Vu+xEo8mXSWVLp7R/3oDgIBmbqo5+eQsF2suQqqtECL9pP6GP4dEF5V
5nCKSK8W0zT7HC4nRTqIN3S7wVPFctiPsGrxVSB/2kdQUYHBB7pCaOWkw9TEulDZ
n0DU1ipwXk0Z3jHNm6wTG/YeONG5465tMKgSjsNiLPjc+cmIHKnmtRzghKpkV8rl
7y7GyFT8NCFjYBFKyPfWA7KCA8r/WJYO4WQeyEhhFekcYTS5yaVb3HZCtTqqoRSq
1G1G+piT4ZAqf+Yg0NBuxrkCtKFIjqXHtnh4dTA1i5t+XwX2g5IG7meQlELXzVa4
Zz/8Wj8o6kU7pek/g5CJJiTHZZxUaNJF2kf/Rc6fnyTtyrTI/ZhM6B1hunjwO4A7
Y1+haiaTWfkQByD1sE2sxUPfCcCMRxvXT0aq0EQz2trxeWWvTBgEFiSNMDXLKVfj
odvJ/BYy0AFxNdA2BXH2eVxUNJ+5iXSyQUwmrbt8hN225qd6oGugba9+2qZSasm1
l6VIE5KPfk5+XuWcLIUzwIkZEkqlKuxFGLHXem1mccWkblG89xcalPCM40YbouTq
gylxPm2FMNns89Yxk0qMCSPZpmsNFa1SAdulngt02wOTBVOHPyXdGXbryZRb+AAS
`pragma protect end_protected
