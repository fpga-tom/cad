// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mkf+iu26Itk80aKSOTDP0qNWYTYHw+r7RF29nfwqstdnNGTL4jXzY/D3Iz4r3jx7
jXQ76PyBy3fILRHGhfQz95F7td/bI32n3s2Zj03tGI+On9W2GVkoHK0lzK0VwyJa
oxvQS8Dp4+jKn7Q9uoWCEuG0F/f/wLHFwe3wxEa7Gw0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5088)
jo89TvuQMiBZ1Jb00SELO0QyAGjvG+nsrYHmvEyaGW7f1geNhsZajvDdtJc+I93Q
EoL9nl7z0ErwBFTvIl/CkSULfmysUGcsQco46zq7K/WHZ+T9vOZoJ9Nb5SPMR9KP
DoB3yVeEJRlo9+zzV1X6XwB/ES/ivossOEdlB/dvn7pPEDOntorWDe8DSFeSOEzJ
jLcFKFLjTKC3OFqneaLF6bwmyTh/2VcUigTWt9jzq44o38OK1vYPl4VIIUUZGc4T
oFojrWNbFaxHZ1KG83Uf+iMCRXhddtnJDnNDMPGQYu2SyFOFerpvum9TETWYZy+O
t27tMHLFu3ggCk1UPZ+dFOrwAMx2wjRl4FV5aTzKfxbwuMZjvTNTDwtRR5samKWt
Io4ORQ7sKlVfboFpXiPbHKDRIIRjKpjXQCM6Q8kgAs4kR4ZiNDSHILJCaUgLqJfG
1N5Ju/KNPqYCdD8iTCE+4H7pWJKPC3niY84FTG3u+3HGRSpAaZctKB07vWg1PvHy
byOeLsM+vXmLMbuuNmksliisjYo6AhqHe75/zjyIJECV6xAcz6XiePd0hlzvLnuq
BbPXhIjPHnxzuJVCsjWsZeKv17y7YLYEfDjDyW6MSfjSPKTl7CV7Ory1gz3HQEu+
feXSdyjMDQnq2Qpj83FwB0WaWCFqASAI4G0X4+QfQA2RVFXrNnBMKMug7n2z3klb
nmkTBq5woS8rLHaebRr4uR9A2PSYnCngEMh5wWkICjVZxxqflrTj3oznFlBSvYp1
33xdpKXef/3VnHr90vGUGKDw+GOhulAUNUwYvvkXtxDGX6XhIOKuRiZbiVMgw4JH
2KfrR/bJvRzE0k39g0BnjJfaJFzjOBVNvNT5o3T0MaKsyVC7hPCybE5+nwRz1KQA
Mf8mgIuPhrlDkyoh+pQ6dltWhCbvYXIWj650tZmqTrKMQg2832DRMNc9CU1IXP1H
PJY/hOpuZBmQzwxvbc/9zmGZ2CedZyh269aQV5B8Dwfdr4q2I1cwng/GD0LchEDp
sTLknA/9DqefI6pGPbV9dCYmdSUwJ8aAvawftSYbjFglAXISy4FdNe/EMplwP9UX
02XewCPgNOIshP/du44rm/ouCWk3/ymYMqSmBykB1ese4gmwuBt9QUcYZc3oudXy
VCoa3m/oOEQDsCjy7jn9ofv5/nEqQbYwMomsaZ1CzSOXoCk5AYiM/7o5VGjmG84B
92SegQFQXg2tGVYsfd1SGHXCUvgmB43CR+HuzgCAFVQlyr/wDSOl08IqGShveFTl
uiDQw3eAC8tUeCxwZe0dI0f1z5V7WDPi9nOHhRtUzw4NDb+Ez7BVsLOzh9CZjwmN
7P8dVNVZ298l81oBn+gxTRbjRbOCRmWj49k3HHZ/BduWLej5+oRf57CeIx8mCYnY
Tn/sC/b7/1aqKklQuu8xGn+fHMqAZBcu9talP36+LWBLEPn1LNkTMAUYbSUlHQWp
z9OCjzvF/bmgX2oDp2v5ZaFxo/Y6gbP+qpDU8bWSC6jdeT+ffBLeHJHEqdqslcXa
S5dtpGF4eHCMspTV60DGXpOBQafXx8d1IHUJrsugfxH4wJ2hoMAVHVe58yH/xcY2
7hCreYf+0zHQSPyjz39jYfz/mpQj+4rSp6o+ZWIrIuwDM8uzE1/8lBkquF8F+j2w
waJ6OlqZAIvOPc7gz2O8cKA91xg0u+SQndroKdDrNOjkt8hUghn6Wxx8VgR9vcuX
8bO+LC63hxWlpqGNJwzo14mYA/V650jJcwJ6S2WTs9+OgUBoZlRmG4OmLs0cr1x0
50aHK/WY3BvFeSXt6W+gD7cxYBnNozijqffDkhXQ/4VGCXXAmx+rlizmoB0b/sXq
CdJ1HyGJIbuMUEEmZBEBNWrSxY7aFGjCY386RjSxev8evXBUA4x/uk24hHOtHQCY
oL9vjBsCfqiJ5JMWE9rp9mIZVAa9Vrg/XIi0HpMClVPkyURDUYACLhgRHu3xmOSf
0xQb36wGeAlZH496XffJ7ceERlvHxW3MMqDKkhvBcVOMjVNvJElyK2Kc20Li8QUV
zakq8CNYIBWe593nlqVs8KsXzVPr9bwIxFkdCQe+GVd1ZcflSXUquBHu25IiaOI1
r9+uKL70knLql4ncDiWg20r30qkvLdgOvmyorfNjDWMUUaN1a3zXJjxPW2yBCYc7
Ug/sLQiI2c1SlulgMduqEKWvFmy5d/tmP1fAHMSs+zcscNUWAIj1zNGvs2NFPVQF
4aEFTvCGDGIBTK+EN9v3jUrfYwF8QDvM9c9jBi/sRkNW/KLrP0Ytz5FzLkPD0MZN
RGbhuacwJtxLAD6PvcHsfRes+gn6fgV7hRnN7a7itKJAcADaR2ktQsjZ0vCZY63P
g5l8FEpRpHJUMiKcdK5CmL85KLMneUcFHOsmNXuEQ7Jr07fEJIhc5T1OQqN2JUyc
DYeOMyRvQf9fTh4LNuIFUCzbwDYMkLF9z7v8hrRf5q3gnwkyEXCx8b4V9X3fCMnb
BQ76kNg/4RQoRKSrCyVwMpWzCXYzMPBAphJHkzOG1I7hH5pP7HN7f8u45FF+8wf+
KlybVLU+LkquFgDYKmxlSTxfmQopZIA9WLvfu3Zqylk5d2HhtOZr8jBuV42fSaQs
99UfzK3WZhtu6758zRODntxEksOza6sNHZne9eEvExmgVsfKxvaVLJ2jkht1zAck
oK/80n0H77nlQ+0hBjZYTdaLxMfb849pM4WNWO+ChxTVqIJ4DTx1tnG6qIuhkbSc
ZZvCaiAmGz3aRr3Mxn2cYmWhvc47sL4Lzi2aU2edAG4lfxlfTOn4ETbIvGJ1Ow9Y
Wj/jXkmVrkXfuB276MrzOZb8dxFIKJs+GR0ggtDE89e6wdAqfzFBo6iNkZew0UXz
W9Y75zNUmuUFp0fpDb/dD36pf+RvaUuhDCY/GcMxSn6dzy7Yq5rwquhFpeEcm8NM
89W0zehA5ZgYy6xdMazOXctlmaezHejZzlfTHrvwW6a+Ws3bAoOWJYRiiX/DTtue
lqv0QL74PFZAnQx9E60d+fmaJfPfx6jkzuv5gsBpoKn9nzTHuDyedbRcGVj8LqKC
BGVEtGpDjhznh2Z1NAdDZEV9cYbrmVRPeKN9i/Me1MMUISVbDDUBsXbe+9stFhdi
4EZcwClidxTa3kFMQNs87pF5c+U1xmk6aaMkcin56D9SACB+F9sPq36wuQCHzDAx
CMyK29CxSn+fKcLs2FTMpas21Zx76NnlzrIIJ4pfvf5z8xlHb9fN6yTA5M+bVUKf
9nH9sI6UHdlcPAUOJHFxEl3rIv3sUHh8hDXg6otoL/bV1yA8NCcelxzcvXxNuAaF
UTLaSUhl8DMaKX52lvUSKRS7eXkhT4aZpjZ3xptGoCJSVBqkUHLBiiWABlZABLl9
jK28kjs7OaoDig9PORxFuH9fXZxS0T1Dh8s8+lxqkOMl7Hv2kY9dWq+2booLjF5v
+W5zG0+DtL6lsR+EpKN2UiuAUYS7C6EdVdTpobKyqr9eg1DqT4VNY09+zbIIovN7
QO5oaah6HQqMAIDgHuXbRSs/pqRHNlgXnfpS/pBTjbu/EcRgwtfoPJC6n6/+hvcG
Lq+MIBIpS6E7d86AsHvJ+kjj+ZdrSWplNfuo4SkOI7PkPL2BtRh95Kd/pkcp6nGB
YEi5ZOq9jxYUk00f7Fy0afLiAeSxIQBnMBGoIk3ea0TQzzRMxwOTdu/vnMaw2OTG
6nUQK6+es71s0Hzk6f6eMcS8VW9SF/DxOgYj+OeHNkV8KGVb6ktm/dkR765s+z/i
5oLce5pktvWPIO7QZU+GXrNuPGHnx8mNhSFe9vCnhSLEMJMeHcZd1+xOvqMIMU8m
V2yK8Bp+LoypfnL/jKYEr9fN7lZj5T572zDUZLYgyZXMfIcEobqOUwOjBqhwkN37
g1KO3N5yxuQHQjY6+MO1GPHz2M5hCkLZEMypHXD/SHYpG2Y9XSb9pTiOQKelQ3LX
wxIshRlqQDgHH9hnIEuwLCapOpnwhOmlRKTNQpDkT+TKaPFGIcjLdlHtpb0F19AI
oJ5SAXdiBoqAgZr3nSGA3xgk/727DH9UtI3jZuw0Zx4aynryBCsuYj/QqhBw45i7
YLTxzFQUoIzOcdLzw33L4jBdG6dGZ1z7+g/x/I73x64nXHzEXl0QbDCtWKPVm9Xh
1aQiR+qZmGvNKcOznok7hiGSrrMsLWZexK+Pe4Fkiwyp9O0cfSv3UBp3LH4g9axf
0N6mQT7kVmCvPaW9CpCs0XkmVGgzHjc/NFKPgInznjngwlx7cJ/DWVFmunkgZSvk
EVI7I5OrNKqWP89H9e5PwvHYdTMugF2QnuAtSRJn8LMe3jx9D/SFpw+r99YlSDQ7
H/gwLCCMwZG53eZDpbBdjFw33hPnJ05cqKdtZkFGS5IJnOBoSLSuR8W1P6dbZm1g
Ol2feH+ARfCDgbu2uJWv/4oaFM3ONGrKiXqUPrr0ug6XH5EvIRdP3TMqcFCFBSAA
En4ahttpccrolUkjgI1Wc8NtEGiFvYpbKkHBdOMj5SA+ozvtpuv9R7x+n0exjjOW
OzVJsOkJQxXRFSB2CirX4hFP0EMBOwRnk0y/0jy2F0Us8GY4bsgAEhfe0GPoeef2
XbL8hNrW0kz55IYXYNbQtvKCVISnqX49/Xt9DKY/lvaDHaRaE331M6o3dFLy1ITn
EaE6ZkXMTgmQnfY1wh/5SgcYvfM1s67kJauW9LI4efZ/AqVfVV/BlgbP9nacnQlB
CT0+7LNlunKtPkIqvYchDdJtGib12gyxdDu6qleOCeUGVgMbdDq1dx/SCA+gDXnS
QgHn/z+CVjhZqcAZIjUVHO1rvHRzW5L0ZhEVN/4t4FHcUQX+GAJyeMOnMNwTZ28F
tMwBFcZN7VZacRFKjKVOt0Q8PovTP6j6/oNj5JAg+hn9lGmroNUxbRRkNdOnJE4l
YKsojDwo0rzNIGGsyzO1PNkz2lrSaUzWp/X90CyqBiEB5DtAjR32UmXum4pTcNBK
Gy1RUuEHJKHb1Zk3cgGDpKIr5iNDxeoYJ1tpCPAL7w6UeevZ949YxPv1sPqARj8E
A/asGGjWwzAZoOps3dbSyPsgdk1e7MvA4e3JQ8QuWh+MHueViDE8U/kezFE5V7ns
eCajosR9OeF3nDnPhkYzroSOAgDonhjHFtFpV/H28FCSd7AfX26dv9gs9HPVbk79
PA3wN78tIhlb0FRYv/xqGrd/3hawTiyJQ2ycdhgmB7D4Iuc5yHNz9WxESUb45lij
9M7lrDhapLEslMiXSDhlpubGhbQSSr/1JBvsmrnXHanolTFhDodwWKpTfTKeJxWL
nfi0q66GVLffFHkuixAMUwlham1hXczTZr3cJlivVQ5vfTNkDMLV/L5P67eEhTqK
9sFALlC85LSQbPcVWp5lMWcuA3xKdjPvMXXal3pBUo0mqHVHdKUo2b4ehZ99TSEE
i1PNbv3x7yT4cH8RBjOg0YGoxN3RaylCblQYioOVW7dKwpNvcoTevsKCvMm2CPhj
PMp/qLryu+4CJZDH0Qz5f0v19CHgdUW/NclJCMlG3jpvjuB2LVJGWphWf5km/TOi
CObMGAIFl0EsRPJAtDmjEf/6BZN/XqlKueT8MS0mvQLnPV328HeeK/DkihVl/++S
zvMDFu1nclLZImMmuvKMKL/VaexGxQv59BamTD65yTieNU2QXoyTE/zcp2qIBkX7
9B4kaOxpMiksZF59EPjhf3hKX/DS5g5SGAhaqoUcZVHoBZFbzGtNW/tvMztkpFAc
FliEpjisR2SbIuRDMrhlvIbhug/j+GxzkK3ZwF3Iz7fjE2zxxV1EMBLlJKCnDVHU
+Gilus1Y+PMR9E2kh1RtKHipGKM9UYXzXR75xjjGuEcX2GS4nvYEZUkIkLXcd3nv
KIfSKbjx0PKnAKKFG7vzsrFN+FDd9vHMOkIT/esBlZqbm7Ay+F/HE3u4xFDzhSyD
d5+mDGRR8JRnWGIw/QZbr65f9pi4kiV8TUukSpD6h2KSTBqWfq9RvSsQfMaS8o2q
1agqvmorF+6l2rbapCyDM+8VWuVMMKajT3HXcVUqjkbwgP4ohHaaW0Ua5qMZfGk+
Ct/xpysvqBpqiiW8jXW45eS5Jijglk4M3qUX2Zi8CIO07YsCcIMociOXjDkJPcte
qAabrJD9fE/ejtvfmEDahQvM4ZNY4F3BI4JCG8jboxdK2cIdQ+JktA718z+tp4Hu
O4r7fxSL1zC6gv9WajdEFKEFkZbiR28IZWqepUU+VykUfhlGyZNb0546b/B/3T/X
Pl6E30CjsI/uS9KAXRHLpXtBiEXVR6NhJHj8esoQuFaevbaVRCYrQQZbr8FKsGKN
lF+wtdcEKh25IlQdLidqHMR1vKsAu9KkWgNNbHTBEAiVvP899smdVHIoUJiOopUs
Z+0j6e/34VnKmFMr+1jMbuBmUXdEKYjYQem0JnwvdV08gP3eGc7pb5cdf0MftZwL
KIOihg2ts3VcrEJ1EMXyzsjr2zOIM1uI9/8ASCB3lOZSgFYz8voPHwCJNXrP+tzp
f9ZXFiaOTfFt7u8nx1/b5Af+6vNdoYv50HNqcnqsl2SANpeVqIb5dl6EtvWqV+Cg
wheyRR9rFfrdcrAegF4MH8txda6MTBwFmWYwKSgu4cIKhKVT5UB+WdX8TENCR/5j
O2lx5lfsuIdX6GP/4xDq7jL3NUs+ZhBwlwPBoZdJ4w/I3SDYk8ep1QweVqmG2Rpd
VUKjLod1JVkg8myFN6g7TK54XKtbtETHFvyNyiCowL0+yzEIlBAIa8UI7jbIgHus
`pragma protect end_protected
