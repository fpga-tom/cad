// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:33 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dauqeakoS/kfoNOcHI1XnUxScTM5eHgZg2I8HH7b8XFTojJoAYqM6ZWwc6Jp/Sz2
zXVIzdu9MnPYQQ03p04/BVMC/R8kMvBV8gYhqVm0ixCHL9ArGsKkml0EAbL30uIe
BYR+O7ZeGU42BDFr4ppu9lD9VlAKNNX2Z7w4WgPgtnA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3600)
3G+4Fik7EqIwpD4KPws7fhQSlePgJJ/T3j3VWJu6fVU0uCC/O2CZLK5wHn1NFVbf
2HQ/GEH6UHPxeAFyWmmGoqz9TWB8Hts/E7FCH3g0cOMdNVeGYpkcdsEqaspelHzr
LNc0EUq4PZDcKnio/xEZ9nXwsW+jqYC16uCQTPasKusQE4QXMMjJks80He8CgXS/
hoBh31kiZTEQdCWZnAvh9dwZSGJIhJXXfhCdMswIzoAkWjbYlC5ztj61NV1irVQe
k5Cz1LFyaQ+OcRoxgynBgcfH0D97NODNIyq9qCJXVDFWfG0og43hCi7lGpstwNQe
BybTERNyb/j6ts7RDiRP7zuZK29YBPY/N284K0vFT5GjobpX9/hL7gg9v6nFII9A
mi2+ZxLT6G9K+80Mpvjs9YkIUy1N5KqSK3aPGvJFH/sJWhe/0fZ1Ta6s6QJs4lpH
DZciuVSooIAcr0dDphGcmq0dSr405NlHVnUc+pf0wyvKC3rl8KclRjdawrTH2R3Z
jaf8ByZK9YwLxyfPM+fDOkPssg4k0SmQe/RLtkseilUwy4sU+UmX3vTOnwecP3Sm
w/AvdA6c0N9IF4vvxsC5uHwxrg5JUm+ln5R3R1E1xLhlVMrqPe3y1I+W9axbh9zz
HCvOQ2nbTnV49O9e4mdjruAf9TABMiA7B3vwXHtvjBAK7mo1HvKXCZ25OiCAOJwN
DhhyrlXzAPCdAt5eZBYSi3tCoZDMV3jcwLRdNfO+CEqYPqb9SW3Xwv0MCIwZyCEE
DpLY7ij1lAZkCmp9SMWMHbvvBnzufaaa0EnuvJOaUlv0U4wFXOcpi/MSEt2WliPm
F80hZHEXwceSBd/fuNkRVquK4VgYNxEI4dhahmVdM1QuXlRGBRa4gi4oCdSej0yF
X6bXbvAWHX0dpmJcXKX8faGd6qWswB0tlhk8/whLq4S8ilqQhuaCfNxFSthWx3P+
UsQFmFSjDyYXi+N4MCL+LoRqMevpqPbUe/zhMTfFmo9JmDyCZHqaoEfp1wCw8uXG
MAAg0V+jXRwBdceeQ4iqPRYM+d69n91wl7FlPWKjwOVK/hytCHAdxo6HmIga5niB
ydxu7X54Fuq7KnlX/S+df4qlRD6pwAqyrQo3ZKDI8C9Yni5WrkrkI90bTmdeXTCI
RKUCupWQv0j8OKghTtQAkhByKe9t1X5R4s5T7PFu6o4OLI8T3wguGhAPKwgXFg6p
EymG1NnKd1VoPmXwOjzPfZZlmyJZQ/K6/WFg9cVrsx6VSsAdNcdiNVVjIh8jS1cI
PBAS+URNM0ys6+GIv7atavQDQDqebt6P0yKoJr9JoxpL3T60AalNRAtXU7xdTCek
ckS0fx7sLn9rciuL6bgYyqadRl1xVOHFvCi5hi7uFopzrOFXE0jSAOUkyMSC/7Kh
GNsO6PECr74CRf1QwNf7KqWTYySW+e3186UrFbOmLBkwht/MuM3CtObnFueqoJvL
LIo3Cvu9depkajVr+YF3BjTreLda9qCK7PWFMLfNijNwOMDLSq/+5cWPebk+qyre
6o4ja29J6TB2oMabYhNwJAW7LbS8/OzzQZlQAY6LeZjOPp5IFXVf19K+gJc6ySeu
fArHq9ekyQbhLrlbDWhHQKfXJXeF9L9sk7C+C9fuTQa+1nXPjsM9fStHgI+ounep
v5bJIlzBpC9T4lO3b0jsz4l0YVWIz0suCRj+QmnckwB6UMvxD6e+j/PArNg09YAr
+k3qHQLpBg8MQfb6N7iOHh3FVA1uOTlltKFgPCuPXiKEzmnpIyYo4ULJ9xTM8/Ev
4Z9MNHIttF2rEUbRtANWOKHQqKIJgAu3mrtk4iTU1yEdvoVUrQRxHPHGnKeCSLyp
cjPc8xwNjr8zOBLKjR91ssS6TGAPfaG24h5xKr+lxr53oO1qHEA0hA3pk0Ksj3sN
oPv+RW1yvOE2l6XYSQY6K2U9gEMe6Algnw8mzdoj9vRg7t6hlwt8yLnBtN1lRVWt
cYAfID/AjaNepyMQoV3wS2eRdqAK5ISwsCviKEvzX1SsoSJ9qZyEIvaeeUA2u0+2
lWEN5zzBhoNPmuk2l6cmZd2Bi93TX2uBfwUlxmvzJj1xhgj1hGPWduZK24jFErog
2cjhaaZ3lDa5in/+SYJ7TctVAtxYVwMxRx5b/lhzdbePeAIVBYE62ruZ4g3Co4nI
uhRZAegKDoakleMWguQP54WxY00nfRG6K/hJawJ9Z/UH4cjDDA+cEumwY/ebrWEA
E+PAnwQmXpaR2C3d26fFl9X6bCiPhtZWTXAvs1u8lLijmeMK4YPuKwNZg4mN0nMZ
JtiYWMctlzt/mycB4BmKzve9l80X3VzaNcEc20N8w0dYA0jspdk8JPtBfLv7Oumq
u24FeHZWJg7PCBSDztbb9F3EuZN8qYk51pqZ8qqyJHm9MQO1itjuH2mRsED8mBuw
0i6pG+fy4RuiBVG16cumtu9ORzDqlEuj+EfkadAI18q0BTpva9em8SrLD1effVeQ
WnHx97pN4fenLyvpFonnkm1woHZlZH1H4gVbyKuyN6pNNIxnfHjCnR/gnlWGT8Lw
M0iva+pr/bbHWxs+7Xe+Xnp7fNTexGJR4h1C9Y8Q0EiOx8LPwM4j5ZSymLN7OojW
3HDC3za6fj9DS+Mh+/EQigoBO9dajSvcxUMaQMrPBt0dPu09NaYcIsUthpuHja4r
ucjhvYNO+aQCfSZdXWWBE66H5HdnvjFLBC8evWGZaua032GKFCJLohwunL1kbeAU
99Idr9YdxQSRGxnxHpmxUm4/sR2uldvAgthhcdmbys8YJJgA0LH31Tm8nsvblXgE
jqFn1rzvnKbgJL1YAm78MfABmv69HggKA+QKu8Re5pgzaN2VJONiftyngHsdeuh8
wg8rwyoGzQWG9FeVB9tv0G/dEP1wfzcC2aUcSXXzm27j0o43CsDOY+8tGljtyubp
wgZLqzr7GkEmjjAGr4gPou+Kkkc2NFvypN4c9u2XKOVY8XHCTrxWVzGLJlqiM7YW
4VGhM0mEizmPxASM3e5JZxZIdCVdX5/0PtQmU4+t0FBkhoeN3ufVhwmVL1VmcnlC
4WC5wrnl4cY78zf1MTknlbleToVAymTBaOAB7WnEmKp9+8GQaEUUxe19S4NXRheh
wOypHnrrrVGgDdWTNz1NoNsYF5yvdxYTZEumkCkJIHDLlv5ISk8che7+MDLjHsnc
OFZKlGclXMkGGv72pRqJRya6gBdpTaYRvqcORTDpP2kzeeZpAFCLqCi+6XBfaVyN
X8YyVVFCufD/sPQrCQRAqk3vdN1IwcpnE54lQgyaRB068Ow7BNgz3b12BUxQ93Qh
jIxCPCy/2fsBRA/Uzuo4Ggrt55MfrIYRBhEdRzbJ8OlMG8uN/2GUnCOPMNoZIi4l
J8x9d1s1vimapYSzPzO2CQ8Foe9/y0g2Y2QVj6q0zK2sw37EGHtPPKQyYNhOLuMQ
No3IIYFhXsBp7PtFX85ApuQOI3n3SSAnhQUZ7vZEYkkUhFBlZhwXRc4l1ixIs52j
xBb66KdVc2s8Lbhfq9+y36kurdMSZYNg5G4rViy1I+et+dcoPW6wiQudvBJmBTXu
mdo2OKVykgrvf6Bd7NaZkWeIC26CQiJ1aiV/Ihn+wtPz15xESZKLjWZoSGV3jOBL
c1sHwGjSVf5wjW6R6Dd5T2iT3wCfqj2oJE7wsRrP2HZwByUzc/5FzPmtL6jE59K2
YGYkDmLIu04eL+eUVBJH4AEbrzS8fg7PYL601OHkPMlfv3Evlm6UU6pks1nFlRlh
kivfz6iDtuts3YHmZVp0GCDMcqhJ/PX9gyS4DUuGYv+6hV+LCqmJucFp8HEGqBgz
Y8xXgs3rpu8/rFZaD8fZZGVq8EkcEKqIojw6/ZKSMhgVe1Zj2QeRUCXb3DwMFTJf
sLtbczeNNaFnTf74Hcj+Nq1PF9elpPiSsBN1nIy5k6Qve8xKpfWQrv7RlYqxi62Q
RAQ9GGRs9VglYwpbucm7b2WK2ePchF1lxjYX8E1+HcXQJmnyv+3NGXF8FkJnU8hC
AOZ3YF8q3t2GuhHQPnUgr2SyPpc/JVDXySviQID0p6zR7h04Tsht4PxYRosbNR5F
YJKs2m0DNZglyToQKs3b4NXvxHdRtNX8pFbZA3eYwuYUljEpQhF4lvrBl67dCCz5
WV/2xPucnk7OHR6YU5tWg8AlQ/UfBaFlHhrdQAetQ2hLdQXlHzEMGS+r0kcrXsRh
I4UCzdlSGu9B4nyn6AJydWaJIqrk8thsjlhR6Fzfw0FrniklO9EWBc8ZjHUCJ/5b
ztTeUFL2Glryhl2Z0ewyk1PGAi84zr0q4Wg5xIszh9ax3LeYNzfS1ANl+Xpjovb+
yyqRDwoiFKqJr/sr/OoWsq5IPGi0v+7s1UTPSzA0N4Oo/ufZTHw8WkYabm3TeUQP
pO7j6oV98QIU8OkgCv9QM6Zu7twSmKc/ItT+I26LxdGVOO7NvxPiqt+QePT2jL/C
KcUNBs84+Z5KiucFMcw1TAbgahDyarzNVwMM/i4dYEcXV2j/0aKdUOqR7TWNwrFO
wigOK9gfXrNOWDGazvLAncFizirGmYvZ+9JtTAh+A7O9cB/o49TyxcyY7kU5xGve
VWnSbC2rCy7PMSlgDxSIUJzjQCKbdq9t3CjryXJf9eNhcjRmsSSb86FfL6oPPkvq
QtYr32mu+EVjWhaQ1rTF9yL9pxlhj7KfZchTIVkh1yWyBZRIOD6IYycMSXKkVh6P
5FwPwd1tIUdIwsXPd/GWKUzOjqcvgCI3YWt9VQLbEtWn9s/TP5kWCZIpf/j7WqOs
`pragma protect end_protected
