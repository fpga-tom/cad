// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:27 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GRatEPNj+1KetlunjilVQx1vRXF9ambosDhLgEhEuLY7jAjy3vQX7u7GFHYWI0Qb
t6iXyC+8Nd3SxYJvLJrH37GT+jr1ZP4/qULm5IeA95ARvqhev6ME5CdD7Gow91eF
oFFKG/6EV5OxKs+aV3NOCEIOjf/etiF76fB7PIbBDDA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19632)
EbhYssxricxp6fYgJTjH+JEUCpmSSRHzQ+LcjGqxoolYspT9vBhWXZ+Bwf2LdmOt
4sDgCbVv7rbiJOKFFBbIVJW7xJcDFmAojKFM99gaD1eO7QrkWYL4Wza/RrxVE+Ey
TXe8A3JfARd9sSn9FlzS9uy6sSlaNrg8LV8DiXAbJ4cjhr0RJ6DX28ikvsBttnkZ
H3QQ5CKamkGq/3mHBFqftezsiMcm0LyMsKRqywmug1XC2Dk7/rB4CfXakptZ6q/d
ElJ9RcDMffZ8ZilEOKgdeUNoW26qN690pE+Y7eBdDxokQhO3q40ZLbW24hRWV6yc
phW/TKi6oxl6VDe9w5rWXsHRDkVRIe5lvE/7MmcaF3lzROkrDL4b75rq5yW73GBD
X4WUoZBloyP3zS2reRqla3BllR54SrQyEcYIz6VwDk5MR7YTjnFyw3ct6FUhBVyj
3pwHahiukUdWlu+yHYBtondiGipT0TikAYHoFgisXZpaXJqA5Ks5ilkPKkISoCAh
0fLtSqy37Q/s9hm31AxLJY+49M59QC5twTBs435eFd0toP9nafiYL44Cs8dIhFtd
Az8qdb54MxqvYmLlheiS++z2FBPELtp5LdvBPOkTuHGYgl08ovrrEKdh03a6XjlJ
6wc8Pj78yW566sIZKWc6U3lbPvDsiGqwHxyiZ+t7jyrk2ArgwpT4AZwLy5SDDkSE
/l77uFW5FzHbxfYQQzxxiA4rttcAuPtuWEajyAXtF64qGcLz43kmSu20ISBIcs+M
VATTMyS4jsMNwKHh9CPsMSIcTEnRBU0YguOpyyIhpe++DrVdutqbiE/q5PIUqIlo
02O9zkKtfM983zFhqz0icDgWWedpjqIgmNSaZsDnxid+AJuDqHVDGVqP0M1h4Vzt
KyB3AwZTePetYGEASOmJxQNZC4yMYzlks/W4HFQ9dVOA3nVkTZOhhRoRoRyrjelA
KRc/xA4khv5cbYCP+RBr5V2oKRUDM/xAQFaRcUrsYM4dLBnym3YQsO0GQmrxs3jq
2axovU7+ou8ybHHUL990JZhoyGSx9LzCaGk5zcWRn+seCGMFNUbJUKaaLvnU+g/0
mo1WnRtwlhjMNL9HU2t+g5mPvyBnhPN+Xkpk1eMM/n06Gytex1Vi3xz2I/ocwR8U
aUe154lAh48wcwkLbSX7dwo8fLQzfMU7CHud9f+umejdDKLdY7vpr5QhSBYEtITs
JjzSNaQHviNpwrIJbRmMG9vhZiwmvg1q/iuiqn+FG9J5ovDfYR3EMCx67W7CL88V
l186dB75Ak8V2HLCemnEKCEEfvJCSRkkUoozWeQKcRYrP7uS8up1jxcLQB3lxNzf
l5sYms2LMy1O0wfMvev/kGCVdrQ0pqw+JFbWk3hW6jcaz//U1/DydUEiX9hLZCTv
7RVhVo1G5QhIuOFGeA0TDbHtekQvvBB4I3CntG5qOXarlhFLlqBIN1J2eqA4PD0L
0HpemiMFW9jYmRu/oQfZME3bkaFWp1FWqLG2TnZTSHa22YGF/HsA6W/ZuPXuvMg/
6R5x1GQW/dsU5BBuyT7wdbtSrTGaDb5R6Nsh8DIgSGretYKIGlxOqI5L6d10lzCO
Wb49x0z+pp13yLPROIw3oBvKqp69WQBJgNqXbaCLJ64Lm4OrdasX6yhDyjGmSRLM
oUqbv9Qf0Nl+cdFkQGe1/FVXggvyUPV+1n4s18P1Ld7HoS4rhz13D6I15qG0/jWQ
kKlscaGne/LhdGpf1AzoLJbuIkO+Xu1dWEtPJnC7OPAOu4+o9j4OJeQp056AjXEM
Z6CPG2G80fpQzUETYfusPrDSISE6nz4gOhKcoJtwWXHIDIElKDZM4pgx8k6tDzZM
uMpD4l2TDkGh6k4Xmy3IgB1Ro7hfOKp2vgCp/+O+QwqScHC5bO63e94uj7ippzGY
BiKLLjx6aEKqQGF5Bt5QYnLJaiObMpXI2I6wg94WY2Trh2Vy5QCvoA/yCrVEcqmC
/49eHIAmr27+zF5JC7wD9BmBhm9wYpmRepscYb3Ys1cqrXKfBR4mJQ6ZQpEX32Xh
ZdibJbKSodRhvM4frD1iF+v0lWenq9BTpPVlO7srWq88EeWtGgr3iy+1oVU7Pyo3
Hf2d+7CtsZgkLHZ/S6MnDq23srk3oJ0aGlrNwbeaECy63io6R2gyoe1G+JCPWWGI
za98GqFTMr9AA3iGbqVwZiw/sMNO7m/AGVDxI14QYQVSr0dSEW1ikXl3+9QI92TW
goHUSeQA5aF/z8z8H60BzsU6yU8PHA6tc1AO/U0kBB0/YdBU4Px1+uXoCmWZsecf
yOCg4KGaiXxJtmd6ZLf2FlwCSAzlRwPb/KsjvByINHwswVEQyMj0YasrDNMlacR5
J/tF6StMTuOwnb+7hnL0bFjeen3264uap41WK5Kxwr6uh//O4FafcFTnp8ImlfqA
6HIAoSqu+PpMAiz2CyxKlfTzSp0Ol77LZTMF6zCbmlw0E+s+xKOFffG7PWYfzNGq
hUhkQenmVsZrhBs2o/G3VW5KoChvj5mJjEewIjVRilunw7B0e8iT5S5tTDfpLU3t
kCro8kjiRVZiTnq5jO7qPZZFO1RbA1F1hoFp6Gal+h8E5N40LCQHeC76THaLDqEX
Fz+d/33OVFInCZfe9xb0KSM9/YP+3Fk1FVvf+I6/9IG/gf12CBEYn8vU3PkPvayl
XjKeSuoT/qy7cZMQJ9vTBEtnnQQUg7gL9LCRyPBxoatOUa+D0fB1HYn2+RPc7Jq2
I1vOlY47t2JuG97wJMb/lAb72nRcUmpwym+dlCzmmR4s6WPJyowFXOOkN+F6sl3G
RHzezcEcEFeKedofilOOD+A/SGN3TQbNYXJKYwr9ifxbbUth/Qm3AOfXIN1BIrmh
6zSorsSG3/QVGKTNB5zUIMWR3Svpe4Clr+z/TL80lEJhhlJ6qDVD9u4wLr8ZxN/B
Hk84tVXkpteZSQaY22R3/bA+DtlrcLbihSgUL/BLce5aWyNcbDJqWMooPmahflQe
s9bwTZ7rDzZS31lk2lq1BGCgNCpcNlWg8zzOPSY8YI0KwDOD1W0nr3abcBWewvXH
oSEWBst5wdDWYpjnSB4ZI7jtIOjD55k/IETtAa54PalyNu14yiIP5Ag96p3Pj1gN
jx8J+O7Br4C1v0jcOv1vFSKJcYNvUHzy4OAbn2mgS0lc0LjhxsWMWkQhf+0469Ac
v9fJxDcO7odOiqBvZzE85uttV1lryyf4BeSNdy7kqxTymawpaQ/D7IJESmfZColv
1HKn3bcmYhHn7s/4fqu2CEysMJwqWu0YhBSL0w9uqjZO5TYu68SIyzQPMuUsKK9+
Xc9Z1lo8/7PT7Z5d7Ec4a6SvsjrY2/ewKTCzpQqRpYKGLtnWYTXWq0ZROAEi+wvm
SGuytET1my3JAWqV4V0P3fjCF4B+ghqgkpCsw/I+AJ8xsohGHuMEEGbZ5eOYLDV8
B+GplEz+bzOp7UeDkycgxUExO6AGjMZsUPlu5FOfull6C8MLIJkfcOOOOY7thjAh
BRMILi/XcYP5DGVKgBghLgxiowXJHNYCNhrMo1+1Nu5p9n2v3vqFv8fkQ2b3qnrX
deCHNy9ZLNYUttIJrRYg2mdL+1hbpp2jwleXcoAJrvq7BKqBoqCNq3cYI+nhX6Ei
HBDcEEn7JiVY8t/pEOHAgyzq4ov2dezk+TKwROJVPKOJ8hYBNt8gHhOJPd8gDpJN
4VQgY6hxhde1mx8YIfkUlHudaCTVTEfj9vkjtQ2KEE909CNKvWeuRPdiHPD9tEUr
Xgj6ThFSV6b2u1iD0XuI6ZLHs8W7pL2jKjTv2YlAmlQug83GAbwo+kgipbH4J0lk
iJl8xr1QOYfQf5gHf7dBFvADaTwFwCV3R1ohu49/AcUXRp4Pg+TFkRXA7HRB9V3d
KMNRObV7MZnnC2jVEI4H1Cj4oFHJ81H0bKOPA55KdeEuyL5pkMC3lyIQjF+gVJ4U
KgYw0XfZyruQeoFSzQ3X8CEE0oR2rg9Fhm2aZTLpURUe4MeLvIyJ2vGc9WcexZ0k
2kKzqkkxT9+z2+PJl6MwJd4t6uGJvQEwG65BwEn/vwYPUqLEsj+DED/1JFybx9ii
xzv5UMG4m/S0ccf4FVqT18lg3m8+QT8hqMyB4RWzLHGjnoPgt/zbpUZhAdIqs3Q6
EpEtpCid+/nuvm+BeVuA1L5/YA2juDcCEfPnTR8LX7tsGgSPcjz8yDpyODJ6ZpVz
lrlk6L0KW6zzawvQEymP0E4+dLRBkckaO63mceAvcfSwNRgjqDlL1PrHn/n5NODT
4uMtsd9jyfrHAKBdRBfhqpDZYnt6Nr1vf18c98Sk4yl9wWdUrbc8mGR0OpTQZvJ2
MoxwBT7ybbq8+Xr6cABNPxC4V5DDxllJsbJgAb0UTVmcmBQ+AT2DypaT+5Y8QY0i
fzIEz7Sl8GCXwv0P5Gd39998lgi7saMAogtQzuyZ8HCk+WFuGbAsxTcUUEAx8x2y
CZhQempURu4Kxj8tmdScYQbFwcyuOhuTg/+s1pD16BIMQCSQlBQru40vvClb0CN2
uavep5dSHe1yp7r0oernuvblfRYth9B969N3EbzpneiPmOlilt5AgySmGTvOKGIF
kxPnq/HyU9Cz1z2SLmM/gdQS0Yg+kCIab0U9697CbIKX0z9Qvky3s1dtNmfMtfN2
mJkBM3yfqiKpKZBbBzNi9ZfT7XtdqP+G3wnKDGE7gpE2MxEYqXQ8gWdmDGRJyI2Z
pUoVifrexPj2PSfiUTwMC2j/UWNAdgm/186eAvaRe5SYz4IuB2U57I2aw6eMHDTU
+Kq6/Z5c9V3GnfHxEgAd2Fok3EzPzWA7ZFP9AnSwEqN7YA9MLdOB+I1YwKFDZxJI
wfDDQH71UnivYdJowLl3XJw+h4oi6WX6jAaSB7GFv2231o889UfSRW2sVJCw+oVJ
epNbKYC3QVYGDRME0Vt4RLiMIli4I5wqpITn+QcY2j4by/aPwlSrDcS8JRCIwZN/
CDr2cjHUE/UjX6kEZTuZz8p3X9aLhAFfIQfQ7h1M6MJrYDWaP7EZppJ2Rj0maElT
tUtEcNAYhKW/A3r2Fw9h8oi0sE5Lxtoztm3PDtHxh7ZuCt1TiODoGoaarBj8oq4s
Rfwjd1/3pB3AqXi8Uo3MQQxljN44CxG+xVynkAxeI1w4OJbqgPT3elKNNUsKaupb
qj5hJ8oiJBx+Yo5+ZvbsLuuPEinCNR6IBMw8q+AFWcDsxY2cxXsoVVkh8IKbOnJ2
kOytCWL3F3ofZZjZYHhpsNXIwqBw0MbtQOYmhCbI91wulpd+4MN3xkyZDSxGdoq7
xne4m4Xflog5eko2x5tIb4gyKRNRiSIevbqL3kt+4wk4Ezal8sOGrg5493Q0CCLO
e209zSCvz/pyjDNBDuZsuqblTGzI2kUowtpOPm2l8sezfXrQf2v+U25GPq3Oa3wt
Iq14kUcd8TPG6S5QS6hboKzYxQC3ACRAHvBFSqPYnapYWjYuxtG/l7KMyTzq1kxe
LPjC+do15nTI0PA6g6EsFSthXmqhNwgBZD/Cj+SP0c2D/jVjfiufP9MvgE9bF33A
GXP2aoIXz9AHOvBUsfrk0pkKVV1SAKzdFEMI8fAT7Tiz3azyC2yjOf8jha113Qej
mHP6VaANBVVuagPvBMczt3t1WXjJYO0diOyr2LmS7EIP/693nO/d0fo2SEcnUkt9
sxYFTleR3GyV7xwIXf06wQnF0aX73DSi4tZlanNGIRjAohZObpkRohpFsuBcUlv7
hr6xpT2BxQOpU6cG0QhuJnIIPtNei5B70Nh/FJfdkQR815y0xUCS/MZVRQTeFN7h
HwU029+5AvM3/ZKF/I5BoVAGaTnXvfJ31xg3ZGP1URMhRbBSAZ8n8+iy3CRNKDW1
9SCuuHt+GX357I/Fo/lY7kemISyb3VniZ021FSvurjBFKLVwXIutYLwWV1efh84T
T2dBBcQ97pjP7x6hHsu1x3dA5zNUmMgmBQiglm3NlmKA6w0EJyH7DOiHGsyfLqWZ
sfSg2w61Q2OrBNvnHpBk9f44ZRvjTBReQkBOdtPZcEKRIsZs8TJAh0MuM4ngkqtg
GD1qqIhRaqVCcZBK0jCQvKyFtN6SZAmKy47+a7JDgWt/BaVpmo8BUPPMNeaq44SX
N1Ncflzon1sKSeQLFJZPdw2qqZiLoT+Ca0YB9EA3YDumdz8c7VS75nQvmUFsPiYI
IcxnJ5dVcISH7OQnyEPlRAvDpq+mdmoGIRKAXJrLbI9/m1/vxn81BC7CBIpggx9s
RsOOy5Hxg2N+Vf42EVnagJGLR7jW+neWqE1V3qOyT4teHjH8w5YLnTMGnyWWhb2h
VZtJCZpflYhSLRIP82YZj1JiVRak9cq48iFMZMl9pZfsOx5NoJrHUJpwiy/3fWOw
UVLIKL1gnx4lkaFZZ1aiC9lydCTbP/mKV2OCSvFRz5Uy8IwomYw0vdN+XN6yH/J9
j8IX+5HDLdP2LWyjgBZfIUdAypNc3AwAGuF8sOgoKb/MO07diaQiho6dM5cKgmsx
SKMmlaqk2SGc05QCvQY4guVxVixNAlH1dSCHrot623wCb36KeGDqZuTnUl9Xvoo0
nYlRWVD0SFOhL0dlaW5T9ux4Np7k4h7gimgI4Mgy7wwukmz/iSlKzDgI74xIape+
PvG0vybOSY3Rp1EYLY5xEDQTOL3V2SlaNnS0A06uU0NsargzXKcq4JpXXrIVjD7c
bnQM5QfGZVNKDpYxQ2tBF8EnG6xfR2E/xLmxFIFFvtb443yutfKJtdvtK/kUx6eU
ts61m5c1oQMR/rBc2qU0hvrR47vbWH3JsXKjJOXs2eAUOSBCdBS2DCOTgJgXqM9D
03F9S8m8L4NHvEYBVwCXNCXXVa1AzwXXd6w8fySWlCPfOr0ymzRwI8DMd2BZzgnI
jY+pIqy/3xpRgmv3aOsmqMMK69BIVLZ3GKmrKI9n7fcC5sIeiKPryy8YNqUK37nB
KEQxUqvp2nqbbXz/xzqbgQEL0vOQA/nAHcaqbrpQw8Blh/ia562BWh6Xl8D6Bq1O
azXLi5Oe1bXVYeuu/XjMusQVmmKk7izyJ2SF6ec27tfp/1C1O5gwqeKfklI4IGDT
vdGJfa7yeSy8xjUvhNSSZDyyWTnqRHzaGEqIotppr0m+oiJjyVIOGVHujM6hzl+t
wvujYmi/WLNVC2QDGooH4/5cqWFsQxNAE7u6CDkmX7xXeNNIqNGr4QkgCoKzdVtG
YxTmS9vewnzLgGWmjgmQHJHnE1QR3RuFpUhkWQZm7kXjcLECY4nICzvAMz+Itb7B
5+WSUHhXjzlKZwzUw4qKbWxza0oMCJX9SAGvAItIW4iWPWBnlSmc6eM+vGtiIXOH
FCvjWsXdNh1na4/++vD2zQkc1fBu2lbD+a/ShrE4wL4WvbU96Qr5rmpvi4O2jZb3
n2L9baoUDzzRzsj/lVg9vQTEL26gllip2Bh9ur02EhdXdszNVwO4e7L7JSj0s2pd
hdlCtzzzqTTIQUw9mBKTw3xRcsG22iYn6dE9fs32/wS2y5XiwoYl6rGsut7Ac8HA
JtWnzDTcvhJ98QVdGoHVRinyh4LGvpUGgaFzv54TNygP9iDerwyv7VPu8PfCNNcN
GgETzX0WCxdv3Yv0atC2KhALyPOWoyDGdTM02Z4K6XHUMp6EFEAA/Abd1rXxTKgG
amDyr+XaL3oNLPI+UzEFLdsfW8eOiJElw33Nuh8cCn/d47W9oyAKdDTaTAF3lKHy
N3eQO9BSPe18POnaM9AmTr2VFP1M01YOM8Viv4NZ4O4Qmf+2owUcp2nJJNcOQGlI
NFprlAN3kljG27FvHG8MmAoHIckou2lZAkLfmoauaTawNxlRgaWZ5mdDH6oT8aDo
87JOuRyT8e0FCTuJ8DoU2Eu29Nscddw4V6az4i3LnQO/hT4lDuD8SxHRAmhMt2pl
AWiueUrxw3EVKpN2yF/HC+X6WaP6rOzJmlglxblJSEHziOF+tpQ/Eajh9hYnGLlx
ZFCvC/5xlfBKc5icmLXhEK0WPmEiUlUsy+sse5hNgEerzZz/ZPDjVfWMsajl62N1
faGCsMhIhN7Hz+m0DJQWPS0Zeitbjtv8zLUlIFjPU1bvLpLp3aLBcdm5bwG5LpmU
qaYstmKRodV5/OK5a+jIKwscKhzUmt0zCxBzmmHx1aJ2FtGIl3N5niC6rbNHTBsU
/Q1eIM3mHOdZCN7Ap1HklTESdk8iioG6YaULIcz8Wm4x2sfH72rMZ5uggmV8Mc7D
ZBM8t82DJtjSjPuXW0do9t8LAKTgpfRm7KMLNZzOoNLm3kt8zeefr1n3qVgQSgyQ
bQnKRTbF6BzXpoOPCrdUZYUxpPX0j0Om5Pw0LDnSv3cXWYjjCTHMz1sXkicdVJjP
HR+eO6M3nQdul8sq/gkfHtHWV+fN8tZzvFFvx5R6DG7G0m/ZE4nYpeXFL53pGxGA
MM5YqBfb04xh9vLgSlB/CN2sTyhcc0gsghFe0SyYWa1hico4z/8vtMNN3wZAq8Ho
tQokz7DHtqTOSWUCSsmtOFQfp21EB54Zj3k2d/AOAC3JtTWabMcS/U5BCUeiX7fQ
HpXo3bI7Zry8Snw7gBWgn7FdQGJFEPK3oza3JK0T9DjLIsmXm8YlqdfA+xu233M7
/kmU8mk6aGXurZOSGUElvA6sCK7RToCcXKcsnpP1X0YcrnOsdOi1c6dcEQ3a4gGF
2vImESSbjzB3P7Rxj+12B0ZeZIx8v9hSCCbUD3LWyjm8aZ+lA0favlaGGF2ESslx
iSptLZMWbCe2/7GuTnvpmuiw1YpBbKUNYeBOiHqO56PyrqEvtuaWUN1+BFfCguJH
INdPcOPEUAJIIao0EFo4WabiD6Qge1ZyFbmVMGCT7aM3NMfhqmMAwO4WxSK+GPS9
hgpmV75hCEkeYNt8+QCLaG3Qj5pKLvk0lC6I+MixffKMnKVEnXoJWrr01Q97xrKD
M86kHHcenBLdw5lBKGciItFkvNopEm/xdKkUCP95P8l5vn+EKSepLeC9ys9DGOah
3/xjOVBbrf32U4cM6BMGiZvpNDZNdM715xAXpMNWPTtSdEK61ZVWHLUT8+fSfKNP
DlmmyxCdAcAu1HYAzuhBOjKn//R2DaaKNi34KNmjdXV1Ami6O0YBGALZPbu4VkXx
rNstdD5bvYrBBLHdkeuDE8p7bVMrhLzJx2NYeTkx0mUJ6NqdrQXKFKRhtBYNKqtN
Y45lRYgLSkDlY5O862zEAT/SNowagknyueQiJdWIFNktcb7DxfQa0eCt9sn9UDbI
g9BMvUzALliD0pYP16sDe8FUhDKl2WD6wyFLiiZqIXG8iOLaZ/jZ4nHi/6jBakQa
zbGlU5+eQc5rSXYp+RIO3JKeW3xYgsLc1IKv/A6UgEuTsMu/cMiha6axT5IW9m+P
r7ddu+g/Jitv+wrznyLAKutCVusxLlALzG6aj5eYFpaigoVZAWgduumAn7kHqtEC
trQCl7pyy7OWytbKK4R6esFt3HIDkx4UCiEwc6OBr0eLaUCvoDdUw1mAHsDB//N1
BARAEX5OQrjuleBLxWcPQIF4iO4ghQfio/Bl276+c5UzLzuWRkJ1Qs/+SqDr9qg9
07njeSaAakcPQCZFzemqRD9/s4e+7c5APpupFq6rcCH5QvI7u4T0DzUvGSPIkPH4
8IyJoFV0RaTNxfS0Feg1rG1vjsvAJ3ybMSXiwXVdczrQx5M8Q/JJquBKc991mLtk
rK/q2DBDwsBCMwpCYtR/nPaJ3TsFnP0PUpa/qWpfo9o8qgqQxpKopfvozfBdZ29w
sP0HKQoBEJodc/WOObGUxaHQqlXs4/mYw8cUnGpXfpisKd01h81DouLAMT6mWe0n
rFzR6+gRoe7OOeMXMD0gXDJdrWZV6dqtH/UeRU8vnSjSZmffh1rGAq8RPC85xhUg
snehf8PAVcEzyMLBdtMmSLT+dNuW/K2zpafTEuVMB3JCF3chYt4RtYvjGWBQtV8c
CtlvD2mgW1t+oxdWpzdBp9u9dRnNup4Gz28JOi7F8TNiDR9a75o0KUeEhC6tsSyH
FbbRiNN/cPaVKaKj2Xq5+VbqqLXZA3CdL8HhuFQHrj9aDwGFc3+d0LaODgB/qpex
9We4lqE51c1QcTc8A5OR5sfkOE1TDd+h6pcTc/s51AvBUpqHfnVDrUyNNNod7Xev
JDs7uu8GWVdU4/7cikAlIZa1il6PcquhlQWhPIPtImi02FlllH9QeVNvuRwMud9t
vPIBew1EUjGC48EJWn4kOp7fdYFpGtZtYTC/DtI60Vk+Y5V6yvfmac2FmJx7aQme
K9/z6MQfjvdd7XeJeHcxCT+rc9mdPsy/Qc4IrnFM7JuINMmYHu81h1aVklV00Nym
xG083d4YhyUt0Hu14SHdTObe+aQUK4FymbdVPDhMbG4ao1QiVBuIEiDw23KdCaL7
lQC/AanY57IHWLQjmA6C6DXoVJGVjY2ot7n7+HgshHgaim5Dn0l75VNPEcyLU0gK
C6b5rU+JVSGK0tLQYsC2bnfslvY3xdz4/0xsBWukCkIRpjyb18TNaxo3xnev52N/
Y4A1Gd+O7e2thBeqBUDjYVckXiZb+cMUdmaS8+cxBA82+9DzR6KxHIMNyra4q9vA
uXLdlyEtc2hPy28oRiw4xDwGuaiaiAvZQ1iyPdvq3Fe3BaFnmXN3R/Pd0aJcjnPK
bmkp6NGlm/I1wm7WJm5gI8zOgm5QybcnbvFzz2aCyOR4QF4zWUxizq0OXvEkmWK8
vhiLV6ZMhqK1j8xmRZXRAB1TJiF/wHBRr1eooGhB+23NspvUm7zlXcga3recasOi
07mXtQXPe3p/g3ZAp5UGL5S8ydwWXS82LnJTVDZlMHxcFeCql2L793xSdFvwURWE
T00P/DMCyOJancgfyKggl0bgxytgwWsB1ftd+uXySHKY/V11XGImTjwE4/+LFov/
oh7VYc2gkWov7Dowd0bC1fq2CljffWicMVgdw576M96HrPIOxKaBgNH07c4VYYnj
4MwDrVhJTkhzAe0DlIZgkH5QBQc44agp5cWgI1TOOVhZNB0mRD+8bMfdXEzOy2Ux
zWi6z5/UnMHF+YljL8N3GjTg6fgBUf3T2xcIN9WIgEoh+jsOSmzoNocdESkdLnka
W2fA+smfu8LXI1p3ym3MZWh4VI/S5l7Z3dYYAmVLDWYCDEeBEhAwVIhRpq6nKW+1
VBqBh6c/4rJB/snwb+Xt7hl90LEk+K6rbSFnEYyCeL3wxojWYojzwUXbHodpWIPl
hDdocrJNJJ+MXbxSU80d80UgQqJvss7I2FDpUOf8zsLgPwPU4qumJc9wBGYhjDLU
ahoboak/2wmA4MS6/qhCI70qRMMxlyiNJF+O/4jwhUBxGQmAmL9sbfjIY/9Eo5ie
10TiqbhxE7Dq28HPE2ViAb2wwvsmKtdb7+7JwPzOli05chMGNECGzTDXQP90Eieh
0AQp1d0QNmTalIAZTsVzu+aRnPtFkf4zVOfCFM3AJEkfSJwgVLcJoKrO5rhY/SQu
REMfzeuXEOWB6UuN4tOcxNd1fqqeQRklqSzwRfSz2aUg68yhWA61k30AkNIYP77s
hdDhS1ss+g6l0szZpMBY3CX0iowLDieJHX0N2anXWu5PfhAvzcUCYvyv8W/jS55V
aJn6eetgy9IzmR+rbWlUbDSNOjSif1OT9wdfHP/8MLkYJmG6bdgKmRmOAlMLCOxz
4sg9hYZsoO2Y/NmImQMmufmBXXlVp+fLA0WpsgzsEmI2MS2C95SQqTXO3CGMj2DS
R81MVnVEiModBgEMhxhbRb57/3PLF74Y2T/OE0l4ULOabKrq6bNxRmiqvhSKx5ZC
AY0swtj4HbO4onwYCPPX1TUpw5MN+4fEozYxD0Yb3qrbMgnCxQKnj6ryQfe75quX
YkSby7uRT8X/fou0M3+IPQ1xT3TIcLzZYaX+dDku79zFIphac1G2Ao8gTV39PJfR
mqVO+cslGiU9SwBhMLNx563G+mj7qX3wgbhi49kyP9Te04JA95hza6mLKj08MDl4
9A3EJhovQuIXU06rXFlBDBlmNK/wz56MhHIrUEGyA8Oe0HfHB232fEIcZI2wQ6O7
6RQ4rlS9vDbcQj426Hmt8J5adw3JIN21r0KaYEc1dolEEMVZtnyfXuSi4ADTOdl/
zoBQ+53BBbgCShCgvTiM9sMp//dYG/F0zFYzFKUtlwdSINbnby667qvLyZyHr0J8
0QlR+bmQfHmKjUkknE0NhBGA1rpkTXmHL7Jq4tGd/UFah8uBtzHfc+d51ulzWRcM
/3OGbuZxWh7VMjAh3c5Pr9YvA7y+AAhWtYn81FdkOFhJcew0fJsScHWc3g1r3A7+
4Cw2RRMp9NtZDMj4MjvNMDNwqC9EZ7SKLlKJTQ23r0rFP9uozYCyF9XjZUVlRBBQ
kkk6uaqrm5qHntNZ9bO/QKEQ6Z1SamZrTxMDhhok3OSUsjqx0TCNMO6peND+rPE2
cNQ8jDt7hpvCIvQZyLt2KjVCB0IMknK2tkgQaCtpUYOBEFx7NT6byWLKlZfJuNrZ
+AFNr85BX3hZzPknGc5Dy1UxGSdujPK2VJVxhIBd3V13GeRWA44cgY98/xS7dSQe
ikJ5R5jeJdJbtNO71xxcygydYh+RUrC1rL6C2NUFlDd9KADMFfBeVhc85oYCi5XO
2s6h7G0GpAhpMtVOeSMqePVW+uGKZCrhrHlliGuIql2SF9oC7W0Il3+yE+oHrsW9
OwGoBWFPb35KC3Pv/DZWgUWwt5ZnbGCGRaF1ooYNMy+z/PdgMgeoDH9B7VOuMXE2
LDQ0/QADU99YKyLaYwM+q6YR6F4Lsw7ekUKHMMLfGwckZ4K7ZL9M1eOXKWRB9ZS+
LgPy2f+O7H9aJEYuGRp8cJWYbifz08N1UXJ7H6IB0X+lccxSCavmXqu0LyzRHJAS
NygBSAcy+Avk1BN+gADkYzLqYXx8d2LpEPIdjphPfFsgvowpxHN117FbdMYkALXF
Vga//cAbbXcJA0TpGZP9KCaRJwE1nebB/hxZHdZ/A0dZ/U2pgP3khzBAyIjApvwA
K9rsTwdP4r71jubefdVpuPZO+13lejZDbqOxpRMuGcez08ZAgn6aOw73AKvwvKoq
jCi4ZjMkTugOpRtYBBDeV7ET53REugPJcyvdyKcIyoJRV8O22VaKg+/KrSx6YFbP
FcR4wwE3Hlxtlt1RTEkLHCZwU2wwWt5xpZ5w8GTWL9Rkx9xM8d0HACem7fZRgrVy
H5Y5rmsPpxqWzQHbTcp5X9iPmxMqCnfYTK2NNnQLMCTnD5nZ6RPpntgYG/0g2n5L
phHju0FSTBWSX6wJbPR046jnzKBJfaG8bYLaVmCbzSNoZl6x9vju+xkGZ8nO8eJW
hRJ3IEKTtMCl74BboPWcOr+dsztn5z1d9d0kx0TG0eHDTHZ+qYXjmaYxmPnzQCyi
lI0/MkKev//lC//y8/kUNlzprPwXa+Vl31TvgPMRw9Pujpxg8vTAM+2DFkHV4emw
Vj3UaDe7fsgb6ZmP/A2Alv+PcGPNtAWupDgvmdWTn0MBbhrMLBvuxZ22tD+QqC+s
PUeiFL876QqulOI3sc0GQVuhgTKq1kR1KAr6tiDBLwQnjjPk9CeVzTCBnUlBrKm4
la3gHvyuwqvB4ESzSNo5qWh9whDXXrkyqV9TfuoposJzHZgmN+3ATPiwpF8HcEb0
MUxmUtIjqHdAD5oY/vaiOFdSQTpWFbDTKOBj3CsWQR1r5vBvZfi0mD4A7uZ1n5xw
78FF06IA9EY97pS6BYwMqaUgPXG1FcFISZOKWoRXFDxsy1DJXhlUGKSk1XqiQROb
mtYK9b+2L2pyBPmBR5httq8kqFXwLuf/ixxYHLwrhTgUqlI5smgA0/U9ZQciNIUX
y6OG8F/HFACX6Z09gMsuSJwjNa7A9HfxF67pc28nm5bnSzAemDlCljopaZ3pAt/T
BsbemZ3PBIMBiO/4rIdxGHq1hZAGWKYUcNcAfIg2GgUKTg9SfDyyEN7rjDP5T9rc
0EFrlKvlgo1bUHWjNpB00f0XID6BNX/sJjrr5New1r0+X/OjwSehX+kAXpBnSIgm
XzwApw5UIwS1Va1SBXFH4AiqqF/8pKBLXrT9Nyy+f48wdNERO17a06ScBEgufhu1
52jpMuV6kSH51gukmRGczU8Icpd/Nw0pGjwSTaHj7Ic6WSDh9bJ+iaRfENw6SehC
Hjadc30v2dNQDwzSRdGIrEKINotaF/pLpaECAhC3Lk909m9HVcyPEjK85OKV7vLU
dAFa5euwlESSdn4C7Cf/LqvZz5W9wkUYp0mp4pCexF2/juuZd4x3OeicO5t5yZrh
NyQA8yVX2/i8RQFRcCrx+WLuWCqphosnjZxELEluMP/YCM4OrPbnSMU5YSlP0l1v
Cw5xLGHHfar02mwyhNQA0cGJCQ1VaDoWPZJBfLrQ9Hm2iLYKPmmcKmDjEgvr84rK
sQPqqk0xv0237wooc+w5oVW9o+rNOdDQys3XQambVWY2o58DHcqdqtsAaJ9RXuIa
qg4nPw716mA+jxlnnTFUrZIp86syKtiPeQQTY4nC23oiuZtCHiKmy8pGJYmyDVH9
ujTS1C56giS/nSDuEaejGFyKQd2OLIxA+0uRehe1546FuXPaq6Lr8CAblgW9nDwq
D/J0bjLMPrQFHPQwxihd78t3Uks4c0t4JHEN5ZAnACexyzvSl6QgWbQ4hqph5rX2
iRT7o4abWyrSKkpgUZobTwxwFzphd5DPDHGHSdk6WHi4Ztdm6G+Tht66pn0s7ulC
snqNG6SuD33nT5j48HilQv1Vk/2kqoG2+UI6+LoQNmClhGZMRYsqfzedLEExKfjp
HDAODf42J+vMa15fusMxLU8LJD9wHHzb+dSwUAwnJl2kZJoRyZ1Cs8BmDHNrXx4f
wgyWPrLQErpFXdRmYmsEbTdd//0fO36A705c5+LpUlcsVJ2z2Ssi1rTgYfSaO8MS
+sawyFv0l99uIdy07STmT02kcYp5HuI2RBlGfVP70Noy+PdEnoFn0sRTxeM1jy+c
/vYUnrRHYW8EQ678X+tKoarHnDQLk5i/ZMEFrRVEfton8T7dmMq9wUyJRigW248O
T2uyXvocWU2k3GvCpO6tWKKJBL0o0WG0ZVHhDC3EjTD3Di7W9RCOdqGtIcriNzRV
KI/jncinFD9DSqNGO3SEDD9k5PXRSykTUzAkciGmzb7lWR3Oauw3SsKZRFFpm9GE
ZgctmphIBFrCx6tT6Gqx2nhzbHaFTgP8nl4m92s4IE1uo23Iimrko/1uEXePsmhb
6biGEQP2c1ff1baM2Zrse/FdaEoHKai2wYc+W7B+gdbngkN3JkH4rctnojV/idC1
NC6Z//tzK3st06WkOXp0yR3UR+1sbccSWrVbQnP1f0MPHmwGa30e24l0S3ZichzC
MppoBGDxdBkWVqfyUfws85A0bCL6mT/AjAVVluBlcd/Rq7IXpwWPi3MLLoK/kM9h
xjEOgHvxPOb6OfDO4SFdvi8mmvsJ/0nz2yJhuCEA3Ru1GgyInsJCN5fFJWSu1A9V
0xu7PBSbEnwcLyPTGH2Bo6T7OtIauEXAToAYcSKqzGlWdhwoyviUiuvCxqVshaYJ
KGk1nRSvHKLfEHtAWC6194KTyamIyj7JSuvA8HG97XxDqTaGig2oQEywfHaXOZFK
fmeqNueYynBbDTqyVwCx+2UgpDDj+wCM7yo08PuEtrPjmJgQNaDoXNjHSu+Lqumz
eE/jNBeb8jUBeu5GMsNdzHSTCFmDLDvgS+92DSvLEzDDqxeD3iALk5jFRDeR2+zO
DAjgZlTS/5vu/Mvaf+vqfoUoiiUI3Lho4p7i/XrmAWAV7L9Z3brSnWsX9brghZvs
byq8sc9+qyGfMrI1DyCcJO7XJQSBR+bUUdWO/k3naEYKs+ofun4rPI6JCOZvC/Mr
uCZ4jAH/Wvak3drJ4Trc6Plj/m6KCyDCTgnZQ0rgGnrnvPDS+I0r0pOVc9xamtHq
hLRpsKFZ0mqzgR9+6j4zAxi6hNHkKrLnuFiqBuAjH2NfB45TQxb3RdWWsulY5TVJ
FfmnstwqC9osvR2tVJ06I4zi/B5Ga3Z9c9YiQ/F9JqAL+cFK54u91cSKElk4doq2
JYo1YIxcBevk41z3FgmxgNJk62/BcAx2AfVzZ75cvuD6oZSvrC+mJW/GlUixpBnK
rQ+n4k3Rg15YnsGo1xGSTP1kr1a+k50sfKr7VlPGunQeqKACivpJV4SNmw0BAsAE
zE4gbNoCZxnlLOAvGIIRP/BZJt6kL4kiHiFK15iBtPBeyuXLLZxrwz+gYP7+lYmM
Ri2LvR/RwaJdytNxp7r7zSbQReMFpDTQJopg7U8SoewAOb90D1P6W6sQg3Du8a4r
Dghfb/tDPWFlDNqqzJIdVtuhC6aQDLG6L9b8ROaJS+LbzCTTbYJ6MtQrYKgvSSHh
TywX9/o6MTc+GVqRnpaK8LI2WNwfe3ATAVNj6U502cnei76QyiOfivMRfSx/unuz
6IFIuq4irwfsfJ/bbmVPNA8KY/PST3Gvwv+bqGTmNkxH5FYD8HeAbCbt5KnQWAaY
D9pqzrJiA+V028pDtvLAPqdfxI8k8HWRNmAH0fuMw5tA4B2NbQlim6JJcDjH91hC
k6x/jCRV8l8QRDdXSRJGMpXNo0W6hzn+ouphQ3K1DKxn8q4u55aXHE+MTLHPzSxg
4BTbwmSvdsghFns6YCKyyxWAX/gImxCB9ChgEtEkD3R8/1zdqpJd6qMoIrct5qdU
1hCrTkmIMxJxiu4yRFut8EPC+kQE63YB+Ug+AG2OqheS0apFan9qDxZJJ73aR2tv
qVJR44Njm60wFQyuYQao1jxUWIvaJxFvcmTxib4T51jwrecKSVFPDwq5ZuHacGu3
FNzPhn0q6f/rc2WjzUF1thW5ihlIULHV1z6PXwGd0fDsNWb2Z778sNAtUkWHmhh5
nGjGi12L+PeSlA66EnFTzORNox7CBOAx+nNZys4qkLtY+1i6udMfeFBUGtlgAbu7
tCguswUAIhafYsVz9CL8fYzxt4xHcWL2PRJ5CyCPvBLPWFsuyNZefudKcF8Aj1VB
hQzUYAp2i4QM4h7aS8LlJBfrsnuc8ipYPVFSgtTwGRLN60Y5tA1vH91cjVKYa+f6
lZ9AV43aWKhi8QPoEZIirngYjHyvabfcxitYFXKl4Fuj2WiV1AHJ1H6LmOx8vGM1
A9j4/GnVt6FRhBmG1gkmfnkBUs00gv5HyhGUzvFwhzxVF+j9lnuiv1LGIpAA/aSq
bW8V0YeufPRfSCaqP4sDT7ea2ZhsYK57ra3AbkOAFAC/1qT9ofqOkwFe5UD190VQ
kE0HrmQGt6zDcUifWrMq+i5sUBkmWkJ/NXUiU72h1KWpzOivk02SMP8EJM4Y/5sB
Mr4UMeWOUEdZgNVsfWq9F5KF+1dBiEUXAls92kE2fmPxi4km9sBPC4gsy7hHSpb4
PNy2CW0PrSnVdhVRTxNQFBYupwgV2FCsk98D4OkkRRSyEqp+R8FeWeJFldU9raau
p14ND1RlPVGpZxwjheJXyLVuS4UyvH9brc1XQIcAYU1t6dx6cskwcRQZ753JbTnb
N/kwfTVanWzgNeYS8ON7hB6s6BwqNtWDQBO36s8plemmPEREs9ewb7OLpbYy56Uq
k4iEwlNk5P8h/A44m4NyI9dL6D0UfrRuZ2DhuQcZ+FzHqLLdxDrY3N+ErwF/zkzL
6Wlc4Qno3JtpvL3/oDGMumKmRuKYtG+VeA5Ud4NnXVnnxbkC07SqLuLa3HIezaPk
PxDK+JCcOLf4bnApgxCJeBgIIsDUNUJD0WGIoQ4HcU+CiPuLecS/8zlbEJ4HXkS/
6dPgngimcflcturyL9yeB2hAh9Om68xkkN/U4Ee6RWswguU/5F2GlwvryYk/mGsP
k4mkRLgJubBceaKCFyldD+dGUBNVP6QWebXcJU1tPLVseNlFGpFohi73Bs413YHA
zTLQEc47fz0hesJY2DFGUTIbj2vtwywnaxtO9GQ1Ivnh+C4KojW6CCMe6nS6ZYEb
tadcVI8EuBmAtJQloftgNPec5robPmNveOdbf1vh+IWO39eHxmUvoQAMYjQuIarm
5VrpybUIs9hKHgWHBoIs4ugWlD3cjSlktJ2ajYVncI3pTWPmeNN7ldqehzIN3k24
DDiokx65Xf4N+HcqwDqO5ovrJKVtz45JhNzAJ/U8sBtOrp+/l3t1v8BRFCZvYmJS
pLqz6/UWKJ4Hi1uSI7m6Ibz+TEZQj0CN7lIWV9HYe/8SDS2CLB8BNvygCX3lxY7O
y0hEPo18GoOWfZF+zpQLjeeK61WEEUZDwaxyC0/mxb9VoSBB/uth18OeI36qgOZh
pp9eBcgxrDOuHm47gXIMAECFshYg7NTZsyv+mAX+lQ7abJ6Jo1c1DM9sKrLB7qjb
Wv6BwQZ86vfHDw5Uil5Xg25gxjcAo1ZmZwc5mgF0lJnEYAujgLJp5GhOQEXFu4ru
4puQF5nR3j5l6Mjqc0q+ecTG/bbPKzPZb4rtNgSW3NMRapoCf5P9scpITBVDS54u
2rIJYNLa9B++l1BL8+aSALZ/88jWqtt2xlxs2RsNYYNiTDbyjkR0WsFLl4iJZB+W
C1Kk7g2KPP5t0vkBzIDjaXywtplfnVC5nokA6VySSCJkHdgS1Lt/NGLRTgIwsnO3
dvGorMa4yTMTE0S5r5RAiMuTeix1t/P5L8qBTDtxJNEcNv872OldNWOUNB9rb2b4
+VnMbasOO9GMdIfHwhSE9OnprE4vAqNBbu1gYjUvgyC+K1YOmQ2foLPLItGLrATJ
b7XvvVZPuGuwxXS4RiJcEj7d7QpiUA9ommBoGc9NrO52oC/Sl37iJrSBi8kmNRfe
ufT0iq73ibyoVst3LwZ4y+VHm2ZABn97GF/jsOsj9cSH6/fFNtENxwfUBMKg/dHe
uiFXGzRcmBj6PrRRYBdnByZWxVZoZBYx75gsiEQjKfzVin3g59gA3K6SeecK0AvW
LxxnPasiCB9PJIQRppUXHLa4VHoltLawOlgBv2ijg0TxeTsUEmzYIBHJ2X9FsR/8
fKslFa0Dz/KgSslchVn2Nb9MkM9Lv5SMlQA9eMsF8JXupMSIde0dhWUaJV26O9s5
iCSEQR2JHw2STMyd47E6KO4kBrHuDJfv3NyYij2vVpYyOcG0eKiJ8Xpm8cQgfUdt
xvc0tVuID3R4rrZT3sjaduzAOccnK4l5YihtW7oVvT14oPx57Ob8uBaCKcay5qqF
MwL3JfY86Otaixv0g6876ci3uTLXdDxInsoneRSlQx9AZsdK9+WqvfangCCIexuB
t/cXEVVL7IoPHSJQxRsArJZLZqFUqw2tcdBPUJZtPtpG7YrEcxpC8DWvBLpsATjR
Ik9iqqBOMhhwEzt8T51ycQY0TiOcRx255mkjzpxwrj7Ket6joKYaWvJZmp/YMpF0
oPEITdcXkRicJWrOfYEuA+Lb3FFjPoDK+P5IAeaQnqZRzVwUPPla5Wklc/C4i/Yj
pzoZlGF6wpztILBnaPx92XpUwocy1sqwe92GxRgcecLnwpNgIecxJ6TlQwd/JHFL
7+aoWI4KNrHZGcFbfdlwBtx9Z5oqM/WIGza56SNHhro2+HL1D/vMF4x7XzDH9wTG
hSkY/0ZkE5u1HH+s8OKIs0cM57PUG5yGUjjUqwZCkwCORov8IIRxi8/c/UWbX1iO
XHVjdGSvtW+dgXWttxKwvamSJmEETJpfrUNt2C1MsNoCnuiFCQQ3k+dXpU4pBWwI
ifnYdOI4ZAd/7GvPCtft9cMt9y4A6BJdapUDbLBDhPs27d05zOSETQQY7eYppfoS
jx0tA202GGwC2r+EOfgvH/CTzypxcCqqMgGRVo/O6VKknglhGOdMp53oPqH8CC6p
Qh/L5xFqvNNBUgDxBsLmqCf5j/oI39k9YiwiAPc5qQDmUrniNa7JVfL0IcLKi+DG
nQ1YvC1ynxxQA3bdlGM0QE+oyb3N6joCE4eZs/0z3VRn5zQ95LBuTbHkDN8Vtrnr
4JP5mHcnKmrdwtnki5HMt1FQ41xe93PhxEJUf0P4+LwuecL/2VUU2n/lMEmOuK5/
DpnPOptgG+SJUxlkSCkjxseunVO5/DqMQBuwl4E4vICSzH1CaGRQCeVC1cIow2hs
TfdMDQZlOWBp/4FNEGV74/fTlYMqBeNPuZlVk/t7M2RnPai7PaGT1DqabPW23VSV
qLtDA/G9pe8v2wefwqpLuZl9r9Yr14kVpATXP+eekLcUxGMJR1+LTmo9I2qLNah+
UQQUT648nD1ZKErO+veBd3PjFlJaJM4VeKZIvVBUpMa/E46l3znb4+8vOm9tX3J6
9VVNrPOmrfacAcEzn6QvhGgSMv/hZjJR9o4IN7aR7ZeVH/wIWnABr381g1H+2X+T
+NdOzWxIK12Z+C6EDzKyoLeHB1fsZ0HjK305zxwEH6QViNCtieGwlEPj9HFuydbB
QfZckWCg/15TRDyYHU8TDJBYzauyfqs3dfCKd3+2eisZWqVTrS6gZ4sisxiGk2wR
Zji4vElG5ULIBRye0nHKY9qfYN6j2y5zHrZ2zO6zlWKiUJPNV9AJeZWOy+7sS2Yv
6pc4LIYhpxiPq2pewCp0Fs1qLvOBOpGc/eaKZsHWWA+ehj8navE/FzFYVdCYWfil
XVqB/NyPJfCQKV7bqQZFMSNkdN/btczEDZKGwIHwrg0QXBScdqVDKwgBwb0393IB
omj5Qa+Krwg3Yd8DuTpe0xQgOIpoqqQ3xLj2ACq90GYh56T3LpPnvDQWI9PWjuA4
ZmkFAjzaICZo+ZCC6+CEVMlZ1fp2xl3UvDDbBTIvSN1hd5T/AWUDgvAwCrYOc6ZS
CQmx91zgvtCBlpJKN0dLJUMRN0ib12Fufrh1qWLwUW+vgWOFguvw8ZAHqvohlA2I
qpUTeI2kzaaH9JNqAUP3OAS4MIQI+Y2WKECYrZSNF8nRixft2mhliSPmem0vFQLo
UzoIrz7iF8e3cl37vOl2js4XL8l2ETxu+0Y0wISOkDT2fOicFm10Bh5nwuqx8B8Z
uibPX12/30S/9oB4j8cX/4xfBI71BmCefpbDrmHsPAtlEEQSfsPoFSjvMPgq9noY
2oWmvcbWVnCz/cUkHVjhvMOLtr9TT1s1sSBklTXU1jJX9npYwgcsZXGr4xr4YRjm
rzq7Vt2sXm0FEc7TikegWJIxg6d0RWsWnV8fNLRxR8nniixOj7YTZxHXX9fpuxWD
PigfJkAsJRrjFPROnKlQN6/F2Qy0G3WVKTvhl/87NH/USWEfp7RahD1J+Hzk8ZOJ
9OeEUWkSXknArKDGj0MenIiFJxpYes/EM+tPQULST3G2uIw5K/6wBqT7pc2yFW+h
QZETAPWsDRREi2MKF+Qw9ASIxurp4+9kL9GljfqU6l+Wzxu2sFkxLSBG9WViFdxo
VAGx3d3Fz73biEL16uz9iWs1zZRmWWwaowBvsA7Tn53HqOK8ZTLqJjsaNC2TZPRs
L1SzeUhUlHt38Jm2nfmGwHSMpB/L4UWIIwLJSTNhLHbZu77t5VOU+3QmE8XzJZGp
TDzq5NemvkRDrxTi3JmB/6GRfhY7Pcn23CeVYaXlsEb8CPqm00trXYaJFyen2mnJ
wRAP8iXtHGF0Yv253Zey7sybU5l2SX/L/nfJJAMRzL9mNMOAe4pTrRsv7gRmBS71
PJ2WwA5iRhAEqag1MCaK05HiJeuNCRAycOlsHLgOYSQjMqw87TdBjHd4wVvF3SA9
Zjo0Qcx6+hKIK1TdpKeZZoB7514AQH1D2JjZxuhMxGBzYLxUOb5VsHsVgdm2hZJk
mDqRu4h1E0gdLaQyc+wvce0xt8InkX2fJKbmRh+BgvxpWu6NU3gOSGTQ4tsv/p/n
o7902IkM1vnXTkPK1Mvp5l8NZ3HF5Jo7HKnLf1QZRc4JNVjZ59TKsQymxAox08r4
WZqAnL1jBYYJoYxTVAszz31jzpqeHMkT5M6/ugW/HgVTdo4RgBLf5LtNjmMGWHRX
7PBKEFTPu/sR8aCHc7UyNUB2CwBDgziXy5gmjkLvZE8+LBilHhk22R8E7E9cG57J
lnC1yFBHiMaFR6U/TD28lOJvRHrFRC36qRPLqLkV/TicFbnaLaVYbs3UAcPIuIdW
/cG3CyltnYrhS/SLQe7/d/arCdYeuutb8A2BcdtJzmlDCp0iab7BOwLKffPbAgVX
n12Yba0zp4+Dzd7aq4iRs5UK/W3Bm3zBvRqyK0Wa8gtRfk85aD/mAObkzLGX+xmV
TOqHF18ZpODDB/y/BN/VLuJLgm06ZwVjRT3oUOiT9ePNQRaImD1u0u2SKroRQNtI
o7lbH3pDLnUAq/pWCcRo7tjmFWUasEs+tUVMESjAcU1tooVuDlT+rW1boudkiTpA
1wet1zdmDYT4f2+fwiYoTPqE9ippp/2OeHoAhryLdLMwZz0VsHmKs1YKzlyPKbU/
mZhHc65CUdOZ0ma7Q76Sjalb7FSH61UTkQQ/3RE7qxncErOnJ0vXAts95a/bhCTu
BywqubRFWlqMXJYaOgyCzV9gBnPJ1a2o3jrAE4Xsxm7YwKN3iOAsAVoIqKaG9K8F
lJ2eSrRfvDnaL1BFhPbWWm7fgSVPIh7IMB2kK5qTD/TYdXJ54S1IMli3VBKs1I7l
FzK/CDYDg0K5OtFWm8Nn4GgoS6ljZNGJoBmcu1zXN/dKwb35CVQV29vjtCNiQvAv
lnJ4BRld6XuiJCEQYj3D1lQaKPiXcy3KFoG9Sx0g0fs9AeTiUBvUIRA3S/srbKyu
rEIB9RsMMIGqM7VkaoowabdIidf10Xr/0bdG5soeBXcPJxAquusgwtQem+NCYMoX
JYe5Pyy65dHSCGP4jRiTTSjda7gm1FZQTGgatGo9jfTgunL5+zcb4T+vhjkEe5q4
OxY0jcqUuKIPS9mfm5jbrCyvac9TH0JgNUyJEDBSQZdQkWwXlzlALbKHjYRuq5Oz
I2EOWoiesPk4mCUBPHJZvKz5tPmfUFKPqvOtUGaYappZ3acLYQ7FahrMZonIhb09
oqesnd9xl5OvRR0nOKgTCb19/AOF2crWZL3BFuXi1BMbLhlJACHhJ5qz7166k8Rk
Aqh3V7IuU05HklDJ7A8vJICkzqRrfFbZyWVzxVU+1jk5jNKgEEkp2W1MzxkI591z
xnv4h8OVfBLmHgZee6IVhYtuHk2KWo7Fd0ueymLwG5XplpAMYRpjqweQ/VhbXgfa
x1KK2vGtIazftkNFiI+PPuP766soc7MriDE0di57UbtuvTL68sXxQoROj+ckSv51
p+pZlCidH7/l5y8MWG4woMUrGsgxmhHgtfrtY5SDyblBwzidk9F3t6I6Pf3zt98r
nBJwTgcQE7EQKPDRpsLPnRPvX1vJFYtPeJEATCl6S+wq0lJ3SJa0KRG3bcR8Fgwl
23K8EZL80UOQP9oDpCz4rk9J+TmGPo5q99s7EMwvVUB/dz3CWT0lSC5YxnlHVF1Q
oDCMNm2tOevZMGzigteHawwKmyz3RVzsYSeAzx/bMvuYKAzIk3h/oN1iDvG1pCPv
iT3VrftImcPJ6Vby20YvLX3280fgjN3DLf+iq+fkJ0g1J4khPoLjAPp8b6HNhtUJ
QLfFYep3dAbB0/Y+lNNw85Rg/bCDUfWinFuUln+KXVWonBq2og9/kxxcIh4YUGJl
Zbmo/TajXPBUYWEyJWClUYPyH0AR13LpARsLGvZPzdPcFmZwEi3Wv2n0UeUxFZE3
YMbJLmLMQGi89TzE8gn4WSpVx+LZZA6L+IuuXp4Zq/kmKJ4mf4xTuO4RCh8f+AUL
qQmROa6HIdOo0RjeNd0icy/G1YcyG9RaxT2+SvChlDPd7XMtxsjHl4oCLE68WR8V
1XBIoSlp+fK5XPhsFy8fmKjrjbz8HfOB+We28tMM+yUGKcgzsjpE6PTJS7MoVZpy
DvXB/THLdX0aAvWMgCyP+kLOppIF9zgf6f1rSLeWGzGy54s7Y6CfFA70qOraJ5tu
k3pfvvdzwzH2rvZdbrCICpVSNdeHYkVfgo2PwWbNdW3X+TE7HD/kE0XbQIcHntEA
T45njSuMH3j6pEyT89cjwJ0ubG+aWMTje4fLLap6Bt6dk8oylNgaTGTqqGjVey8V
S4Nqudu8lKMqfUopoLLVdDjUWsdhdDZkhtm8dbP0Nq3SsEaZ2xTbbe3M9NE6J8D1
saw79yB1YAn8KR8bZ6bUCiqpYJFcpSHKtEFVQ7baFR9cWx0Dee8LAgAZRMwdWwh6
3zQxRsLij5RfzC/bHEPuplR3eeA58vBsysz4I+/dCar7JoE00AJc5cDe2XrtClkc
6QPnJ4W8pXl3Jwwxaiuh+IZqd9vt4+Q5uRX2QZkv8W5RtCmJzWJxIe2yE9RXnHvJ
reyGoDCfcYXqZiwZmJwT2Rbqw3AKZkn7G6bF93ByE0uwtajvjNsSwJ9JBdMZZyqz
zyXY6wLgixfBRIX7ZjpzsJjvcSANchIn075ImXhoDWGn+rchNiDg2kMsCKgA5lKG
NgPkxSuHLYcXyiA3izNivjjqt6hXUKBicbvPyHM2eXZtb4XV8+6FQI5uolbM+Ft/
LxeYcrp8Wg6+cKDk2keQx9QnqzAKOvWhe3k+eMZhVg5v7QU9NnXMsiBDEwdQOW46
6p7enm9yQB9fZTeI/BBzm2p1cJBc58WnpDidQnW9dLo72DGL16x/u5GrC3+x1fiV
td7cBHB8wTR1QIiDvWFR1nevMWDnXNLnrmMQ8xT+eUJfOkAR0RojXSSO3SG9IkVc
C+b+3vNvhxiDMYxbKIYUxR3OZ8nWxPhiOcT6JcK1NNrKQsNJNLwIXEpvpsLDRvN5
wOlGhrUpjZePe1qEk2DjPGt3XC5rb2QrhVES5ZGjlVKA7v+3pgGD4ajfdgizU8vp
Kfc93XUZPO2YvTmwP45bh3Fn7I/teK239RctEauBPKISQ8NIZMekzLeLSTZbxN7N
CVBxZQVmFlCQYvH/1Qg5uhGhOXLQ8yMBjS1uPpdpUYI4gnKLRuQcZnsMocknz20F
+BgJlfZsM8w/m1KJJgsZBXWUDd6Wv46N9EcmnUbKLtOUvYKwUI/iV3RROw8/L5o8
vyxMNGEv9yZxDCquPllYA0EyRbDv+UXNz5m9AqduxVEaTTAJ1h9LOoIPYhK4Ic7I
6xdcYY3Ms20d2ciRNV0rAeVO/5WA7ZdyB+dxwTpongZ1bu9qP1uQAd/apdaTwxh5
vIQ6uhjLS13JuugcmMAITiLoisIVVGEbJkK26uC6BJbACrfHn40mZxbppR3za6YL
ooFbDM/QVGhZcowpp/lElN44NgluT0Dc5FXuzucBZn8IAHPlNjSiWSVZ0GYrdKSY
LRYMl5uoavdHh2Id9zzFN2Dr9Y8saCPpq/GJnG6OAbtvCCbAdnOOvmS/aOavHDtz
3ynq8Ssa2ytMLnhB3e2raLWLZALO6xfuWDEKccHD/JPdsgv/dlau1Q1mOu67yXcI
ZYNJ5NeButh85IQ9x0glBeCZrUvQUcHQ+FObHFBlfapANT1+BqAF0UG2hR6C2Xdu
GLj013nK5a4f0vK57xWtzfcAt9Qa2qmk9lOPNnwYcm3ZFhnCPdmmJKi6D+8+fLiU
ivqDLZtfJ8JgzKSWSg7kMixOlW3ttb0u7SY92ghMECSKG5C7qrwu9tmicIE0esDC
X8rnV7LBkX0k84Fr68Ze44L4EAjtNHmRDCDeyo2tyFAg5Nu74RSOUf3n/cCUZaC/
ysUGgdsWUw/PTLvOEpsVL60s7G6VYrKleB2bubnxM9tJR+9JZkzbGZcnm5XYLS5I
WutW8J/WDZwlFzVi2u3wfNM7SnK0PKO2yJZSa58teuisqK6ZWnxeeoPubbdWF1vT
/nqtKdFdJopID0M8LOgUKR+Nv/yzsldXP57Q6+WOJyJuELKeGFIONCfCC2+2y7We
KJISp6a73VhNMiISwIn5IyQU65hOzNz0RMmCWQMwDtwIPY8DNug4cVST0lcQQK01
5rckPBPVr2vn83N9g9wMh7g7WnxRitsh/Ntmj9xS8IOff1RgQz+W00PKwSOOi/EK
cVFniO/F2dtBG7VvRr5KwBnazv6XZ962JYgPasj8XK42bLgSriyFLjupt/Gu9WsB
a/wARmUkGY+ZDbaKUBhomSvtJ/I5K2JP79I9ULB2iwZaYeGY9CnM7KxUR67XJfKQ
`pragma protect end_protected
