// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:29 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bvLoGwDbFevRiMjFs2JbGB6zfYcT40BYPZakSNZAMBaZu+P6ARD7bAks4pXKE2HF
nay3LW1DZ2s3vXZC4Ot+nuM6g8EUuiQssdltr+awwlNhKhun8OFvVkZVHDQdpBTv
l9jZT3ilJmHY6jYu9iwVk13pL3LV02ZpOopm2oI6yQ8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8160)
Nn32NEe11lrD7XNbnmaUd05NA59d5hcQexySYdneRyJl2BCx3XpQ2YsJDGmy8u87
gCZd8rinyAxQrtsr0MhU0gsHdo5aIxVec/tAoZGFpIPc3GEVQhn0SFztoHDGZ+N3
fQPPN+AoJwSUYETxf5/4E7Zlx1DkBuyeOSfGohxafTLt7bV59Sry3BISPePtgPHc
jMU3GVKd02+MTBdZfMuzUX5SDNyIPBZ+6g0cDLmf6h3zqXH9S+ALEngeqoTqzYqY
xxmYKPxRPYWUHq3MfaaEaeHFyo/+ULu8fLkw2kwlEl4YMwmjG6/u2c1KxLpmSW/A
UCyAtOa4TJvZbnMa71QXCGRZBHM3mWqdW3WMx+kEPjM9Xt4zR5RhzH4jx1ZMP1eN
Qcij2DyMYxywt1UQ/MgIR1dSRfP9E+JYK5IzOHPzQGEzj8Bcy2WKizzUmofWlQHt
fr7S38WVwg15vWp+a2cc/JGUKCJX8Lj6NrgruFwL+zTKIF51I5gkFsnDDWwiwX1f
5RL6udhYbiKE+QzxyPoiEaqd5jn1qHnur/H02XY0ipbU9cardtVJhUoNkyWupxSb
c18gUkokVJeGgLn+YEjDkrUXGnODJM7rsAeZOKZs3yjo5HTdnzf5a0oBcyxY1h0E
JfcWxjthpeZDg8XKJtc+NVZ6XqGx3ISGvGTK9jXvDE3Kl48ty5Ykw3eqTBxq5uV7
ZYPMOnTyKxr8YTo7ohgh8T5xcVLkV+DYkHJaLAQrofT7cM8T9DAB7FGuSpvI4LWy
uELI1trjfpVcrFfkot9GZbHQ0W6Vzx6mEC79Th/wv9+dFB5dN/0ZpSaeSji8ikG/
yZE1Jtu9JrpK+NvzTpoGT6qwEAw7FMpKTZMmRCquuolP1MF6hy/ppnDp7+2rhffT
nVG/CXk4nrWmVr3Ini0sxOA2MsHDdY0Ed7b3D11QG9c6Qfok8xB3djj5mYINZWUE
T9HpmVRzJC0StAnV+oQmQuC0xctGYlaw9d9vZizuT2YzqSXyYVnvsd4y5ueesPaC
plkIxwz5/RwJmuKHQMtEG5HDowuMdscSImoVtysQWmy9wYTS9eDSdBUJT9mdowfL
nZCbdcgCtv2P+tzHtLp4ne0D7IcOLUkcCc9XnGXDUc8oDUQ8E90PuBLByxlTGKN8
uHBewlDs9oylL9zlSWVaXTMYDtLpwhlR9Fg2CXePenyDnXhwt/zZSb02G4UcVyFs
pQ2Yj8Uf0XNTxyHG60GyV2yfUj4nObptTZLuYvEH/JKFOGRVRp428PSsTXa5N7yg
gshrpiRDqcSR8n/agSNsAT9uDgLwfSrNdK0RD6etWXYx2NkpNKnZvEUJoGTflpr3
d/LcMPAiVyBKnQwiLgRyOdvRAlaO+UBU77/r2EsRNCM53l01Cf7enz2q1hbQTSDd
dQ2bKQLLsZ1X0znhSVkrLvx/libMa4X2FLbNGH8ACuxCNYz3niVc1QTN+S32WGB8
V0B89KREroygFzbhzbr8k2NEVGbfGnD2YZ0T8zptusT6Qf3zFq9ooNgRkoO9x3jG
atDz4XKSr3CI+ZHxYg6UsxaHQudAjGB9yMle8rLil5RjcxDAEWjHsILMzaMLMsFL
frkwgh196YrKrG0w7TI1Tbm5OA2rCH9oKsPGqaLaPXg4x7MBpH7SeKoIY0EmIn/W
G5VzMtHH4NTEs2SD5cYVOU5iFrqqUNJFmr8jdN5HPxDAJHk4JsBNSf1gGmmo3yX1
5Npb8cU/cwwCcIEw6t90xc80SODp6J2Vmrm1jw53zhpWWVdkQ1jEF4yulONnTd1I
pSmQrdeAXH/6OpYgwQB87tcZK08xQH6h8MEpXRwQYr566BnYDf/gyFkUCpPTblwQ
TPhIs3CXMIPj/HSy7P1muM0++S4Wc4JmH3DS9HFODyvKMziG4R93GMTgCG0IvunG
yPIk8nOQG/yeefrFHRAp0zxW8KbGPFlRfRMZgTzQ8kisiWqxYbDRAzB9/PKZ04rh
Yr3U0y+vyR6X7i3hsGaQqlCTg1xAvdrM3H/VB6HWz8Sk7vUAEkoOBGtC54uFGn6R
9YCb1h3VrukJESmSBJnFRJN6ofLAPWbpcjdDQgKkLvPz0heYqtUj8Y9ewuj7VE80
jPUo5Lh7xuOe2M85kfflVcWRpAyDLEnRhZ4csZgDEqCluIMqtOSt9JUpiLT6vkxG
TfqC2AZw1zZRZ48xmfCpxmwvm0tn5h3lnUWc6ucM+tsBwrgONlhaaPS4WQ6hVVmd
gtwF5SyCBVk+NtYpgH2AMOApzm0vAd5Yp4ER1j0iUIFooFxK2WOHn/NCeNuCKB2J
kMGGpBhHvaUyhmFBM7n5QLA39WVSynMDZTQl9l6Z5Hc9a4SQHl1/W1k/ukf7XC3h
b+B3JItUH87Kmzf3NEAEj/pqUv3MgQreSQCaryvZJsPkZaKyDYprnopZE5bEeMPO
2ez8/8MqfAmvpBjVuq3K8Mlimrt7grbICiRkUl9rbIRtA2vu2cSsa/SP4rxQeTKX
UUYnGUU/HfnJKBPQ+Pg05MMDIwgCU8qljnN2vvgp05qOaLm4m1iKuhyc4/hIVH+G
s7PhHDqSl75d1MNAKB6CmxrtB7jIDAlEy5ATcesEvYTRZwd1ORmNWdMrMQ9kO3Dj
42VLOrpOZ2WZ0U590Ci4qa1W28JostjIKoWiyjyAbmmEpqqjroCXDlaaFj/HXeuZ
sFsOXXakoD5GDhFsYHr56R2zqXn9o3+wi0yrpSFy8Tz5pEZ2Ho/VsEMK7l98eEch
FGenuYcY34UKA/tCmzosil6UXd6N1xvv1sW6k4/XHhMVAHCBr75zftwslh9VYBVB
WOtMW87bzq8p7DCo40XH0Q6MyklwnTWKmTkjTSARif8qTQqJSpU6ivd0HR6cCC9p
FLXiQSadBH/exPCqk49n3P7r4Akot2uNojusJM5jQJIkvQrfsevlqydANcNUuxUt
YAjHjcBwUtNy2F5mIUrln3Wo44xHctreT535lW33xFlNty8ko4hViVURxahhGwCs
j66vwVKY/MyVCb0aXnofwP/EJrmypts/GlcyVE2sisIe0NAfIeX1sNaIt7snapqo
yypODjWR/T8X6AIXLZTCbeEIT2JtxBQ0QpBfDlMMdCYysbiwL6wpwHh1QDCjmhuP
c2kXvnS0wYjHJAkW20AICS1BC842Uc1yl9EGupe8cn5MBAzid4xEZbdk5CbyFuxg
5HBHKLDE00wiRbcGJzpuaaUwUIPK0gYBW6SN9+S0Nw0cHCPgtDgXAh7NYVY+PoDt
mhQW00sL/coyOmPQVXfGd22MnLfQ11U/lxjWIQW5wRxAfdiD8qawne+JpryWmytx
xEsBvAvBn7Y2S+HUm0nyWK5l9Gv12sx0BZvW0ndYg52NtKkKskMtCZMVQYbXx03I
Whavbljh5v8g7RGvVmfhlxv9veXs0uRpBW3RvkXlBcGCkcd2xOATfMovwZkEBb3e
R3xze8IbT2W+wXdG3n6EPcPLFdWuGiNCBJLZOkSatI7sJGkfsXQmxv3UntVOH26B
kjhHW/ealiQNpS2Tif14AOqWAeFu5IB4hObWh7nGfT2kL53WUVx/j73+14as5Hht
ekz6KWO3lcWnP2CEeX1gsbT8IGM9pjYZgDHlSUjB9pSBMlgiMggeKbmEnexeyluk
lTt0AcB8Lwo1TWxHd+wiRVCf451PTqrWeBBQIpRUgG5jJHpxAA7uMu/r0LVCr2Bt
W8u5qBNJE5v4dneNBP1W97ezZ15JPsChcn/gjE0Kv5miYUdqzk6No4LHMwwo5D53
C7WEdnuDeorLNNzqaNa8n0cc7WI89G5MNJ/6NjGHP6ghfHjfU0lByINVM0dSShhT
8say8ZzmvfkmDk57turH1GOTXJxnMJVkoIKxjqrxzhLaf3Ox6yO5saXj/p2/ndO5
oI35dwuYeKUrHpkGHCHpGdUuwuLBuORR7Wj/clWeZWllcwYohqrHMV+R8dnGs5ZD
NKAG1+inyZ19i9VQsXSlHTc9l+Y1usmJkV5k9t+/Uti/3Bg+JM+edg1v3bxrikVQ
cJk/iYzG8ihWNPpIWaNY1KGTDwoEE+OkbEHVx9BZCjxr0D9j3ywMzxEA1MbJJ1uF
709EHSjvImGPusN+v+iLWecUPtzZi2VEr2Hr49mf53OpgbfzaSD5TRkJq1XjzOyJ
jMvtzP6NTp+jjSIqZ/NXq+OmVpQPkhHG7NaRgJ7jmKIRlc+Quy5P3QM8KPF7D9eA
d8cAfGAij3UEUsukGaskCYRVMUNOKv+oLm/UcdCOjt5Z+wkBLgQYAEe8dPMhqT94
GruCwrY9FhqfbSquvHUT4yDol/yCrBxeLAaWcogl99pbWiHXkyxDYzRqEs9c9X13
ZB2Trxk6p6FNcgdOCy3P25QvC5cKAEsijegx2ebOAaK4MhH3GE8Wz+G/+Wg0X7N8
8q2qPuR0YHbSE2n0ravqInH6MCFRYTfyAxunI0F06DeeZauTLAITL3XrCsu1JTwc
OQtzO3AwbqJXBmxDl2JNzxxx/Bp4p3H4TQVmyUwJLmWSXck+Tl+CJgzhLnmw9rhZ
HqHkv9PSTK7JXsB6WMCHmZy9bNEJCV20qWMBf+QlqVC5/wugshnqq4+sO8QBUchy
Ry2CWVxnGXBT3+ysc2RQ6Jh8UzNc+iCLhE9j3J5NKplrtEbtTEQ2SUZilCRv2fI0
1sZk4waNuXzeGn15T0zYrPQ3k93u/oCip57H3dJk9sGvY/C9bVqfjLZSfXfhQCQe
06DvLCN1+Zf9okNc44v44/W2e07DXLt7GH93kJ3iGhvv7D4+gL8Fwpd74p4NbE1l
EcHHA8F//ySEme/76tMF59+TdZNubNOAySKYGXf2iJ60NPnbYXGZIbX3kvtNcEAO
Xa/jc2NuW4exOqwJTys9xwo0YKIUnqSDv1ecDe9F5pE5K2hJW5bRD4uKEfGA26T/
i1C2/oIF+Nd6daKjagqL0ZijOWGzb9dIr6P3k2y+5aaELlERB8ilx5EDRyDQitXL
LsQHNLu/E86KZJi86JPKtWd1LqQjYyfLMMD0P7WzVLSghjdXmlGG8G8YNwMTTecg
csATxLmtZDiNdROM2WpVv66kveuWMTxLfqmK4BMH0kqiM2A3P99YX3QT1rgCCmX1
5bcQOdiWXW7RDdh2sj02DUKB24nZuieJ/K5MndkYuhIujQUZnicH8/t1XZaiJXOP
sY0pOGsKhdcYTMc3Bvh5IGcIc6qDZNFCr77dCPHdenJARFZntA4Uf/vIxZtocXrB
d6tSjyAho7CimkZ1J4SThtj8mJz3el1HpiKbkEMM1pAtFIrl1OXpFMUt37OHgxbB
x5FP77938o0xYytvUNhji+47QNDLG1IUW12vo2xf98tBrlSAcKRzapLCsrXqSMUc
N8JPzW7AJgtZJxoZ30QvjA6fcMloukG7oM0ESRiqosOJ9TYoJHtswZyVtwT40rYF
rpHYPBMSsA6p3N+jhCCq5HNx/RXAGjd8EpIkDAGDxT9l9cxQApr/gQKWiD5re/vT
Tt65qAgNydXwQeLj6gazw4tSPQoQYJn0w5L/JxD67z8EVWGmYrUseKxfpE5rH3Af
oT3Zs92Ja2zrMyMkAJCIkNCjnsh/I3Ib60WerEEQIqIJGMcR/epqG0cbhzOnoxl1
tZSiJmkQjqAE1wmRywCQIWQF/OKyvRg38ybMiWbanccTiFIUcAyE2HAqCkI+Tcgv
a+8b0819k5+GLYyl6jM28ZRtojuJx+8EV71MLG0A/lceSU+p0/VZEGF/hnpQQz7f
X8nKcWU1x0/ZQCr7rSt1EN0dlS3Z3Qz3e6Hj1vt7kpnlDkAEogeWtGiUf2HMq/6J
0WGr44wj2N8TMRI5SHGPu/D/i4+OKL+CzxR6Yatlgf9rpFhXPGReCrt+/RsY2igb
d4tJ1mz4x4blTfB3ydjVbqh0GFYqb1X+cc1kyyGrDBIklUyp+ZNRlQiAqFbpBBm1
ZgZGLcNpF32kLnKwTjB0NA3mdbx/BvE1c3kjcgzqsa7zMSUzNl872XkEF4ELM3ll
0hsG6nz9okqJktC0UVWyB9LOYKheHzADOq4Bq7Mkv+rYQYYb859/Da6ltlMkhgyF
X88L720mqZfP7yaV5Idl/erRB2w3IJXqhrwfQZ/IWzKdnTS8qbMbF8wbjnWQeg0X
IZttFMKg0SyP9RLn7CIjhCpicrQstcklHVqqNCTuxcbJstHLYR7M0gWY58VtHrhg
MHFlRoxnO4qcO7vJXvzmd3hiWDkl2WyQK9eKkxxxtguciPwBGD1AG/wd5/lEpei9
B3BioIOPSisXWi1lycfl08mkqLWeE2KAC6ArbP3xPj7vSRYvgMV2GnWznnwwF2sl
5FQHIRwqjz0abGVO+SWmozOj/IYMin1PXu6sT8ZtVR1f8Rr6iCC4FVZqVrkOOQ4w
Ph0tYKb7T0ZjQh7KDKQK/rOyEIWhjK1l+wGc+X9wHYhD7pfKhi0//VeLuPJiuOMJ
dePB3WgY4dQmOKNWYu43woxkgKIoF7jEhgAYGCwrrRR5NDFqZIJC1G6MM0BJhRMg
fIcEQ0CgHGFC4Wkani0p4XzbXNSGymnLMExqeA6di9jSnVGXtXhk78ZoUQ6sUtAD
g6/K+lGRE/j5xooZG4eOZmvDUat8BZ+mR1lECVwZxAoempLaie8i9sEoULX6H6if
+auU/cTQ3g5DrK+DSjnP9SPSxiCqMgb4J1Hu9M4KJhBjNxYbSVucjDEwHxDp63xx
kyK1RsJBB+PqY5wwBo0Mk73es70WYBn5QgItUjxYJjLqJnOfp3Akr/rEbIfZJjJX
5hxG1Q0e2mXnO+o0mzoT7aTguLfKt072t2K1F2LKmQMeQpO7BycnvM+U8mNzjdBB
fXYpTNqKD/5ADjf7MCQ9jxKZpHnGE8L4N9RNK+2pr4qNGKPJ6hBFJayjMzBsLyFK
QcJiVgHqkfs4wciTtQwoQ5BplTikJnAl6WPpVGTW/OFnS5P9NCgDFKdE/e4b65iD
MN5ohTvzeQQFwTK5E7qP1dEQ6ShwJs02R1xoE00uyAv5EB7nEAeBlaO8x1ozYyU5
5Bri1PMo0W4Nz1X6ZHf5a8ZGpemlxhI3yvCperceIo0FdrNo7MLzLCyfDarXFe7r
s50sPX+8ej/rJuVHIBzVSxHuCr2qYHiVvvU+5ms1EmVOukNSweSvMP/3aSw4kDOH
jLWGbgoZ4hz4FcMuO4MOU7Cpvq3OBxK8cHcHsRrJ9NG8LgkFFtI+KPyp6B4P0iCw
MH6+BEn2adMnhFShHGOvns+ca9Z0Iya+4oWKDx6jMIs061rxMwWS1Ov9Vmo/vXPI
u5uTp43nzYDbSviwNI3chhVbIIHuS8K2Su09qWT+vvr7Syf0L/DK+/ZZPqbeUHTX
i4mhQidulTxkHRLdUMwEyWVoJPjE4GRg2AH2GhJsSIMZtMvOTdjmP4kfBc9DHoJZ
LNB2gaSzWYAcnD/7VmmOKPhFOfuqk/BweI+1FIcrbkbcKrDqjdI+jDEJnnk72aHn
TQhln9bA8Y4Z+0SIOZXd+hGdePybd6BsK40vEXkSVykQf4BTD2kbFnyel2j9psG/
kUXQrNh1N+mNKlu48LYwudYV18fBDU+0jIA6owES483v0NgjiEg8xmsLIGbsBCA3
S7zyx8xxVTOqes8D/gsmFgRgkEl67Ni+KyIYta9IYxwMoG6MKLlBWQPwHkzVRqlj
l6xvPmPedGMFAeGoRyL5GpScAd1cPa0OySLE0q+g2ZETppuSGLAmgJNKZff3TKV9
kWEocHvd3i9spGkxCX1gjyir1q1h8fUL4UwGA4/qFV2/I2/7zZ3GBIGfzONuru7a
xr5b6mbba6pkAcaq55FI9tTbAfWdA+XDRjnUiC/djFOBA+wkA5W7mGM3eZwwUFmG
Oq1Zg5Y2hYvPeXQ+963Lr2ga9TLueoEvgJpeCrktBEY7FvxnYOFAsyLw5cdDYuxZ
6iokT9o+gVGgD7dGKZNyJldvFhdH+7I4DhAqGiF830q3U68nyC27eOzPEa4BD8Jh
C1aQeXCrhYlj3K8ontJtkGoyW96n+TDbnq4vmb6sg0po7N5mNU3Ws3ZP184FssDJ
oD1E4gcX80CcLWlD3kvL3ocshqZ/lgwSd0oMRiLTjLlnj9c1tnFs/NA7L9f63XG0
YsRgzqc48Alq3A3AOR8iqHXs/hfDY0lb57p53ysq0fCMC8fzahxXgEDWQhmGjDc6
7DuWsEyeK8PFeyBcF8VGO43gWbeOYpXij/oF18xlxlvGsVUwzr9x23nzeE3xkXKR
eaatfwsYYUtIBEAe0jM9SP6xKTQiNbEncH/048NueIoFlH/EzCT2ePB7/1yn+cnB
2MrP6UphiskC0vGQKUb/NeKMs5ypfypwr0kGSfQOnioBqkWDvElZU7RDwd0GH/bd
geNqAkEo3La81YlNtD5SOib+5Gwmj8ROG0TbR62aabes9ENss0PmblMdsuaSIJIA
xywm1XTIxLvpfvAixMVpWzYw1Ib2KYtDae07zLyED50Ll+8fyQPbNOH3TNw9ba1Y
/6jEBbT82h+Jz/zBGlWgjAix0+b/vrkb40MYlc91elQPo9F7b5ei/zSih6UQfFkY
SB8SylzKgk5Z8qn3YQt0pnn5fVBTkY5tYVbqbAiYzhvUeiV1zVnyJmsv5N2hHjdt
akguHGtKVL6jwgcyAWqwmVJpL5m37YiWeXoFlnlkenmO6X85PM33EvX6dggmZ8PM
oT0HbOuGwmYV9BFMBw/US9vfnF8s4JurIXP5dmWYr1Yc5tORI67JPlq5iFIZ22sX
onvvYGAS1lyBsOzMCdR9lqNURmEHvLoX44SfRZNX7Obs+MCoNzU7xOydBxT3kksf
UL8RBp6Pl8kRUMIFY9Pjl4u65qggbiubskcz10QBFdnIi/y7bNGQTldzO7Oge5S1
uaDYdfHFAaXsGlXlHMHxOLo1kcqI9IHUFUUQ63sTy3YuByjwyT7biyCohxcEG6QB
TX1NyzsNBQrkYoODGMCbzyChPR720ObhlAp5pZI9471WLfKLofUsaSylqEhUZnvA
8TImOhjtVOCWMUu8uSBRoMqxLCthaxxZ/iw3y3v9DHOy3FhX1sOFEqouclelSSTM
ISt4RNVH0IlTfekvHN0gd7KuOwkVwHTnpkmNsnAHYoAmN6FKiVwmYMhcQEzm22dA
akLDTdpSI480j0gVolUcnjTQycI1o+TpfQf4u2hA8D/ZigHqWz2/P8SlQQU84UA7
ZT3J3/Yz60e6qGtnsc6k5Cj2nzwBNGcegxjmcwtFNVZLO//YLNqd59yP50489k4B
e8KiDiFmQrrLbEILBIY/X1xh+NuHIuYGq278Sa5teyn1fcFp68TnYWowZC6xydIA
wlYOR2kBPvIUfEbj2u4CfAOcLCaRUDiuHwA67dHCaD7ZOG/Mca0MnlrEjzKgO/4b
YRxDGr5iL5yBZLpDMb/p7tj6ZBhu3fegyuRg+CCNqiE1zynaki+G6nJtYMBexl1C
1LbewK1GdVvwHNmlCq/kDqww2+y3A7/hCjvQJjENMhHE4PjcaTRKeXkueHPe2BWs
gWyJdX2ydFEG4Kx1wmjnVLSPKe+HeYvWnWmWPuDw/Qm05iCWV/3mmkDnv5WU0hxg
Xp6PeEJKDuUWc0mtNZqs1wGLXGeZ8+L0vP1bF+ON9J+8GfddMaov6xQq9QDeK6ie
x92zSAG+LEJU/2gJpU/b9BUJXWz/xsEndTi/xvN1g5asNHN7fAbTrGsIPwZ+SoRN
3Vbm6H4MfAsqm8ydC1GCNHVWrWiHp907XXOQDH28OGhF7dPkSGqaMHZQMX102qat
ENpjEEPpqqyb2bHNkMIEiAUtUSuuK12Xg7054okaufL4zp5khJoALOcFmfVmZOIq
DeVfInKHXGiQC454IoHqgakFgASOYOLxqTI9TvKo8JWzvFaZtjPTrQIwwtF4nrhz
9QtAHByms18LBNWcnzqYpeehCcsfQKtBlOb4ZEEjF1LAysHtJAOaiKqvJ4DukOTi
wEeCwl6Ficcr+VNcstLHmG6hpEDkB7jAVRNOT+OCeM5Ap7w3B/irMTnmzpudVSrP
ViW/huU/3tnKcpMb4/baweZUgJ8Tgo1A3uvKiW6SGhGbckvHainQQfFfPzgj34KB
TaWS/aHh+L36U2ROt7/Xiy0ktn92n7QDESTFyBWTMF1aO1s43LIaqmOtty4YxyeE
wE9JY70TNIHObZts6gElCHbAPM4tb3fwosZKJETpNy0AJO1exNgVePcviJQcKjO5
iqtOtS/JotvYDh5WlIZ3gTFUvWPCdtLLjLjJRIErtliWEcdVN8/m/83qy3HaOEdO
f8pWX6S3PE2bc/veW+kLWVa5CEEa64NpFesU2bHeXjsm3J57rVyvpYovgvVYATDw
wvHPoks2/lLtZRvMXavAkLKQWmoVUsNLQW9XEn84Ag0vPr9AQwxgy1JI4akf7Dfc
RE4yQr6B7fQJa82I3WnvU3RsNK6IvGel2rc7UL2hMobi9cO8jq3jeY2YNKYuR6cm
kTAMGC6aG0SbJBrLciEyI+7akcnVkrevAi/noHTP6tfEZeIgKkfnvfZ3aEsRTSVh
e9KwImHGE70Xie7QYdxvOwco3PZv1YI374VFIk5qbj8ELw/6rIVERTpgb0sjL/e5
kPvJObHyVXsbmgcL/mL7hE6sbXJu9CVZDaUgFIxWETRkYt8eKFMgn3ygs7u+78Qc
5lsZ5HvzJ+vOu1iWGxnNQSUC+yMvOkwoGvViACTTm6gT3jOb2M79nLtne6EyvcQ5
RTBhVfj6eHj0iClED5L3VqnyWyHwxPPqBFryvvywKdPhxtECKLxTyVHE9gh35nl6
kDAJ82eFXu3pOCvarB9cUSx1ByumZ9GyYhmQWTqBr9HRD9rc/haMEd4Pi71wyNnR
`pragma protect end_protected
