-- system.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity system is
	port (
		clk_clk                                                    : in    std_logic                     := '0';             --                              clk.clk
		clk_hsmc_clk                                               : in    std_logic                     := '0';             --                         clk_hsmc.clk
		led_pio_external_connection_export                         : out   std_logic_vector(7 downto 0);                     --      led_pio_external_connection.export
		mem_if_lpddr2_emif_0_pll_ref_clk_clk                       : in    std_logic                     := '0';             -- mem_if_lpddr2_emif_0_pll_ref_clk.clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_mem_clk               : out   std_logic;                                        -- mem_if_lpddr2_emif_0_pll_sharing.pll_mem_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_write_clk             : out   std_logic;                                        --                                 .pll_write_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_locked                : out   std_logic;                                        --                                 .pll_locked
		mem_if_lpddr2_emif_0_pll_sharing_pll_write_clk_pre_phy_clk : out   std_logic;                                        --                                 .pll_write_clk_pre_phy_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_addr_cmd_clk          : out   std_logic;                                        --                                 .pll_addr_cmd_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_avl_clk               : out   std_logic;                                        --                                 .pll_avl_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_config_clk            : out   std_logic;                                        --                                 .pll_config_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_mem_phy_clk           : out   std_logic;                                        --                                 .pll_mem_phy_clk
		mem_if_lpddr2_emif_0_pll_sharing_afi_phy_clk               : out   std_logic;                                        --                                 .afi_phy_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_avl_phy_clk           : out   std_logic;                                        --                                 .pll_avl_phy_clk
		mem_if_lpddr2_emif_0_status_local_init_done                : out   std_logic;                                        --      mem_if_lpddr2_emif_0_status.local_init_done
		mem_if_lpddr2_emif_0_status_local_cal_success              : out   std_logic;                                        --                                 .local_cal_success
		mem_if_lpddr2_emif_0_status_local_cal_fail                 : out   std_logic;                                        --                                 .local_cal_fail
		memory_mem_ca                                              : out   std_logic_vector(9 downto 0);                     --                           memory.mem_ca
		memory_mem_ck                                              : out   std_logic_vector(0 downto 0);                     --                                 .mem_ck
		memory_mem_ck_n                                            : out   std_logic_vector(0 downto 0);                     --                                 .mem_ck_n
		memory_mem_cke                                             : out   std_logic_vector(0 downto 0);                     --                                 .mem_cke
		memory_mem_cs_n                                            : out   std_logic_vector(0 downto 0);                     --                                 .mem_cs_n
		memory_mem_dm                                              : out   std_logic_vector(3 downto 0);                     --                                 .mem_dm
		memory_mem_dq                                              : inout std_logic_vector(31 downto 0) := (others => '0'); --                                 .mem_dq
		memory_mem_dqs                                             : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                 .mem_dqs
		memory_mem_dqs_n                                           : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                 .mem_dqs_n
		oct_rzqin                                                  : in    std_logic                     := '0';             --                              oct.rzqin
		reset_reset_n                                              : in    std_logic                     := '0';             --                            reset.reset_n
		tx_0_led_readdata                                          : out   std_logic_vector(7 downto 0);                     --                         tx_0_led.readdata
		tx_0_tx_serial_data_serial_data                            : out   std_logic;                                        --              tx_0_tx_serial_data.serial_data
		uart_external_connection_rxd                               : in    std_logic                     := '0';             --         uart_external_connection.rxd
		uart_external_connection_txd                               : out   std_logic                                         --                                 .txd
	);
end entity system;

architecture rtl of system is
	component system_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(29 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(29 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component system_cpu;

	component system_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component system_jtag_uart;

	component system_led_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component system_led_pio;

	component system_mem_if_lpddr2_emif_0 is
		port (
			pll_ref_clk                : in    std_logic                     := 'X';             -- clk
			global_reset_n             : in    std_logic                     := 'X';             -- reset_n
			soft_reset_n               : in    std_logic                     := 'X';             -- reset_n
			afi_clk                    : out   std_logic;                                        -- clk
			afi_half_clk               : out   std_logic;                                        -- clk
			afi_reset_n                : out   std_logic;                                        -- reset_n
			afi_reset_export_n         : out   std_logic;                                        -- reset_n
			mem_ca                     : out   std_logic_vector(9 downto 0);                     -- mem_ca
			mem_ck                     : out   std_logic_vector(0 downto 0);                     -- mem_ck
			mem_ck_n                   : out   std_logic_vector(0 downto 0);                     -- mem_ck_n
			mem_cke                    : out   std_logic_vector(0 downto 0);                     -- mem_cke
			mem_cs_n                   : out   std_logic_vector(0 downto 0);                     -- mem_cs_n
			mem_dm                     : out   std_logic_vector(3 downto 0);                     -- mem_dm
			mem_dq                     : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                    : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                  : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			avl_ready_0                : out   std_logic;                                        -- waitrequest_n
			avl_burstbegin_0           : in    std_logic                     := 'X';             -- beginbursttransfer
			avl_addr_0                 : in    std_logic_vector(26 downto 0) := (others => 'X'); -- address
			avl_rdata_valid_0          : out   std_logic;                                        -- readdatavalid
			avl_rdata_0                : out   std_logic_vector(31 downto 0);                    -- readdata
			avl_wdata_0                : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_be_0                   : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avl_read_req_0             : in    std_logic                     := 'X';             -- read
			avl_write_req_0            : in    std_logic                     := 'X';             -- write
			avl_size_0                 : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			mp_cmd_clk_0_clk           : in    std_logic                     := 'X';             -- clk
			mp_cmd_reset_n_0_reset_n   : in    std_logic                     := 'X';             -- reset_n
			mp_rfifo_clk_0_clk         : in    std_logic                     := 'X';             -- clk
			mp_rfifo_reset_n_0_reset_n : in    std_logic                     := 'X';             -- reset_n
			mp_wfifo_clk_0_clk         : in    std_logic                     := 'X';             -- clk
			mp_wfifo_reset_n_0_reset_n : in    std_logic                     := 'X';             -- reset_n
			local_init_done            : out   std_logic;                                        -- local_init_done
			local_cal_success          : out   std_logic;                                        -- local_cal_success
			local_cal_fail             : out   std_logic;                                        -- local_cal_fail
			oct_rzqin                  : in    std_logic                     := 'X';             -- rzqin
			pll_mem_clk                : out   std_logic;                                        -- pll_mem_clk
			pll_write_clk              : out   std_logic;                                        -- pll_write_clk
			pll_locked                 : out   std_logic;                                        -- pll_locked
			pll_write_clk_pre_phy_clk  : out   std_logic;                                        -- pll_write_clk_pre_phy_clk
			pll_addr_cmd_clk           : out   std_logic;                                        -- pll_addr_cmd_clk
			pll_avl_clk                : out   std_logic;                                        -- pll_avl_clk
			pll_config_clk             : out   std_logic;                                        -- pll_config_clk
			pll_mem_phy_clk            : out   std_logic;                                        -- pll_mem_phy_clk
			afi_phy_clk                : out   std_logic;                                        -- afi_phy_clk
			pll_avl_phy_clk            : out   std_logic                                         -- pll_avl_phy_clk
		);
	end component system_mem_if_lpddr2_emif_0;

	component system_onchip_mem is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component system_onchip_mem;

	component system_sgdma_0 is
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			system_reset_n                : in  std_logic                     := 'X';             -- reset_n
			csr_chipselect                : in  std_logic                     := 'X';             -- chipselect
			csr_address                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			csr_read                      : in  std_logic                     := 'X';             -- read
			csr_write                     : in  std_logic                     := 'X';             -- write
			csr_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			descriptor_read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_address       : out std_logic_vector(31 downto 0);                    -- address
			descriptor_read_read          : out std_logic;                                        -- read
			descriptor_write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			descriptor_write_address      : out std_logic_vector(31 downto 0);                    -- address
			descriptor_write_write        : out std_logic;                                        -- write
			descriptor_write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			csr_irq                       : out std_logic;                                        -- irq
			m_read_readdata               : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			m_read_readdatavalid          : in  std_logic                     := 'X';             -- readdatavalid
			m_read_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			m_read_address                : out std_logic_vector(31 downto 0);                    -- address
			m_read_read                   : out std_logic;                                        -- read
			out_data                      : out std_logic_vector(7 downto 0);                     -- data
			out_valid                     : out std_logic;                                        -- valid
			out_ready                     : in  std_logic                     := 'X';             -- ready
			out_endofpacket               : out std_logic;                                        -- endofpacket
			out_startofpacket             : out std_logic                                         -- startofpacket
		);
	end component system_sgdma_0;

	component system_sys_clk_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component system_sys_clk_timer;

	component system_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component system_sysid;

	component tx is
		port (
			clk            : in  std_logic                    := 'X';             -- clk
			reset          : in  std_logic                    := 'X';             -- reset
			tx_serial_data : out std_logic;                                       -- serial_data
			data           : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			error          : in  std_logic                    := 'X';             -- error
			ready          : out std_logic;                                       -- ready
			valid          : in  std_logic                    := 'X';             -- valid
			startofpacket  : in  std_logic                    := 'X';             -- startofpacket
			endofpacket    : in  std_logic                    := 'X';             -- endofpacket
			led            : out std_logic_vector(7 downto 0)                     -- readdata
		);
	end component tx;

	component system_uart is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			dataavailable : out std_logic;                                        -- dataavailable
			readyfordata  : out std_logic;                                        -- readyfordata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component system_uart;

	component system_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                                           : in  std_logic                     := 'X';             -- clk
			clk_hsmc_clk_clk                                                        : in  std_logic                     := 'X';             -- clk
			mem_if_lpddr2_emif_0_afi_half_clk_clk                                   : in  std_logic                     := 'X';             -- clk
			cpu_reset_reset_bridge_in_reset_reset                                   : in  std_logic                     := 'X';             -- reset
			mem_if_lpddr2_emif_0_avl_0_translator_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			mem_if_lpddr2_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset_reset       : in  std_logic                     := 'X';             -- reset
			sgdma_0_reset_reset_bridge_in_reset_reset                               : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                                                 : in  std_logic_vector(29 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                                             : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                                              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                                                    : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                                                : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_write                                                   : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                                             : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address                                          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest                                      : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read                                             : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata                                         : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_instruction_master_readdatavalid                                    : out std_logic;                                        -- readdatavalid
			sgdma_0_descriptor_read_address                                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_0_descriptor_read_waitrequest                                     : out std_logic;                                        -- waitrequest
			sgdma_0_descriptor_read_read                                            : in  std_logic                     := 'X';             -- read
			sgdma_0_descriptor_read_readdata                                        : out std_logic_vector(31 downto 0);                    -- readdata
			sgdma_0_descriptor_read_readdatavalid                                   : out std_logic;                                        -- readdatavalid
			sgdma_0_descriptor_write_address                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_0_descriptor_write_waitrequest                                    : out std_logic;                                        -- waitrequest
			sgdma_0_descriptor_write_write                                          : in  std_logic                     := 'X';             -- write
			sgdma_0_descriptor_write_writedata                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			sgdma_0_m_read_address                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_0_m_read_waitrequest                                              : out std_logic;                                        -- waitrequest
			sgdma_0_m_read_read                                                     : in  std_logic                     := 'X';             -- read
			sgdma_0_m_read_readdata                                                 : out std_logic_vector(7 downto 0);                     -- readdata
			sgdma_0_m_read_readdatavalid                                            : out std_logic;                                        -- readdatavalid
			cpu_debug_mem_slave_address                                             : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write                                               : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                                                : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata                                           : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable                                          : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest                                         : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess                                         : out std_logic;                                        -- debugaccess
			jtag_uart_avalon_jtag_slave_address                                     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                                       : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                                        : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                                   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest                                 : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                                  : out std_logic;                                        -- chipselect
			led_pio_s1_address                                                      : out std_logic_vector(1 downto 0);                     -- address
			led_pio_s1_write                                                        : out std_logic;                                        -- write
			led_pio_s1_readdata                                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_pio_s1_writedata                                                    : out std_logic_vector(31 downto 0);                    -- writedata
			led_pio_s1_chipselect                                                   : out std_logic;                                        -- chipselect
			mem_if_lpddr2_emif_0_avl_0_address                                      : out std_logic_vector(26 downto 0);                    -- address
			mem_if_lpddr2_emif_0_avl_0_write                                        : out std_logic;                                        -- write
			mem_if_lpddr2_emif_0_avl_0_read                                         : out std_logic;                                        -- read
			mem_if_lpddr2_emif_0_avl_0_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mem_if_lpddr2_emif_0_avl_0_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			mem_if_lpddr2_emif_0_avl_0_beginbursttransfer                           : out std_logic;                                        -- beginbursttransfer
			mem_if_lpddr2_emif_0_avl_0_burstcount                                   : out std_logic_vector(2 downto 0);                     -- burstcount
			mem_if_lpddr2_emif_0_avl_0_byteenable                                   : out std_logic_vector(3 downto 0);                     -- byteenable
			mem_if_lpddr2_emif_0_avl_0_readdatavalid                                : in  std_logic                     := 'X';             -- readdatavalid
			mem_if_lpddr2_emif_0_avl_0_waitrequest                                  : in  std_logic                     := 'X';             -- waitrequest
			onchip_mem_s1_address                                                   : out std_logic_vector(12 downto 0);                    -- address
			onchip_mem_s1_write                                                     : out std_logic;                                        -- write
			onchip_mem_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_mem_s1_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_mem_s1_byteenable                                                : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_mem_s1_chipselect                                                : out std_logic;                                        -- chipselect
			onchip_mem_s1_clken                                                     : out std_logic;                                        -- clken
			sgdma_0_csr_address                                                     : out std_logic_vector(3 downto 0);                     -- address
			sgdma_0_csr_write                                                       : out std_logic;                                        -- write
			sgdma_0_csr_read                                                        : out std_logic;                                        -- read
			sgdma_0_csr_readdata                                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sgdma_0_csr_writedata                                                   : out std_logic_vector(31 downto 0);                    -- writedata
			sgdma_0_csr_chipselect                                                  : out std_logic;                                        -- chipselect
			sys_clk_timer_s1_address                                                : out std_logic_vector(2 downto 0);                     -- address
			sys_clk_timer_s1_write                                                  : out std_logic;                                        -- write
			sys_clk_timer_s1_readdata                                               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sys_clk_timer_s1_writedata                                              : out std_logic_vector(15 downto 0);                    -- writedata
			sys_clk_timer_s1_chipselect                                             : out std_logic;                                        -- chipselect
			sysid_control_slave_address                                             : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uart_s1_address                                                         : out std_logic_vector(2 downto 0);                     -- address
			uart_s1_write                                                           : out std_logic;                                        -- write
			uart_s1_read                                                            : out std_logic;                                        -- read
			uart_s1_readdata                                                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			uart_s1_writedata                                                       : out std_logic_vector(15 downto 0);                    -- writedata
			uart_s1_begintransfer                                                   : out std_logic;                                        -- begintransfer
			uart_s1_chipselect                                                      : out std_logic                                         -- chipselect
		);
	end component system_mm_interconnect_0;

	component system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component system_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component system_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                    := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                    := 'X';             -- reset
			in_0_data           : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                    := 'X';             -- valid
			in_0_ready          : out std_logic;                                       -- ready
			in_0_startofpacket  : in  std_logic                    := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                    := 'X';             -- endofpacket
			out_0_data          : out std_logic_vector(7 downto 0);                    -- data
			out_0_valid         : out std_logic;                                       -- valid
			out_0_ready         : in  std_logic                    := 'X';             -- ready
			out_0_startofpacket : out std_logic;                                       -- startofpacket
			out_0_endofpacket   : out std_logic;                                       -- endofpacket
			out_0_error         : out std_logic_vector(0 downto 0)                     -- error
		);
	end component system_avalon_st_adapter;

	component system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component system_rst_controller;

	component system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component system_rst_controller_001;

	signal mem_if_lpddr2_emif_0_afi_half_clk_clk                           : std_logic;                     -- mem_if_lpddr2_emif_0:afi_half_clk -> [mem_if_lpddr2_emif_0:mp_cmd_clk_0_clk, mem_if_lpddr2_emif_0:mp_rfifo_clk_0_clk, mem_if_lpddr2_emif_0:mp_wfifo_clk_0_clk, mm_interconnect_0:mem_if_lpddr2_emif_0_afi_half_clk_clk, rst_controller_003:clk]
	signal cpu_data_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                     : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                         : std_logic_vector(29 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                      : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                            : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_write                                           : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                       : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                  : std_logic_vector(29 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                     : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal cpu_instruction_master_readdatavalid                            : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	signal sgdma_0_descriptor_read_readdata                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_0_descriptor_read_readdata -> sgdma_0:descriptor_read_readdata
	signal sgdma_0_descriptor_read_waitrequest                             : std_logic;                     -- mm_interconnect_0:sgdma_0_descriptor_read_waitrequest -> sgdma_0:descriptor_read_waitrequest
	signal sgdma_0_descriptor_read_address                                 : std_logic_vector(31 downto 0); -- sgdma_0:descriptor_read_address -> mm_interconnect_0:sgdma_0_descriptor_read_address
	signal sgdma_0_descriptor_read_read                                    : std_logic;                     -- sgdma_0:descriptor_read_read -> mm_interconnect_0:sgdma_0_descriptor_read_read
	signal sgdma_0_descriptor_read_readdatavalid                           : std_logic;                     -- mm_interconnect_0:sgdma_0_descriptor_read_readdatavalid -> sgdma_0:descriptor_read_readdatavalid
	signal sgdma_0_descriptor_write_waitrequest                            : std_logic;                     -- mm_interconnect_0:sgdma_0_descriptor_write_waitrequest -> sgdma_0:descriptor_write_waitrequest
	signal sgdma_0_descriptor_write_address                                : std_logic_vector(31 downto 0); -- sgdma_0:descriptor_write_address -> mm_interconnect_0:sgdma_0_descriptor_write_address
	signal sgdma_0_descriptor_write_write                                  : std_logic;                     -- sgdma_0:descriptor_write_write -> mm_interconnect_0:sgdma_0_descriptor_write_write
	signal sgdma_0_descriptor_write_writedata                              : std_logic_vector(31 downto 0); -- sgdma_0:descriptor_write_writedata -> mm_interconnect_0:sgdma_0_descriptor_write_writedata
	signal sgdma_0_m_read_readdata                                         : std_logic_vector(7 downto 0);  -- mm_interconnect_0:sgdma_0_m_read_readdata -> sgdma_0:m_read_readdata
	signal sgdma_0_m_read_waitrequest                                      : std_logic;                     -- mm_interconnect_0:sgdma_0_m_read_waitrequest -> sgdma_0:m_read_waitrequest
	signal sgdma_0_m_read_address                                          : std_logic_vector(31 downto 0); -- sgdma_0:m_read_address -> mm_interconnect_0:sgdma_0_m_read_address
	signal sgdma_0_m_read_read                                             : std_logic;                     -- sgdma_0:m_read_read -> mm_interconnect_0:sgdma_0_m_read_read
	signal sgdma_0_m_read_readdatavalid                                    : std_logic;                     -- mm_interconnect_0:sgdma_0_m_read_readdatavalid -> sgdma_0:m_read_readdatavalid
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect        : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata          : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest       : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address           : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read              : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write             : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_beginbursttransfer : std_logic;                     -- mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_beginbursttransfer -> mem_if_lpddr2_emif_0:avl_burstbegin_0
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_readdata           : std_logic_vector(31 downto 0); -- mem_if_lpddr2_emif_0:avl_rdata_0 -> mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_readdata
	signal mem_if_lpddr2_emif_0_avl_0_waitrequest                          : std_logic;                     -- mem_if_lpddr2_emif_0:avl_ready_0 -> mem_if_lpddr2_emif_0_avl_0_waitrequest:in
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_address            : std_logic_vector(26 downto 0); -- mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_address -> mem_if_lpddr2_emif_0:avl_addr_0
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_read               : std_logic;                     -- mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_read -> mem_if_lpddr2_emif_0:avl_read_req_0
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_byteenable -> mem_if_lpddr2_emif_0:avl_be_0
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_readdatavalid      : std_logic;                     -- mem_if_lpddr2_emif_0:avl_rdata_valid_0 -> mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_readdatavalid
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_write              : std_logic;                     -- mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_write -> mem_if_lpddr2_emif_0:avl_write_req_0
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_writedata -> mem_if_lpddr2_emif_0:avl_wdata_0
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_burstcount         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_burstcount -> mem_if_lpddr2_emif_0:avl_size_0
	signal mm_interconnect_0_sysid_control_slave_readdata                  : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                   : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_sgdma_0_csr_chipselect                        : std_logic;                     -- mm_interconnect_0:sgdma_0_csr_chipselect -> sgdma_0:csr_chipselect
	signal mm_interconnect_0_sgdma_0_csr_readdata                          : std_logic_vector(31 downto 0); -- sgdma_0:csr_readdata -> mm_interconnect_0:sgdma_0_csr_readdata
	signal mm_interconnect_0_sgdma_0_csr_address                           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:sgdma_0_csr_address -> sgdma_0:csr_address
	signal mm_interconnect_0_sgdma_0_csr_read                              : std_logic;                     -- mm_interconnect_0:sgdma_0_csr_read -> sgdma_0:csr_read
	signal mm_interconnect_0_sgdma_0_csr_write                             : std_logic;                     -- mm_interconnect_0:sgdma_0_csr_write -> sgdma_0:csr_write
	signal mm_interconnect_0_sgdma_0_csr_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_0_csr_writedata -> sgdma_0:csr_writedata
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                  : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest               : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess               : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                   : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                      : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                     : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_mem_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_chipselect -> onchip_mem:chipselect
	signal mm_interconnect_0_onchip_mem_s1_readdata                        : std_logic_vector(31 downto 0); -- onchip_mem:readdata -> mm_interconnect_0:onchip_mem_s1_readdata
	signal mm_interconnect_0_onchip_mem_s1_address                         : std_logic_vector(12 downto 0); -- mm_interconnect_0:onchip_mem_s1_address -> onchip_mem:address
	signal mm_interconnect_0_onchip_mem_s1_byteenable                      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_mem_s1_byteenable -> onchip_mem:byteenable
	signal mm_interconnect_0_onchip_mem_s1_write                           : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_write -> onchip_mem:write
	signal mm_interconnect_0_onchip_mem_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_mem_s1_writedata -> onchip_mem:writedata
	signal mm_interconnect_0_onchip_mem_s1_clken                           : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_clken -> onchip_mem:clken
	signal mm_interconnect_0_sys_clk_timer_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	signal mm_interconnect_0_sys_clk_timer_s1_readdata                     : std_logic_vector(15 downto 0); -- sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	signal mm_interconnect_0_sys_clk_timer_s1_address                      : std_logic_vector(2 downto 0);  -- mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	signal mm_interconnect_0_sys_clk_timer_s1_write                        : std_logic;                     -- mm_interconnect_0:sys_clk_timer_s1_write -> mm_interconnect_0_sys_clk_timer_s1_write:in
	signal mm_interconnect_0_sys_clk_timer_s1_writedata                    : std_logic_vector(15 downto 0); -- mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	signal mm_interconnect_0_led_pio_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:led_pio_s1_chipselect -> led_pio:chipselect
	signal mm_interconnect_0_led_pio_s1_readdata                           : std_logic_vector(31 downto 0); -- led_pio:readdata -> mm_interconnect_0:led_pio_s1_readdata
	signal mm_interconnect_0_led_pio_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_pio_s1_address -> led_pio:address
	signal mm_interconnect_0_led_pio_s1_write                              : std_logic;                     -- mm_interconnect_0:led_pio_s1_write -> mm_interconnect_0_led_pio_s1_write:in
	signal mm_interconnect_0_led_pio_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_pio_s1_writedata -> led_pio:writedata
	signal mm_interconnect_0_uart_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	signal mm_interconnect_0_uart_s1_readdata                              : std_logic_vector(15 downto 0); -- uart:readdata -> mm_interconnect_0:uart_s1_readdata
	signal mm_interconnect_0_uart_s1_address                               : std_logic_vector(2 downto 0);  -- mm_interconnect_0:uart_s1_address -> uart:address
	signal mm_interconnect_0_uart_s1_read                                  : std_logic;                     -- mm_interconnect_0:uart_s1_read -> mm_interconnect_0_uart_s1_read:in
	signal mm_interconnect_0_uart_s1_begintransfer                         : std_logic;                     -- mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	signal mm_interconnect_0_uart_s1_write                                 : std_logic;                     -- mm_interconnect_0:uart_s1_write -> mm_interconnect_0_uart_s1_write:in
	signal mm_interconnect_0_uart_s1_writedata                             : std_logic_vector(15 downto 0); -- mm_interconnect_0:uart_s1_writedata -> uart:writedata
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                        : std_logic;                     -- sys_clk_timer:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                        : std_logic;                     -- uart:irq -> irq_mapper:receiver3_irq
	signal cpu_irq_irq                                                     : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	signal irq_synchronizer_receiver_irq                                   : std_logic_vector(0 downto 0);  -- sgdma_0:csr_irq -> irq_synchronizer:receiver_irq
	signal sgdma_0_out_valid                                               : std_logic;                     -- sgdma_0:out_valid -> avalon_st_adapter:in_0_valid
	signal sgdma_0_out_data                                                : std_logic_vector(7 downto 0);  -- sgdma_0:out_data -> avalon_st_adapter:in_0_data
	signal sgdma_0_out_ready                                               : std_logic;                     -- avalon_st_adapter:in_0_ready -> sgdma_0:out_ready
	signal sgdma_0_out_startofpacket                                       : std_logic;                     -- sgdma_0:out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	signal sgdma_0_out_endofpacket                                         : std_logic;                     -- sgdma_0:out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	signal avalon_st_adapter_out_0_valid                                   : std_logic;                     -- avalon_st_adapter:out_0_valid -> tx_0:valid
	signal avalon_st_adapter_out_0_data                                    : std_logic_vector(7 downto 0);  -- avalon_st_adapter:out_0_data -> tx_0:data
	signal avalon_st_adapter_out_0_ready                                   : std_logic;                     -- tx_0:ready -> avalon_st_adapter:out_0_ready
	signal avalon_st_adapter_out_0_startofpacket                           : std_logic;                     -- avalon_st_adapter:out_0_startofpacket -> tx_0:startofpacket
	signal avalon_st_adapter_out_0_endofpacket                             : std_logic;                     -- avalon_st_adapter:out_0_endofpacket -> tx_0:endofpacket
	signal avalon_st_adapter_out_0_error                                   : std_logic_vector(0 downto 0);  -- avalon_st_adapter:out_0_error -> tx_0:error
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, onchip_mem:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [cpu:reset_req, onchip_mem:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                              : std_logic;                     -- rst_controller_001:reset_out -> [avalon_st_adapter:in_rst_0_reset, irq_synchronizer:receiver_reset, mm_interconnect_0:sgdma_0_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_002_reset_out_reset                              : std_logic;                     -- rst_controller_002:reset_out -> tx_0:reset
	signal rst_controller_003_reset_out_reset                              : std_logic;                     -- rst_controller_003:reset_out -> [mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:mem_if_lpddr2_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset_reset]
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv    : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv   : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_inv                : std_logic;                     -- mem_if_lpddr2_emif_0_avl_0_waitrequest:inv -> mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_waitrequest
	signal mm_interconnect_0_sys_clk_timer_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_sys_clk_timer_s1_write:inv -> sys_clk_timer:write_n
	signal mm_interconnect_0_led_pio_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_led_pio_s1_write:inv -> led_pio:write_n
	signal mm_interconnect_0_uart_s1_read_ports_inv                        : std_logic;                     -- mm_interconnect_0_uart_s1_read:inv -> uart:read_n
	signal mm_interconnect_0_uart_s1_write_ports_inv                       : std_logic;                     -- mm_interconnect_0_uart_s1_write:inv -> uart:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [cpu:reset_n, jtag_uart:rst_n, led_pio:reset_n, sys_clk_timer:reset_n, sysid:reset_n, uart:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> sgdma_0:system_reset_n

begin

	cpu : component system_cpu
		port map (
			clk                                 => clk_clk,                                           --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                              --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	jtag_uart : component system_jtag_uart
		port map (
			clk            => clk_clk,                                                       --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                       --               irq.irq
		);

	led_pio : component system_led_pio
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_led_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_pio_s1_readdata,        --                    .readdata
			out_port   => led_pio_external_connection_export            -- external_connection.export
		);

	mem_if_lpddr2_emif_0 : component system_mem_if_lpddr2_emif_0
		port map (
			pll_ref_clk                => mem_if_lpddr2_emif_0_pll_ref_clk_clk,                            --        pll_ref_clk.clk
			global_reset_n             => reset_reset_n,                                                   --       global_reset.reset_n
			soft_reset_n               => reset_reset_n,                                                   --         soft_reset.reset_n
			afi_clk                    => open,                                                            --            afi_clk.clk
			afi_half_clk               => mem_if_lpddr2_emif_0_afi_half_clk_clk,                           --       afi_half_clk.clk
			afi_reset_n                => open,                                                            --          afi_reset.reset_n
			afi_reset_export_n         => open,                                                            --   afi_reset_export.reset_n
			mem_ca                     => memory_mem_ca,                                                   --             memory.mem_ca
			mem_ck                     => memory_mem_ck,                                                   --                   .mem_ck
			mem_ck_n                   => memory_mem_ck_n,                                                 --                   .mem_ck_n
			mem_cke                    => memory_mem_cke,                                                  --                   .mem_cke
			mem_cs_n                   => memory_mem_cs_n,                                                 --                   .mem_cs_n
			mem_dm                     => memory_mem_dm,                                                   --                   .mem_dm
			mem_dq                     => memory_mem_dq,                                                   --                   .mem_dq
			mem_dqs                    => memory_mem_dqs,                                                  --                   .mem_dqs
			mem_dqs_n                  => memory_mem_dqs_n,                                                --                   .mem_dqs_n
			avl_ready_0                => mem_if_lpddr2_emif_0_avl_0_waitrequest,                          --              avl_0.waitrequest_n
			avl_burstbegin_0           => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_beginbursttransfer, --                   .beginbursttransfer
			avl_addr_0                 => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_address,            --                   .address
			avl_rdata_valid_0          => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_readdatavalid,      --                   .readdatavalid
			avl_rdata_0                => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_readdata,           --                   .readdata
			avl_wdata_0                => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_writedata,          --                   .writedata
			avl_be_0                   => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_byteenable,         --                   .byteenable
			avl_read_req_0             => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_read,               --                   .read
			avl_write_req_0            => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_write,              --                   .write
			avl_size_0                 => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_burstcount,         --                   .burstcount
			mp_cmd_clk_0_clk           => mem_if_lpddr2_emif_0_afi_half_clk_clk,                           --       mp_cmd_clk_0.clk
			mp_cmd_reset_n_0_reset_n   => reset_reset_n,                                                   --   mp_cmd_reset_n_0.reset_n
			mp_rfifo_clk_0_clk         => mem_if_lpddr2_emif_0_afi_half_clk_clk,                           --     mp_rfifo_clk_0.clk
			mp_rfifo_reset_n_0_reset_n => reset_reset_n,                                                   -- mp_rfifo_reset_n_0.reset_n
			mp_wfifo_clk_0_clk         => mem_if_lpddr2_emif_0_afi_half_clk_clk,                           --     mp_wfifo_clk_0.clk
			mp_wfifo_reset_n_0_reset_n => reset_reset_n,                                                   -- mp_wfifo_reset_n_0.reset_n
			local_init_done            => mem_if_lpddr2_emif_0_status_local_init_done,                     --             status.local_init_done
			local_cal_success          => mem_if_lpddr2_emif_0_status_local_cal_success,                   --                   .local_cal_success
			local_cal_fail             => mem_if_lpddr2_emif_0_status_local_cal_fail,                      --                   .local_cal_fail
			oct_rzqin                  => oct_rzqin,                                                       --                oct.rzqin
			pll_mem_clk                => mem_if_lpddr2_emif_0_pll_sharing_pll_mem_clk,                    --        pll_sharing.pll_mem_clk
			pll_write_clk              => mem_if_lpddr2_emif_0_pll_sharing_pll_write_clk,                  --                   .pll_write_clk
			pll_locked                 => mem_if_lpddr2_emif_0_pll_sharing_pll_locked,                     --                   .pll_locked
			pll_write_clk_pre_phy_clk  => mem_if_lpddr2_emif_0_pll_sharing_pll_write_clk_pre_phy_clk,      --                   .pll_write_clk_pre_phy_clk
			pll_addr_cmd_clk           => mem_if_lpddr2_emif_0_pll_sharing_pll_addr_cmd_clk,               --                   .pll_addr_cmd_clk
			pll_avl_clk                => mem_if_lpddr2_emif_0_pll_sharing_pll_avl_clk,                    --                   .pll_avl_clk
			pll_config_clk             => mem_if_lpddr2_emif_0_pll_sharing_pll_config_clk,                 --                   .pll_config_clk
			pll_mem_phy_clk            => mem_if_lpddr2_emif_0_pll_sharing_pll_mem_phy_clk,                --                   .pll_mem_phy_clk
			afi_phy_clk                => mem_if_lpddr2_emif_0_pll_sharing_afi_phy_clk,                    --                   .afi_phy_clk
			pll_avl_phy_clk            => mem_if_lpddr2_emif_0_pll_sharing_pll_avl_phy_clk                 --                   .pll_avl_phy_clk
		);

	onchip_mem : component system_onchip_mem
		port map (
			clk        => clk_clk,                                    --   clk1.clk
			address    => mm_interconnect_0_onchip_mem_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_mem_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_mem_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_mem_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_mem_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_mem_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_mem_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req          --       .reset_req
		);

	sgdma_0 : component system_sgdma_0
		port map (
			clk                           => clk_hsmc_clk,                                 --              clk.clk
			system_reset_n                => rst_controller_001_reset_out_reset_ports_inv, --            reset.reset_n
			csr_chipselect                => mm_interconnect_0_sgdma_0_csr_chipselect,     --              csr.chipselect
			csr_address                   => mm_interconnect_0_sgdma_0_csr_address,        --                 .address
			csr_read                      => mm_interconnect_0_sgdma_0_csr_read,           --                 .read
			csr_write                     => mm_interconnect_0_sgdma_0_csr_write,          --                 .write
			csr_writedata                 => mm_interconnect_0_sgdma_0_csr_writedata,      --                 .writedata
			csr_readdata                  => mm_interconnect_0_sgdma_0_csr_readdata,       --                 .readdata
			descriptor_read_readdata      => sgdma_0_descriptor_read_readdata,             --  descriptor_read.readdata
			descriptor_read_readdatavalid => sgdma_0_descriptor_read_readdatavalid,        --                 .readdatavalid
			descriptor_read_waitrequest   => sgdma_0_descriptor_read_waitrequest,          --                 .waitrequest
			descriptor_read_address       => sgdma_0_descriptor_read_address,              --                 .address
			descriptor_read_read          => sgdma_0_descriptor_read_read,                 --                 .read
			descriptor_write_waitrequest  => sgdma_0_descriptor_write_waitrequest,         -- descriptor_write.waitrequest
			descriptor_write_address      => sgdma_0_descriptor_write_address,             --                 .address
			descriptor_write_write        => sgdma_0_descriptor_write_write,               --                 .write
			descriptor_write_writedata    => sgdma_0_descriptor_write_writedata,           --                 .writedata
			csr_irq                       => irq_synchronizer_receiver_irq(0),             --          csr_irq.irq
			m_read_readdata               => sgdma_0_m_read_readdata,                      --           m_read.readdata
			m_read_readdatavalid          => sgdma_0_m_read_readdatavalid,                 --                 .readdatavalid
			m_read_waitrequest            => sgdma_0_m_read_waitrequest,                   --                 .waitrequest
			m_read_address                => sgdma_0_m_read_address,                       --                 .address
			m_read_read                   => sgdma_0_m_read_read,                          --                 .read
			out_data                      => sgdma_0_out_data,                             --              out.data
			out_valid                     => sgdma_0_out_valid,                            --                 .valid
			out_ready                     => sgdma_0_out_ready,                            --                 .ready
			out_endofpacket               => sgdma_0_out_endofpacket,                      --                 .endofpacket
			out_startofpacket             => sgdma_0_out_startofpacket                     --                 .startofpacket
		);

	sys_clk_timer : component system_sys_clk_timer
		port map (
			clk        => clk_clk,                                            --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           -- reset.reset_n
			address    => mm_interconnect_0_sys_clk_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_sys_clk_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_sys_clk_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_sys_clk_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_sys_clk_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver2_irq                            --   irq.irq
		);

	sysid : component system_sysid
		port map (
			clock    => clk_clk,                                          --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	tx_0 : component tx
		port map (
			clk            => clk_hsmc_clk,                          --                   clock.clk
			reset          => rst_controller_002_reset_out_reset,    --                   reset.reset
			tx_serial_data => tx_0_tx_serial_data_serial_data,       --          tx_serial_data.serial_data
			data           => avalon_st_adapter_out_0_data,          -- avalon_streaming_sink_1.data
			error          => avalon_st_adapter_out_0_error(0),      --                        .error
			ready          => avalon_st_adapter_out_0_ready,         --                        .ready
			valid          => avalon_st_adapter_out_0_valid,         --                        .valid
			startofpacket  => avalon_st_adapter_out_0_startofpacket, --                        .startofpacket
			endofpacket    => avalon_st_adapter_out_0_endofpacket,   --                        .endofpacket
			led            => tx_0_led_readdata                      --                     led.readdata
		);

	uart : component system_uart
		port map (
			clk           => clk_clk,                                   --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address       => mm_interconnect_0_uart_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_uart_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_uart_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_uart_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_uart_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_uart_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_uart_s1_readdata,        --                    .readdata
			dataavailable => open,                                      --                    .dataavailable
			readyfordata  => open,                                      --                    .readyfordata
			rxd           => uart_external_connection_rxd,              -- external_connection.export
			txd           => uart_external_connection_txd,              --                    .export
			irq           => irq_mapper_receiver3_irq                   --                 irq.irq
		);

	mm_interconnect_0 : component system_mm_interconnect_0
		port map (
			clk_0_clk_clk                                                           => clk_clk,                                                         --                                                         clk_0_clk.clk
			clk_hsmc_clk_clk                                                        => clk_hsmc_clk,                                                    --                                                      clk_hsmc_clk.clk
			mem_if_lpddr2_emif_0_afi_half_clk_clk                                   => mem_if_lpddr2_emif_0_afi_half_clk_clk,                           --                                 mem_if_lpddr2_emif_0_afi_half_clk.clk
			cpu_reset_reset_bridge_in_reset_reset                                   => rst_controller_reset_out_reset,                                  --                                   cpu_reset_reset_bridge_in_reset.reset
			mem_if_lpddr2_emif_0_avl_0_translator_reset_reset_bridge_in_reset_reset => rst_controller_003_reset_out_reset,                              -- mem_if_lpddr2_emif_0_avl_0_translator_reset_reset_bridge_in_reset.reset
			mem_if_lpddr2_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset_reset       => rst_controller_003_reset_out_reset,                              --       mem_if_lpddr2_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset.reset
			sgdma_0_reset_reset_bridge_in_reset_reset                               => rst_controller_001_reset_out_reset,                              --                               sgdma_0_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                                                 => cpu_data_master_address,                                         --                                                   cpu_data_master.address
			cpu_data_master_waitrequest                                             => cpu_data_master_waitrequest,                                     --                                                                  .waitrequest
			cpu_data_master_byteenable                                              => cpu_data_master_byteenable,                                      --                                                                  .byteenable
			cpu_data_master_read                                                    => cpu_data_master_read,                                            --                                                                  .read
			cpu_data_master_readdata                                                => cpu_data_master_readdata,                                        --                                                                  .readdata
			cpu_data_master_write                                                   => cpu_data_master_write,                                           --                                                                  .write
			cpu_data_master_writedata                                               => cpu_data_master_writedata,                                       --                                                                  .writedata
			cpu_data_master_debugaccess                                             => cpu_data_master_debugaccess,                                     --                                                                  .debugaccess
			cpu_instruction_master_address                                          => cpu_instruction_master_address,                                  --                                            cpu_instruction_master.address
			cpu_instruction_master_waitrequest                                      => cpu_instruction_master_waitrequest,                              --                                                                  .waitrequest
			cpu_instruction_master_read                                             => cpu_instruction_master_read,                                     --                                                                  .read
			cpu_instruction_master_readdata                                         => cpu_instruction_master_readdata,                                 --                                                                  .readdata
			cpu_instruction_master_readdatavalid                                    => cpu_instruction_master_readdatavalid,                            --                                                                  .readdatavalid
			sgdma_0_descriptor_read_address                                         => sgdma_0_descriptor_read_address,                                 --                                           sgdma_0_descriptor_read.address
			sgdma_0_descriptor_read_waitrequest                                     => sgdma_0_descriptor_read_waitrequest,                             --                                                                  .waitrequest
			sgdma_0_descriptor_read_read                                            => sgdma_0_descriptor_read_read,                                    --                                                                  .read
			sgdma_0_descriptor_read_readdata                                        => sgdma_0_descriptor_read_readdata,                                --                                                                  .readdata
			sgdma_0_descriptor_read_readdatavalid                                   => sgdma_0_descriptor_read_readdatavalid,                           --                                                                  .readdatavalid
			sgdma_0_descriptor_write_address                                        => sgdma_0_descriptor_write_address,                                --                                          sgdma_0_descriptor_write.address
			sgdma_0_descriptor_write_waitrequest                                    => sgdma_0_descriptor_write_waitrequest,                            --                                                                  .waitrequest
			sgdma_0_descriptor_write_write                                          => sgdma_0_descriptor_write_write,                                  --                                                                  .write
			sgdma_0_descriptor_write_writedata                                      => sgdma_0_descriptor_write_writedata,                              --                                                                  .writedata
			sgdma_0_m_read_address                                                  => sgdma_0_m_read_address,                                          --                                                    sgdma_0_m_read.address
			sgdma_0_m_read_waitrequest                                              => sgdma_0_m_read_waitrequest,                                      --                                                                  .waitrequest
			sgdma_0_m_read_read                                                     => sgdma_0_m_read_read,                                             --                                                                  .read
			sgdma_0_m_read_readdata                                                 => sgdma_0_m_read_readdata,                                         --                                                                  .readdata
			sgdma_0_m_read_readdatavalid                                            => sgdma_0_m_read_readdatavalid,                                    --                                                                  .readdatavalid
			cpu_debug_mem_slave_address                                             => mm_interconnect_0_cpu_debug_mem_slave_address,                   --                                               cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write                                               => mm_interconnect_0_cpu_debug_mem_slave_write,                     --                                                                  .write
			cpu_debug_mem_slave_read                                                => mm_interconnect_0_cpu_debug_mem_slave_read,                      --                                                                  .read
			cpu_debug_mem_slave_readdata                                            => mm_interconnect_0_cpu_debug_mem_slave_readdata,                  --                                                                  .readdata
			cpu_debug_mem_slave_writedata                                           => mm_interconnect_0_cpu_debug_mem_slave_writedata,                 --                                                                  .writedata
			cpu_debug_mem_slave_byteenable                                          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,                --                                                                  .byteenable
			cpu_debug_mem_slave_waitrequest                                         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,               --                                                                  .waitrequest
			cpu_debug_mem_slave_debugaccess                                         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,               --                                                                  .debugaccess
			jtag_uart_avalon_jtag_slave_address                                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,           --                                       jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                                       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,             --                                                                  .write
			jtag_uart_avalon_jtag_slave_read                                        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,              --                                                                  .read
			jtag_uart_avalon_jtag_slave_readdata                                    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,          --                                                                  .readdata
			jtag_uart_avalon_jtag_slave_writedata                                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,         --                                                                  .writedata
			jtag_uart_avalon_jtag_slave_waitrequest                                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,       --                                                                  .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                                  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,        --                                                                  .chipselect
			led_pio_s1_address                                                      => mm_interconnect_0_led_pio_s1_address,                            --                                                        led_pio_s1.address
			led_pio_s1_write                                                        => mm_interconnect_0_led_pio_s1_write,                              --                                                                  .write
			led_pio_s1_readdata                                                     => mm_interconnect_0_led_pio_s1_readdata,                           --                                                                  .readdata
			led_pio_s1_writedata                                                    => mm_interconnect_0_led_pio_s1_writedata,                          --                                                                  .writedata
			led_pio_s1_chipselect                                                   => mm_interconnect_0_led_pio_s1_chipselect,                         --                                                                  .chipselect
			mem_if_lpddr2_emif_0_avl_0_address                                      => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_address,            --                                        mem_if_lpddr2_emif_0_avl_0.address
			mem_if_lpddr2_emif_0_avl_0_write                                        => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_write,              --                                                                  .write
			mem_if_lpddr2_emif_0_avl_0_read                                         => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_read,               --                                                                  .read
			mem_if_lpddr2_emif_0_avl_0_readdata                                     => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_readdata,           --                                                                  .readdata
			mem_if_lpddr2_emif_0_avl_0_writedata                                    => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_writedata,          --                                                                  .writedata
			mem_if_lpddr2_emif_0_avl_0_beginbursttransfer                           => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_beginbursttransfer, --                                                                  .beginbursttransfer
			mem_if_lpddr2_emif_0_avl_0_burstcount                                   => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_burstcount,         --                                                                  .burstcount
			mem_if_lpddr2_emif_0_avl_0_byteenable                                   => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_byteenable,         --                                                                  .byteenable
			mem_if_lpddr2_emif_0_avl_0_readdatavalid                                => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_readdatavalid,      --                                                                  .readdatavalid
			mem_if_lpddr2_emif_0_avl_0_waitrequest                                  => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_inv,                --                                                                  .waitrequest
			onchip_mem_s1_address                                                   => mm_interconnect_0_onchip_mem_s1_address,                         --                                                     onchip_mem_s1.address
			onchip_mem_s1_write                                                     => mm_interconnect_0_onchip_mem_s1_write,                           --                                                                  .write
			onchip_mem_s1_readdata                                                  => mm_interconnect_0_onchip_mem_s1_readdata,                        --                                                                  .readdata
			onchip_mem_s1_writedata                                                 => mm_interconnect_0_onchip_mem_s1_writedata,                       --                                                                  .writedata
			onchip_mem_s1_byteenable                                                => mm_interconnect_0_onchip_mem_s1_byteenable,                      --                                                                  .byteenable
			onchip_mem_s1_chipselect                                                => mm_interconnect_0_onchip_mem_s1_chipselect,                      --                                                                  .chipselect
			onchip_mem_s1_clken                                                     => mm_interconnect_0_onchip_mem_s1_clken,                           --                                                                  .clken
			sgdma_0_csr_address                                                     => mm_interconnect_0_sgdma_0_csr_address,                           --                                                       sgdma_0_csr.address
			sgdma_0_csr_write                                                       => mm_interconnect_0_sgdma_0_csr_write,                             --                                                                  .write
			sgdma_0_csr_read                                                        => mm_interconnect_0_sgdma_0_csr_read,                              --                                                                  .read
			sgdma_0_csr_readdata                                                    => mm_interconnect_0_sgdma_0_csr_readdata,                          --                                                                  .readdata
			sgdma_0_csr_writedata                                                   => mm_interconnect_0_sgdma_0_csr_writedata,                         --                                                                  .writedata
			sgdma_0_csr_chipselect                                                  => mm_interconnect_0_sgdma_0_csr_chipselect,                        --                                                                  .chipselect
			sys_clk_timer_s1_address                                                => mm_interconnect_0_sys_clk_timer_s1_address,                      --                                                  sys_clk_timer_s1.address
			sys_clk_timer_s1_write                                                  => mm_interconnect_0_sys_clk_timer_s1_write,                        --                                                                  .write
			sys_clk_timer_s1_readdata                                               => mm_interconnect_0_sys_clk_timer_s1_readdata,                     --                                                                  .readdata
			sys_clk_timer_s1_writedata                                              => mm_interconnect_0_sys_clk_timer_s1_writedata,                    --                                                                  .writedata
			sys_clk_timer_s1_chipselect                                             => mm_interconnect_0_sys_clk_timer_s1_chipselect,                   --                                                                  .chipselect
			sysid_control_slave_address                                             => mm_interconnect_0_sysid_control_slave_address,                   --                                               sysid_control_slave.address
			sysid_control_slave_readdata                                            => mm_interconnect_0_sysid_control_slave_readdata,                  --                                                                  .readdata
			uart_s1_address                                                         => mm_interconnect_0_uart_s1_address,                               --                                                           uart_s1.address
			uart_s1_write                                                           => mm_interconnect_0_uart_s1_write,                                 --                                                                  .write
			uart_s1_read                                                            => mm_interconnect_0_uart_s1_read,                                  --                                                                  .read
			uart_s1_readdata                                                        => mm_interconnect_0_uart_s1_readdata,                              --                                                                  .readdata
			uart_s1_writedata                                                       => mm_interconnect_0_uart_s1_writedata,                             --                                                                  .writedata
			uart_s1_begintransfer                                                   => mm_interconnect_0_uart_s1_begintransfer,                         --                                                                  .begintransfer
			uart_s1_chipselect                                                      => mm_interconnect_0_uart_s1_chipselect                             --                                                                  .chipselect
		);

	irq_mapper : component system_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk_hsmc_clk,                       --       receiver_clk.clk
			sender_clk     => clk_clk,                            --         sender_clk.clk
			receiver_reset => rst_controller_001_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_reset_out_reset,     --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver0_irq            --             sender.irq
		);

	avalon_st_adapter : component system_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 8,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 8,
			outChannelWidth => 0,
			outErrorWidth   => 1,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => clk_hsmc_clk,                          -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_001_reset_out_reset,    -- in_rst_0.reset
			in_0_data           => sgdma_0_out_data,                      --     in_0.data
			in_0_valid          => sgdma_0_out_valid,                     --         .valid
			in_0_ready          => sgdma_0_out_ready,                     --         .ready
			in_0_startofpacket  => sgdma_0_out_startofpacket,             --         .startofpacket
			in_0_endofpacket    => sgdma_0_out_endofpacket,               --         .endofpacket
			out_0_data          => avalon_st_adapter_out_0_data,          --    out_0.data
			out_0_valid         => avalon_st_adapter_out_0_valid,         --         .valid
			out_0_ready         => avalon_st_adapter_out_0_ready,         --         .ready
			out_0_startofpacket => avalon_st_adapter_out_0_startofpacket, --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_out_0_endofpacket,   --         .endofpacket
			out_0_error         => avalon_st_adapter_out_0_error          --         .error
		);

	rst_controller : component system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_hsmc_clk,                       --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_hsmc_clk,                       --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_003 : component system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,               -- reset_in0.reset
			clk            => mem_if_lpddr2_emif_0_afi_half_clk_clk, --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset,    -- reset_out.reset
			reset_req      => open,                                  -- (terminated)
			reset_req_in0  => '0',                                   -- (terminated)
			reset_in1      => '0',                                   -- (terminated)
			reset_req_in1  => '0',                                   -- (terminated)
			reset_in2      => '0',                                   -- (terminated)
			reset_req_in2  => '0',                                   -- (terminated)
			reset_in3      => '0',                                   -- (terminated)
			reset_req_in3  => '0',                                   -- (terminated)
			reset_in4      => '0',                                   -- (terminated)
			reset_req_in4  => '0',                                   -- (terminated)
			reset_in5      => '0',                                   -- (terminated)
			reset_req_in5  => '0',                                   -- (terminated)
			reset_in6      => '0',                                   -- (terminated)
			reset_req_in6  => '0',                                   -- (terminated)
			reset_in7      => '0',                                   -- (terminated)
			reset_req_in7  => '0',                                   -- (terminated)
			reset_in8      => '0',                                   -- (terminated)
			reset_req_in8  => '0',                                   -- (terminated)
			reset_in9      => '0',                                   -- (terminated)
			reset_req_in9  => '0',                                   -- (terminated)
			reset_in10     => '0',                                   -- (terminated)
			reset_req_in10 => '0',                                   -- (terminated)
			reset_in11     => '0',                                   -- (terminated)
			reset_req_in11 => '0',                                   -- (terminated)
			reset_in12     => '0',                                   -- (terminated)
			reset_req_in12 => '0',                                   -- (terminated)
			reset_in13     => '0',                                   -- (terminated)
			reset_req_in13 => '0',                                   -- (terminated)
			reset_in14     => '0',                                   -- (terminated)
			reset_req_in14 => '0',                                   -- (terminated)
			reset_in15     => '0',                                   -- (terminated)
			reset_req_in15 => '0'                                    -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_inv <= not mem_if_lpddr2_emif_0_avl_0_waitrequest;

	mm_interconnect_0_sys_clk_timer_s1_write_ports_inv <= not mm_interconnect_0_sys_clk_timer_s1_write;

	mm_interconnect_0_led_pio_s1_write_ports_inv <= not mm_interconnect_0_led_pio_s1_write;

	mm_interconnect_0_uart_s1_read_ports_inv <= not mm_interconnect_0_uart_s1_read;

	mm_interconnect_0_uart_s1_write_ports_inv <= not mm_interconnect_0_uart_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of system
