// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:40 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bmis7y5PviwZtNjbtgfB5xc4H55S5qRheCU2R6X+6ADN51+3V787KaOg4chpocu8
02wbqyipF1EEVT6MBhTQzgPO6+Q7lyYfG1Qe4ZCdCzXaBj13sjbmDkbt9A4guAwt
5GLDlGBfuf1GVhJDQtvGGOWxTu5uVeZgoTkao2k2UJA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6416)
GeJ72GbCIhb7tekql1OASHxnwH9lPEUZHhI9C336F1B+0eUqVOzC3hbz0m3WNXOk
zkTBHyRMYT7vpG6AqcHMKq1j6ZzefGgVbndU3ni/azaBcTEpr+ZG6a/I1ozI+PGX
Vsf1iOVqSfKsbeO5j+wjnk2+tDlQ370t6bucbe0oi+qUKcfSC4nNW+cSv58IZFPS
g2Foo6YY8595fB/eBz7if6Vgxea84tAW8hpioy3G2iVxABDVu5QPcPnZhS3ZnNTM
sFvPfyDJvN4HXs8li7DrHBPtO5p+zMBVlY415Jo5/w1gBFUTWQYR0QHkQHzJZKt+
GkdzYO1+dWMcwtKR27eHlKRR9mHVkazZh7iIm33kujYR8i5g/XWlFrFMq0jWZLRs
zmEwzAHcY0Fe0AiuIlxEq3wwrPrdTDMPUX4axtqSO7t0oRv+jJa7yz7zrTmyQSfY
sQHqSfwhqI/nrPyyJnkgowloVA88yGG3TmvfTLo8o+Q6pYIGlJptelwkIuiMrIJL
3wTnSJXj44LFEv9WlNGHDzEKznZvSwzpd/6vFFDHpVnEHbhFzLWZp8d8Ca2bBDcp
uLRBq4fFgdMltkd2X8aSuD2nauSV1bePhpqEng0L6bEGbJvPKecW5fCfvnUpGEYG
CkgbYENxKoFvzCLYNRTz/6ohHSblBAAyMOPXM3Yg+RYmfJr/D0orsSDBkVLWfDtp
okzjK6IlA2QjyfbnAX4hd5Y349dNlUls54Ij+rV9ANvOrN1waql3yWentgx+B6ko
SN7XP+JSjCJWaqp+++iYndaz6WqfeYslGcKEl0CD/keEI19q6W6moHl2daTaInQC
sg1wfBO9PolUEAf6j6piL4OsXLsi/k4TmHUHtEpQaFjQ6tcY/MkY/6+OjB8Q37FJ
14giAtuqwDsmBOFfqeAMkGBBS0sUrguIBqwA25PePuxNRpU+pt4AbNhMNU0WHdNw
aRKaS6GKxSOxRPXKWn9U2zO9lSb0xrMXd4Cy3S7TkO3cYiRBUBuXw4O8GKSoawDN
ocZAdrtQQk9zQLp9CYrVrUMIDNUK/UZQw9AtZMIIF4WGy1Hdv9lz2BEs/CCQl9K+
6E15nicJuWa/NwlMEFQ/9caBHRpOE1WyovuyAyjyNKiFEe6ZKXXZ53VJh7V64e1C
VfwuJEk8CAWuaVf+bS1/ES/g7KSXNtt4mR6do7qsJFBd/28WBYDpGDcjkp0z+OV5
eUyWcGM7cSZJlxAPD4hSrFnvvDl8oTTwA6HqDNeaRlYsf9N/XGO+w2+KxeFd0yxU
x8rGBw8Ca3TlmuE33ZFa+cLusOgvijL+yJZ57QyxdOmMF+1ru9+MdboY6PuoaYgs
kDvYnlj/j9fW0URgyyYZZ1yfZgPHsaqOnfT5mIjtszAztzRK9eSoJTv/hFn1whGP
OjT68nG0N2xtd5ecpS+cpIOD6ZRL+3yADcgXBEEH0U1GbEuqtaEI9r4PCHPHUn3o
hl6F/DbpOHh/Eld6WIUiyFuV/weOXaWZ7JPyiA21mnXUBG0zuDWgp4+wX1ECM0pd
kcBiRnBhh/Co6Wb3+a9Hlk7phdRVhO9mz+d23FPcB+YC66rJ5BwJ+Sb2aAy5aA6J
jM54GKC4DBr2M2exGwE5fqo85SwgyApKVbcckb/APlsoiYy6/udyLDUK0Ua1LsSR
5jDG6mn+RPbBWcI/MPG16TN2mWJ+Mi5RtOBOrI+1ArFBvPRiKUCQdVv5748NvAtc
V7QjcP9JqAVJUc6clZGv3Sf6018Zq7tMxbzhlGfbpWqjGvvXl9Vk9d2FCgQ9Mr4i
D0PIS0lsyO82jiv626pbi4up9AVJJ5EX03E7Q0LzxZfRITVcvndxwPSygunDzToK
4Tzue/FDZYe9qPL8eFGNAt168f8igd5BZFtybrr+yMkO6OsrRXyK1sDRFUYXwsgI
g3MJK+Z7J6NAXGFcVzkYs/QHXH7iH7p/E4w3ZEIfNYYBffXQn0/4P3PcJOT074BN
TIPcxPzvt5KgmPUg0osZnxTxVh3QG1ZPRx7z8gsUsmZOCLeo6WMvTrthO17QTjD9
opQzqdOief2E14YomGxySes73SGby3R4Q2dce3apoRvTZ9FQGPHeloKEMGrZ7ciE
FTSjZsKHG6k+b3vxOjSj3w70UgU528By5W4X0SEWEEVx/cIg/aH+Nslw6a0CxDMl
Uijq7piAo+MgcGan0NOpBvE+oqP3otFULGHF4zsI5X0atbsa7vNQij7iBWxd3fde
JYt1WqllcdsRlBpk2v43ssdTUvUDEd+a0V945Wp29UcLeUmOqZWeAQvmxW+sTBuU
MQSjuEFmZFc0SL/5KgxGte0xEGfwNa1IL4KP1T5ti6R7xgjZXAqgialHcE5fRReI
MHTfh8Vcv55eYSvYIGu2ephDGebdowjcnAZ+PJrTr7rVa7/illCC6d+EzcWqthFe
SSvcRiXbJwOehgdUaJXJUc82CEbd0VJeTN4kQWqdc+2ilDAM4P+ZMC1DX+XhEeqx
xp7Tc7ysXoXDMulOFOc5aswIhsiywOFJX2FOnRXtSrb/xW0VTugIhnuHeXBSl1ek
RSWqO8emX/FAjLHmsxG2/0RDG1h3fYYAM3h2Q1tKmgd1+c75mO34QJXCKpdvMwAZ
JRjBUtTaCJx8fQT5QpEt6kVSRidSwPFhqQ8Lbs31BwGjSqH1VDsDkfIjSIXCV+wV
2r26AtRpDcZagZ/HC6M1I3za7sTMZfD0CjOJzURofuNGYUVOpI7gZyCOLv07huVh
jeaP6noiVuGWyj/WiPDaAO6azsNY5Y8LtRAIk+KvpxoRYE7N0oVFNv8WB+QI9C1i
TcaQC8HtJIVRZfQ/uGn0StWU2Ztmon+en49AG/++2cUjMeEvzfAAe0ritKi+vG4h
XTJLwJ4hLo2Wf3VJC1dFA8tjQ8D5ZTMjB0AAaW8Ow1OB5LMtIqbqgw1dY0TFLy5f
IP7v0mqFeY5eS77rgw9BM9mXnuW3Al8hlh4+CtzJwrFHKmB9MfDDXxBOTXiyxRIV
eXrA/0OwctHQdV8N6+RWbJqnPM53kjUNwewIl/PNao6o1yvaiCrYf5CKtBHibQ9a
MFECNlaftIUs7NfSngoVWpIVODD4AIz6eLnFHmfSJ2jGqrIP3/NsSh8VMz2+58kQ
faBmMYNlZHa/p0G4X0KHcGwSjUSTch24ro1Y4+5hLKN6fu8hcosuuHU/mdkmhhys
OuElSBuAlbgD/Tamb28rnupqnEV6JxAB3CtABSNuklW5tFEbRfmkWAQ8KppssDb9
eynWwozdNeM4G3IuyIm5OXESThUVHaRGZV7e9IqdJ6YeZQJcTRHhlOKWwWi+yXwA
puYOzexSWGaLfGavlt4xiCdza+9oLyE+P4KkqMigcN7+r/BNVc/S0bfQimT1uLOL
XnnGPSYZzTur+IzWOuKrpwS2jRTU9490ZMran+6eRNjRT1aOJeElpVWtB/f39Lbs
ustZhpnXtYEXecety/Sw7JQW5kvDH+uE+9QMxEafrDx3e1Qjw7wJOcYC4WT06KXz
5nyyN477B+3vm/uR6Op7XjtoCrpY+cCzEuA2fF/Zr6sWBBrcZxGk7rMEsvxS6WIP
PULVvsLJzKvsikkYV+fHBd4vLc2kPe9d6BxSAZixAZaOYnaB47V+XTYq9TnkrfBA
EZ4ej1dgdvTihPZ7ZGWYGawVV6qz4IJckYtugy5iyXYQ9/6YdN7Bu4Ry0yvJQJrv
UK+59frq3W0TgUygR2i3lcLd+qvds7y266YV/TiYovVauJMH7n7Qf5jUiO8lug5l
PA/QcJrs+1lOTrNVDiqw9UzS0U0aIxUDke1G8b8jFlrNsPI4nGwYmlw8ofJH+dib
7GeXecqpx8B7gWLI+vN7Y3tpUMgaJJjUizvH9YqMSGcgqnkoHBsKxJOzo4R6wdRW
7CxyF6qCOY2tVO86Q4XJmt936vUI4+qdM962e9Cekw2ICnSiwti7yqegz3jyInGv
1ubGaPzxlMgYcGZb7tTRTAy/myXpW3TzshdbjSWfgbPZq7PeGg9szIwQd0lgjP+V
vrPB0+o1nOrotho+LsyBRQR/pbhwoDvN4t0YOOgqhtsntG4wDxBCkakKMlZbCsVJ
NNDzjpnDP6KGF9mzVJHnFDEDJZikY09N/UjWveh2R4+aT7TpoOK3hhtubmon7Wrr
xQqFYOw6IpsmfVh+sYLRvOKB6dXcQeVtLhk005kItHnyP11Clkjji1JydUYYH8Kh
S919FAa1nFvvByMUfSi0UuvTaL6em18Vt2xJn1ikRHvT7THjuOJSnVtrSOW1+oTS
x6nibQAyUJtEMyl268Ky1JRcGs9EYvc3WchcPJx9eAv9LlQJoGM8iZOzC3p71g5V
ZvmSjPfAfzVWDlhCVqI4OBba1fC5a3f977+djNEpWpHcauummnORHbG/gf/zCiGz
T+p1U/PxdQqVyfPuxvN9ulhvUQErk7DnwN4AJEvGfWuACTx/QiM9un2Kia7E9PDx
AzRoUjDpaDaAkFxaglpvCP68N4dExGpo1ngtR2T2A62M76HwZvlOW6BNQCPd223f
L7n4oSA8ORrS737sajG2UzNsXZX02jjWAzX2FEUwQKac25kruHUPp7J0I876hyCX
+9JWJi4gkwiDDRIP4ebi7PB+cXq0p7HiyTvzR6VR98MysqNmZtmAxRD+GgHdwEBM
XyAgl5zZuWUtVTg9kWW1o3FMOJN2wZy4RsIbNt0hRJPJ5233qg0Ax+MDOJDXI/Ie
8Zn8WaIhStKqufz6WKjB/nHf5qwMC3VcoeUBwYLiKCcuQpy8RkrvM96qBLl3cCcM
SRXmb2N4DLDrvWMnfscU3JONOqdXkRY+1fI1XDLKbYsXqrdG8kCsKoq6XMyyvMUO
ek/kxxoTYlutiG1KDXxrruERaKRG9WjsGdRugDL5YEA+XqUo6o3dw7IZn+IRFFTO
NzZ6JuoAl1q7oMRqNISMIXFRwPv6YYuX4WVJd5ruU1vrYEwP93boseVoEwLA8/+q
RH/nzfGGrCTy4V74q30uJiU6SYy1ep27RAEeQzj4Eo25hU/qPR2X31ibnF9vNAIT
pQIxr5razXMiNRqgsNVc8/QoxSQGLbO8J5BPywG28tUcVhhenyY/yTIw4v8+F3fW
fErzN+2rRwr2P90uUcRYvfEHYCtyY+G6bFR3/hn4x/aNYLCbECanYxdpzZs46D4/
xpMDaQmfjMaR8sEvCRSzX5s82nLh/4wAn05Gt/P+w4/WapIRffq+7bs/Y6Qi+E2q
Gq8XeNdsZxaApS9VFPYNwlGkFx+8qKjgC5leqOLvs8qdx/dXzgTpW08FTZ/D7vMh
zjCv1RWaaN7sPj+DdutEhlM0jUYlvo9xvQySbLILyaClE0oLaadyk+Js8KQxU13s
uaoPGCICeXLRm/7pAZ8e3lvnGf8Z8WPQvQu/1T59UhiA3mrKYuZ/jUpBTJlCS8w2
juuc0afbEfXmANrJmvHaWL4WEP9nwrMa2AuSxOS362LRJGRHDa2tIXMEbyNcz/cM
mlntZ9WtVczNu9eGk3jJ5bMvKWQz99JryUsI6VIguQGMbu9r/dHAwZj0nx3nSe40
AiZIpvpvNCSQ9lnKnOBD84YXjNOxilcsGfeLQ/oE4jpZUV0QouISrhncpo4Ap05u
4+mzHKgSx3+olYs8dmE0Ly6jY0PQ9NDvNUpNzhYQWtzoLkU4tx0OJQ6bqKrYH0/s
NIosF8RMRLwoddKALMcwppOFlK7mCWEBD0uIFhO1LiWUHaSEMJqpaXZ0Zkz/8o+6
R3T+083YdnKewgdn8ZFoizm9027Pv7gZaNvY2xeJ+wyKwP7b5A14zlJy2rJi4NT2
nUIOBWwkERkNSjTI9237BfEw7pC99kcLUaRm4k3iu9YqZaQ+SkfIVuFFbK+tlksM
NZcvq+iKkbRXtKlmlHSbFyauHbd2ho4Rh0NHaICMvHdDv+swXxexl1gNaGrHtzDv
Yrq0+Xm1/wRjRIk9e0ofbANHP2PyDOdh7jErvpdX6DKtVLY+0VXySC/ODNt77GoO
9xQoIxhsAd3eCXm9yiPeFXCH9X7DJN3Eg+GdkO7eIU8/2UmoB5OD+EhEupSVYOIW
pJWgCAFfDuQ+rWgurGMqOxef6Zx5Wgp3Dd0ItQEHzHAXAPv6kfYoiTvXtY7qQL6u
+kBshygCrSo31vB6FVrfa7jolXDCsegkYBuQgNTL8UMT5J+gHl6BtLE8V704fzdp
q29rs5iiEkhqHc+g53dRvVdMZpsZX4Q5nCffrthY3K/Q7riH6Nl1Auds+lYLqSzS
8zs2W7IJsH0njFdnbkon2JXWr94toY+uvMeuDn0IsA/NNUz8+PlBXT/m3yY4qA5A
rBwT2cfK1zWyUFVdzvpzgdO5gsyvTiME+rqTp8MOT0MgXfe83hVZstzSlC9cV1Wv
0UiV1oJu5/GRf0LlElKlhfV7Mg2SN4RZEZKYI4jkypXIXjwmDwQMs8iL27445jIN
ylpcfDdsD6RLnNBLs5OQ7nbZkYWb1lHlB798decsM0xRLF524lkY5cPt0UqhWdD7
4EyqcPo9VbXy2W7NM6B62xLLSFdafF0Azhqm9/7cvAf8cV5/NZvFLeqOMjt2MHzB
danu5knzj0dFSxE6L8obW6amXlPwEBDdvTX6oVbPrP5lzb5We4NBPRzZ9YCx2u7I
m4HbWCMI0FBMX+SVtv7J2Ll1ACVtVJFtVyABshm334cBhZr0Wpa9K9aPsb+GTVGj
eOiSIyoo6U943Qajj31IcUDhdjDlASbynkYqR6k3TPvs0P8GbNdTnrkbNuCsJPIJ
vr3c4c54qhMh4Ls8SBRuvftZAqWE3WMlWeI2YTNt/+kE0RR4rTv3c9Xu8gntApqV
5p7KZx/4WayPI1syMnySEQyjg54VaNk5oyndfumTkmAFg1cVDYMjMEH9/UdCk7Ey
dHMh2NTFXvwif8qH1DnzNdKRmsfReEQwd3B8UeQuugd5RLiJlxr8qgfrj5+shV0M
Ce+fQ9PyXrbLewWJ/SKdpMBtyrM1ROcEOZ6Ag7rRWGTYoJXSaJWleCuNp6BYlf0h
CrQrRN2F9ydpftgt/2WTvLv3VWM2tQYakm/il/cQzS2JxaVUd3NTrn2BTy5qAdTS
Mv+SLL7BbDgdySsXbdOSZ/Nl13mKTBf+58S1JBwQ2ATpD75ggDUkZpqIq1GVZDF5
efEzlUx/7ssr6HWFB/UkYNqzfLcrvEeoFiGP9zUpjkuqk7WGtOnRW7sF8ZUmenDF
xFbxtIeJtIoA5SL48XNvjCruPZnOXcnNqgfvKST4KSJfWkt3b/PFKrqB4Nicm+Sz
KNuxeilXZm/dYXja+4+U2bekATbbpJepPQZLQarlXyRb5+IqroesFN5bJ5ZPRZ4u
Lc4v6G94VTyxZxGEOGwGz7exHMc3vTRGiL1PJECaq+nHE1XToAJGvoUAcYJ1Ts39
3SNHkcIdmMxDobIL9RYjPXDeYws2CwnoW+kgg4+W+hAj7P1ZTFBEtt8HlRYwT3PA
YLTuk/TCzDq477b1bZFkyosFAflIIu67e0ZdDVUSTAqrXtiv97LS2GYeVG/ujZ/8
Y5NoAQS/7GYg14dsKpbQVV4fiKSsGPeY1WJ9KOV8wxoIFxbDvx48L5xALJo0t2lc
EYl1mEdUIaYQYeZ/DdbM8K3osQaHzWPdG9YM338cAKFdeHlOBvJa6Fsb6NaISEab
zzTgD/TzPJb9Ukp8g4RhYJolk7Pj+R8uqp/U7RtxiYsgA+jYAJSCJA1+WUY9NgsP
Ry9bnEm0oS6FLFZWq73jTe8EwjyfKAQRr8uc18E44vm0/gAD/Vo+ERA43Dgv/cDk
QPTDsM+gdZo7WhMJQX1MZQarrwipXb/29jFeB7ZV8QM3vQN47hUOMo9YyicBtDld
PXVMKl5CWrOK/mH/3U7Nvv9sAqItCo4x2vatHZWvqjTiMzV7Gcbbd25cbyzX6of3
8NI97CrZ+dIqn4wYkmRmWhUbMRw0iW5ZUfIDkR0DR5axs67RnbcTGkCZbhBfT74N
6H7f3L0Fw+mkyvYjug8GbSHO2C9lFMbTLzPr1BhvMTXXlCHytlTDfR/egOy+3wYN
0eV0anTPDSJHnBN9uH+/vCLGhhhP84IiZ5IZbDVTGxzt2dZ89ehNdrFywp3YpQ61
MlvDX1rTRkbUHW6+uwHosv+8NBuyoZ7QDj/iTGoh2faUZgAsXHE7tPXAv1fe9w86
KzwPFRqA3OrhdF6RhRl7WlJsy/+eKW1vr1xaCEb+sXV7KLT5ZGRrzOXubjnn33XC
C4vl/G0BdVc1wFYVrtSDyeZmJasWpCxMU9PyEwWZKwctWpkWgRxzzOFCJRnLYdTn
Tc3uDZXwvDi6OqB1cDePtqaIp7hAAO3mezk/vwnZ59mMkoz1i8QY45mWI5qTPUBr
x05+ndE9OM+0yiQ74HG2s2SE+Gug2BjQ5FgrdSg5cW65aXr3BmR5WlfGzLYyE3kB
AS5++eOZWZBcQH8NeMebIJ8jqn25a5Em5b6HH+LyVWzBE6wUDpWnEjQl/7dgqY2i
1PBqpKUJaUdZ752+Oie285GckZLF2SXzwuj+No6Tn2I=
`pragma protect end_protected
