// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NyUad3xJw0SO+UwpNM63mlkLKx2bvBMe5NOdoyYpQ7TOSPyA1FtbN28xedOtlCkY
NYyWR/Yn0K8vtY4LGDJ1hSHCEEdS+M9SJvbgRLMFrj7XE+9wlSmqM3pjaovBumF7
eb01t13dkqlIWEx+NMsOz/YyhlYizxg4LaLhF6v03/U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8960)
oa2I7M5IMZjAraUK4X/OOK8X6ZNkaqIsj+Z9gUpBPRuyr09Mj4apGhE4rnoFucDU
tq5AXfKn9kGfUCGldT9UXUbVyKaOQQ9ESy8FJDspKlnSzwk7PpZMH57WXR9MC7Bb
rxAyIyR45TzKbti/JOK+NSXgs3iImypZnKISVb9Rx5/3J4p9qn+hnxvn+QxuDrcS
cHcrNIDjmlLCWicm0cNUXRNS2zjnKjphvLXaWeTxdnW5IxDy5GfStsEAYrvHpfov
6V96xo4LR/yC5m0S1KFpBdWtFj+phHtTbjDoMO/x9oJh+EsD7FLvhHdqHfw7RAAI
m/pdjvNkirBIwyoRVXoLW7D9yYM7LwxZUgcTifWictgMDE7UXUEOuJRhPxW4VuEp
CyksK803j3EdvlKPOiNh2v65zNMe1O2wTIfHFczzpd6kMygzSK9LCryT3cvAH9J3
2aJjfZVUZdUFo7lbst7IrzJN5ERP0nFSvO7kN9XUk6nUTBrloJV3v2KjZ/CzQlli
t41dnG22sFtbdvh2khrO6rECXPngPu8gOd50G2+FQLjbtvLwwWaLg1dZLAnjosnU
8fe+KssABYwM/KHLshLLNvuv3NVQbGzcuyPN/hu84xKredGv6FzBTST3UQ+//mh2
zfvythynr7M/ZcsWzWtI1WbDk/L4CCm0BPaJCT4WrHTPF8aU8U+72MiMk5zrJNe7
VhMnEGgdzqLzBr8mBOOKv/e02bq5TqQgR5dZL7dHQga+W+OUIb5FSLHH9oWa8Owp
4hy0r02AOSKVh4umQA7VLlR4rt3B5S2WiKlPxloorUaPdx5V1Rv6MEqi0sI0ZAu3
cWRR2MmY4OaqoRnWIdY37sdQGuFoKzTLR+1jW40xvPB7zsFYHhTx9WrqsXejhPt0
acTCzou4TH2pSsda7WwLJXTUU8U3DcKBRQJocvMLUJXBEC1JBEsgth4l4UNfY18b
Q8CDPT7vlehOT9QEoF+GR7HsY1zB8xSnRd37bstQVbAXxoIj0LWe/m0W0Ycv/R9N
Hd4CvcOArxDUNqjUiGRp+geSlRetZmqsNslGZJHFUKtY9VqfpAQg5tP2WVbXy6tf
rkiIJc7SHIaAr02pdk8fPi+CIlT2hfLxqg6+2eHIakri7dSbFpe6Y30G/EVMgjAl
x4SEtHXs0ozP2ZZnKy37ektyktUx7vOTF24XFIQnFGAngFVjoJi5ZXs+MtuMSQws
EFkyiAaLbV7E5oLUWGA8Ze3jL1hesV0vPxmUQ10mjxjCORDIC4YMyzw7Og39jhSe
W1lycOoltB+it/Ewhmfmo+Rl2uYgaxcTH160CZqw0WtFNLbq2GD7/YHE0kSWUkv8
jKJKnl/rzMvnZBtB/Ca79ELNnhclNNDM+aDHNzJTknSiuTJpSab2GAlLA/v7fhAg
JB5SIl5Eb5muXU/DlEMJRqWnoSq/UWZAMv+eC2q/0f+8Izx+/J48o8rx4V8DCVbD
oNofoiEvUV5LYy09tGEZppnJ/JgYG/hFHd1mE1Jee8DphjLJP1lCSTdxgew7gPoz
oXYpqBcsBdNCI4zmI6s7VF0NK4I2TY613383gk8hAm2EzYJCRn5wr0Cditoy3YpG
/pjCpehj6tTsRYw969zU3fJixAL7YXWJWZLMn4lYbRCS/9R6nKKzAXiDnDR2N9ul
Re7wAA4lw7RuW6vqHCGiQhGRXfBo/iB9429bQr+86jqD3dSYQxXaZI7T4gbvRj+L
uUUWyXf/oD0YdnmHNBf2ZAliBxzYlSgrYPvJ9Zc0b09h7rj14jpgVnGMRqo0EWua
W+8frjLBI9JEvS1tOOuGyqgJti+paU6Q2NPpmwkyVSNqNZi5Yz6emqJQXFlJxpri
iNsjGo2QLFNhXcpsUAKQ1EZHfnJriJJAG72XFnVaGZ+B/wCq4AYMQKPS2JKs5kRa
pkgNTCEG+y7Z2z192eZAKNJtSjcL+sqitQsyiRz5cjfmnU8ViXD5gzBTRT4Co1aE
aaCh1PUJDBQxW5Nbemq1ic2KCj0AyBLja5rUZqlHSBcDt0b/NT6EIt188NgxJg4v
MKRh8URcFwkVY5YkDsMwBB2S8t/7+/FcFDm9ZkxMvULFLJaFj4nO9oKrtwVT4WF7
B/SUwrLaTdeQWQM7Hm5qp3mh3RbFy7eHMw0A03PVj7O0sDrJMnq7lCWlid197TWQ
BptRqOqKCW6hl2VfgogFrpy8IkhWTd9D6MQWOo7CBXcuznYdT+MlKVEoHR7b5sUQ
6Hw/6nCj8G4JfpKp51A1az9QukVqi/nWg8KNYOmC4fl/mEd0Pz/CmYYAHo0Vyaz2
tam8d27HcHfvVVOC2BwoPLYJW4U3bV0cpNf1efgW64/FWWMq3Iv3WsFCgbghaMCY
w9hpYAanVnwYyrhQpy6zpsnt/PO0I7D9MpG6gOeYsn9/zJybfn080sOg/KwRzyFC
AqZya4e0lAUol8T32ka41AFdi/6ErgpW52NHOW6ot/TSShxrzEjYfXlttKeVod0h
IxmUa+NBOSlLrpAG2y4mqY+jmGEoDQ/EV3Ordle3TVkavQP18dSQ2Wz5rwwhBU5O
YDTYTxzhL5QDftL+ak5GsXymIYVvcufCMygp4FuGW/hvIQp+Ci2AaCruP5hPDYob
YbFeKyaYy6PI4ZZssQBelczcDaBZb3GtERmjz5O+A7jyGcgRTdtaEEedMDmrNCJI
5E5b+H3/eCzP8i2GPwU1GvnneiM7hYv967fP+gPAc5vfN9vGOJ+esPZkw+Uw+chc
bfGYee86eb06VsJWW7DpdVDgt7gj8bfrASWS953h4S0EAqkqrrF9x+U1iWfaK9fb
hN5B7SPhQoLLh76ESVsfhQXXeaK6nnW7piiQlwsDO3BcHK6iB2zf3S+0fAhtGyBt
gkwNCl5WlKjeLtqMe102T5kWUSZvGMfGNvV9XkoiAmiAmApufbF/iAfhNegMJQsn
AzrocJ3G7Y7Eymj3lACwDqnoh99JebFe7/lhcBSHze0vxrH87brK0+BQ+TvjPD7v
s+VyyroYsZSQ721gzA2CYPnV7r/gZGLSMrZYXvinH/8wtBR45P5hltQfaQLyfjqM
jkx6SKRxVTkTH5vdOsaTGVQz7sDsw9bNmh5I8gcPELCQPUI2OBXA/ngsuRaLXPlV
EV8CcU9QVLqwOaXACVKamZwMPLoJTeaQc8iV39AG3LY6ex2TGh2+tqdCvk5QyDMb
m9ACgvfufCyfFwK5VgDfJZK3PqIMA9624fnt3t3KdLuuleacrQX15Bu1tkegaQFV
st9rFCRKJMJeJPeVTT1mz7g+xvLWPD4DxyNcxGmgbTbRw3yPTo4c4zw3y7iIEJ0x
OwLmvdXhEHQxTBHEp5SAO5LAU18HH49WRmdK/RPWjdgUKi4nlOCGAkDi60RoV+0S
kEZzt46I4vCrkPHQjYbDsQl7ZhRfGPw6W+FC/i29vQDjx+8WJe6mLkFhR7W3Jzxb
iQ5Xcmlf1zcnZ8p8eoASx8+q2GqrD3yE/PZB8aQGVN7rTsV5voIwovgzK2qmLrt5
0ypr+9sj4jSFPg2mhdbnP3uV49G5KbvlZpv8/1tjkbOStu2Hxix99f2LAfzYHG4N
l+WbU+0Lqtpwkt3xC6I5kNhsvlpjtVVP5QSbgwJSzA2Qy6MKuZOdaL7p4TxCSQUZ
HMtQngeJFrNbW9svUnuojQFdZlQp6x7cBiN8Pf333TAjE+DGNOIM5pN7lmmaYBrn
LKn9WoQQBEI+nAaWqahyhCtbJ+hObOMOfVHErc4TlbxG/ZV3pWjZMtgKbpDdDNmI
Q0Vd1C4+SFf8KzpDzeyUVwpQKkWfxkcrQIoKJslMGOYLtUOKJyojis0zpu4V0JOO
Yf91gUg6c1DV23Yywv+NI8BDVOvSp19SUWU4WZStifYKDZWPz1uQKrgEuq24p2gg
2fVGiWYN7zEpRZ31+ZtPqS8ZV8wgauJ2z2/z12bpZqO0KNmsZrQYUXGNGgHuYtIj
i8tLZOllDXEECbgz+WIbBcppyFqAG4g3OZNCbSL7TLkGORYxrs3dliaE/BsNuQX5
KXF4+CPvacMnH/h7KYwxVsnohsR5CHmE4bz7h24+0XEi90xVAEi5wpo0JGW8yjd2
wzXCxD77r5xWQIXVd3LxRWd3sK5rN8bE1ghiRk8ECmNHA08+Fdb6MkmMwvxKwDSq
GsEgsg3oxqaeNOStJsEpJs+w/g73vkTlIciJCjtA2JCLyTIgrfcwc61ItToKjwrj
nLlqrXbswCB5nYrllyqRI29BKVZdSbqvvNkET0I5J6Eo4n2KoPVqnMVdA//6d16a
BU3ZJoC+E8jR+cK0A286tUP5aqB5SxfaPwSy9gBcIrbnybi3XAT1ZD6pYONUOfrb
N9S6TeZfVr442im2gNtRy3xdDkTjXFPsEzM0N7/uDgPqp9Pz7lBDSRiq1tVUzdVR
pfYMWQgz/5FdLuPnymWCT6rAurwz5q1uSnqwuD/OI/rGTLzKsFmxoB0j9RL7Dn13
CzOhULisCg96h2laxLQrQpH3Lm6pc0mra7XS9JLgLZKX5xYTqyIKZswvzOVqlwHJ
9GvH1XGTwaJDkJs8M9cOqO6bNSt4Lp5RWz4sySwuAT4tHzWFb59/On66EfsJaBUj
RgYFxZQb73Xp9WQekq0vUkETYWEMmu7sKornR2ID0v8P3yF2TM0UY89sJi4UsXVo
yR01lXHU8ePlXQKzlQFWZ301p9aSGkadE0tZ5nRMBIWdCqjDBN3gggp+lMWV8WSg
03bhzSRDdBzAqTeT5Esqc3o14vrcKHVz2OXqQbyTLXKx7t+tIFjU7SpLYiAiV6ad
tQxDlNwP+H+/ZKfCOUlPqPxuRvJ0K5LdHHRzSca7K7MS2OADtXGY58GX4Wrfq4eQ
YMTu3vb9qWQlLIpg9DzfP8ySGwR7OLwFI4F6foI8oJpcDQh+BYoh8GoVG9Pw3si+
+OXD1C8KCApsqg/qzpyb7USbNL/w+uq3kTz5CRWqocM3is/ujJt9jvDgDQHX1i7H
Shc1jWKR3Hb/DDFfnkLZttYG0XNWI+C9uJOrH3HqAelUDtmuaVJGjWaXA7ipn45w
F9cDGR5dHfLJDpyXhaOIOPSyrEORMImuD3MoiYPIdfIeNK42CInifhi0N10Yyd27
T/4rt5H8lj+wK7Ll2Ypc2HgjrdxLPYf2qT/sipblsv3yuJ7pWzh2+mPQpXS3yYsR
5/zKkrTYlpQ6OB7SUcNTL4nWps7QHjZp4nuGFKF38JvUr5IZCNpchtNWE+fa4WFF
2xfOzBe2D2xQMGpj8De8jZ1cSLxK+MA15yI9WwDRR7MzGcULJt82M6mGBIxjKMah
J3rcUOPe4O1X4cQ3ogml6ayyw2/oQfq7p3wQkaAewhyPJSFFINhUnfRd9tb3/vxj
Lp0bHEiaBzGSCwrZQizFNdYhvDD/SCRxbjNUqNBDmW+tZeTl7vZWgWU6MrtVNUUV
2XIIwFOU9b3/gPkcYW55Xn/+YhQOL4SEfgcZoSXDK5cJFjDDdgSP3V0+KzGA1I7h
clAHuJhrN0/evou9aLOVlehghoAZiCJf8nfOHhn2AFn6728krgjcfOXFIN9haack
nb8J1QfKJHnIlglmEjyfX6S80FQ51n0TFYgram1Q0T4m+dWIxPK4U87V1ddhfoFh
YZAXVWLzaIlCAX5XSNwiGOe1pICBv810vxugN1Fsb502cbfGMBOHKwQgGlP/+LDW
fuiIvzx+XKtGv6oLbTEJ9H2gBI8WD0VhQFXD29Rdn9EpHke5nby+kjU1RW6M4eBa
FjIWAO9SDnlij6pahzR8s4xLu+Z70C2aMuMjMGqyrgYcIFjrb3JYt0Z+DpoIsv6s
aolJP54EMJMEPY6kNudlLIpYqOmx6bX4sLQNQR3UC+kiXYMLr6F5QXbY3vpPgr1w
ELZo/f3cFfVdBULOLDveTBjmmhWkFruiGV3DN8zx+AXFa9juXkWWWl5qjVXIT0Mr
yP2tBdH33kf9OweNWxs0Xr0k01dg8Nvl6S48lWJSZPXgiWexV4fZNkMyslqRJqSw
tXNgRNaptXJmDhSKt2VopOPFKvLRN5FEH+6VTCYGMiMZKiic6n6aGuguvHmOdFDs
PULcSDb2ZONLr0P6KbmmYVxXddSxgo8T2Gub5YgkvL0Eij7Gr8eLHWv6oAN/bbA1
UtIJelhyXlKvJF0ICSf9KbrrTaaqXqzHb+bnEaF8BOy7I7oI4bW6OuHZGRqNOf8G
ITVzmFwpRgTtB0Ra/H9T3PAvWj87g2/a+Zdjot/k0Xt/BeVjbEx0XsUo1VzQfoRD
8u5GApWXJuZXU/xvDevCdXsu1YxANxRj4+ti85ojvND+gOAQ3hyvE+Ad7r7fmwkZ
RcUInMTjnvODCUXkujoU1bHL1/FiTaBCSz6MTA3bdsWdq4stCWMDkNpkMb655652
DuxzdRIMhAKrkgThPk6wkBV0djTpZndHEMZUCPMQXq3iTYhHyKG5XexSFGtlOAIt
EsarPZpFgjuCwnbKQX2cO/q3iK41o80YXh+mwBkNSlfrGmFnWy8ejNBRnftoutk7
RUAZ5w+L0vMaEkKG37VhtB131llU2P6caX1wWQ5YLdD6ZLBs0ajRvyrrm1WwUyth
qbo0QeQY6CoPar5XapDhIfloYLW7u+2pI7YMqPfoB8s/LFUtnMlS1kJoR7ugAQW3
aC/k1u6LfteWZolnej20fXA0GL4oW65C0CVyQe/L68TzMPfNaIdr8mW3C15dywrb
A7Qo4ylzvDyhQpPTy/QZviUKb/v48nb1r7+OGb15+AEerL0XtPub7utKOQ7NpdYi
sBfU53GiR86QpQZx3Qw7fK8fNqK3x70OpZ5xgj2cWGefzEK2vLYODBM8hvWMxCYU
PZ8Nlq4KqETQ1myDGHyGIewEtOSUTcExjgRte09CJn+wAevtNAeKkXqEHWDRr0s0
yjUBnjONhkVbyirfizYFJmTsL57/jC8BPOD9aSKkb999ungX5+csLVMrpf6P8G98
RgIUBnEKieVht99nbJWbOuNkAxMKmETGDCFBeNuyGqUtRsTF7bLTk5p+4YckblKT
gstW9wnJasCdM+NlDejlUXm1cVYtPe8LtrBLL5pHzXlu9a0j7wJwXW2qZGVh0Gra
XGd8bMzUwt0yUDy8Wr5U829ks5nHMs48laFzFFHHCEAcVQ3vx5pyLYHmVgq/3Mqw
y9aGtBYTSTLHrmxn+pr3MeJLyf45K8oYG216OSGHbij7LUcYI6dOfDbu8yRc4uPC
1NOPgTI6jN4MNPfMbsJGJyu5JotQbVnD8v0+mnnzBIMIQeDKpbM7iHidZk9AZLBu
uKgUEkzXQMpdep8GFbRGF/GUtxsb9e5f7deWGQF+iD8drIOxvyvoYFsIogfwiHzJ
6Mdh8Idd5B2YO3hWXxZmRnlORQYLAzei26oh9Bh3ntQpE4rZ3fR3GuwcnA/FiwRc
K15TUooVRUTLs2fXeazS0FrnhKK9hHL6dFFE7ein6tCyu0AZHO2ddCcjmDjIPa7h
Bp7dem6OzAu0rZpN9lEx36MAW/lQVCCSzEmQ2jypmA68cbSRGsipJn+KeNSeIIYt
1a0dUwiWKgSib/KZ73BoLsBh/5dsHKBBozsLl94Fmwe8XmCpyoyNpIts9JmMwfvE
oSSnDAm8AMGBVAZLQX0UGm6lkcP2omU1HI8YoLxIFBOk7oDFl04qjRG5OjmMSQQp
hsFVe3bUR/k81V14ekZb4C+VqsN1eSN7RCSB5bmMZe18rCDvR0kMu7fnoOZtJMa2
c+9Yqmu+RQSVpMv8sfBZ/+8Ry7lrqS+i4lsCmj31ivcunSn+IFoYNv8B0UcEzAEc
Y3GnLHZ86E8MrOui2Hx+k+pDZXni3zfu99TCM52/pVy+HjUbSYpgRNOm7Nxi6SWq
zNqaEtUi00e58S70vEJbpdJUeeK5/IoIl5NIzVX0XWCXGLcSFFF6zUsitbjl1r7M
pBfWA0hrT3WnWf1MpY/soUMMBp6/e+9ST9Fr3kXn15tM56qsBAOeg6zVaZ2Q79IT
5NItEHRYwXMsUl2WLCuPRVbG/oHEekMWF94Qsl9+PBfPG6rqctdpkT6tQ/5eSg2R
EZK4XMzY+hwmuMTa5OuJb691F/zzU1sUNEa8WMzu3aFzq+bMeDOtXSdFIg6xXb7/
x1Y5MEvD9fcWBblK+dpunWDPtBdr7Q/0yK4AL/hKCURGqlsYdD8l/jD00RJi0XE4
mNFUtwIo+Wl+oTfAEUl2QWEzRUDMsJCgrhNZ/naQFDSsrMr06bVuQvk6BOmTOIkm
WTCixnOStQKCAop9Au1lcclTma9Vq3/W5w6CasTuVnUDupN7hOQ1TQr5L9ltJ160
di0mdUs6YVh9dQ4r9O8wbqBZAROnFYbkcKjFKUPQyTrIBOmIX97eFUId8Pbda7OO
VguHJd34PAjGYngryTH2F7p+fFLyUsF2BkyaAVLW7vytrRRxxe+2Nf2J+suVtz20
k19qKBa3E3EQrC4vzLybo4b1beHBFgU27LpBpE7QxA4Fg8MzCerFPNIecM6OxH1o
aFUAJe4Zxh4XEBF8Ks9SSQISfrL53kTYJ2dYdY/iNc9dZZo3esa+MWmVfvjyq2nG
6lTNG++f6aT5pjows2TYufxZ+lBqJ9vtaSzy2P4R27I0RfvIAkhmpN+wVh8HeBOp
TvTo3Y2G98tTw8dcoESQDtL3y6biTi2Yquc68lSGiCgKnUf+SM+G+IEE7hLOUXAb
6JZuucfaFThwvWanqOiyyrZw0xJntoQagIapPuO1jBTTdsils6MHmW6gZKjWqaK/
pfygZ1w9qO+hN94T6jspZYwkUIb2LaIJ1TfbmL/AYEgq7TpBX3we2YivMp1d+DC2
ClCJupEL1MyhtcmvB2XPKkvIB0mF2ZTg8n7HsoB4D/EkzRacmH0on55/hNDHIyKr
1eCTWMaX4cRELjbKgVOtxkeS5L3WqO3heODdtx8f0nHOgjQ5S2/gQKE2TFGL54AJ
4vKRdd6ArL+rU4ex6wMnC+BaKn6fzN2X6pABKRdC+L9uIGzjdTZiMPbwF4eSjfrL
O8WIb5Qw/RjjUQRfhJjnyXcafKNX36KuzS9Pbs0xhuD/ML7s73zF6ILk47SpAwOR
JT16gA2unjCJeT1FzjqqfC3oVfRMv3hCSLnP+BmRE25Mybt/nN3A4CvH9K1H7bnO
dAhrs+HxZMV/eG1zf9QkNz8gkdRCVpACMaDU5km3A+NOBHsK3+AaFtQqwIToCA/Y
Ga0o2J2naBro0cVbruW3B+iUV5WwvG13c+qjwz/brnftTcjz3ylx8aPn3XUHcY03
bu6GWE2gph1UeLZVdsORKa5vx+1e1e9Ot+M1zwn/K9MstZtjjRWIIzaE0Mv04eEd
fXbHvaYRkxd+48vsKwATBTVpjrNDhoj25eVPV5t67mVFQD756FOtPsqYz/pgsq9n
g4g4zzZcGGI5W4VY93gzMYr+7825xL6pDYuibFdPYTVyvU1DnW0ke2XHiy70/Hz8
uCpPdTBWqHB1+vHh3W5hiX6HX++HbuJhR22EhO/9+eKf7ORLPq3FTkNTral0DtCO
vIWp6AJBCGk8WBOZsGOwU+X84ARzxJqZ2SZncjXE9uB076fZdAmGHTM0Yvp+wxqr
cpM7xme/qOWJUwl0Svwr9hf+BiDvPnIH0s10TH/pa4ZTleYGqPYJ/oeG7u3ycw/e
oIp2Jfsqb4g57MrwBHAqK+eS/ZOy1/eNR6bzmcJMqyEFYUbPYmRk1tV9pmJngOs+
ZzzA13pFDlReLVcj48SkAJFJiUkbdGI1u+3cVCZQPrtCpuwWMhQEbBMmVS1lIb8s
8OsKR0KVyIAO8gIp13FWa+oEdXEdxr8F0+AhjpGEG37yAy91aBXqrWVvIIdphEWz
3E5IOq+0fraB/2W2Th719wf0ftpzpRH6Wk9ptWhTOrfe3aOCpB1UNfTut2WvvsQJ
wfX62Rc/pEa1INpO9kPuDS1hbeKwNnZgQ5aCATnDwgY3Kohp+OLmZIZrmxqfKumC
x1wFQVMuHz41IxwlMLXKoUPwgxBhJtBcJxl2WxsoQo51fVHgFZ08ObeZS7Aj0GrE
Gl40+ZIHfQgQ+9wOq5/lAzcCAmcJaZsOxP2NElmTzZ2coeVyQPSmA8EUXsw/x+Iy
lU4AtWAO2CcxPrRy0EERs3jl/Qnxx5MuTSS9R+lD6GvavJHtczPD8TuisJTwiHBs
p86iKjBkOFj72eMUqkDStx07BPU49BR0QsvyclGuaKGGoJ1SNfDZ8EedY3voOond
fSRJXNTKJ5iAbYtyFAAS2ygoqEz8hvASuqnKhROEs6NurXlsyuaqogPbq9gMR19e
P51+1T0yh+vvUjjPYzI5CG2N4tkkocB4rHl0T7R8QKY1ltUG8xMcJzFBMV4LS9pJ
60AZ4RdXLdsPC3vnWPWnxQu9bB+EcRtVEAQqx0YZma6v9tq2HffIPL/EnXKJETY2
stWOUF8z7QmEbD3oXZ68M+MUT3RZgg1/Yf9cxAzYOJ/wnMOBJtQKnwwakHExM8+g
ib7Ib8fnCoTw3phnpfLG+YhG1e5Z7btVm0RLLaYRzm9wBG+Hz1nvodd2c2knDMw+
Y/hHPOCHOmijriMytGgEX6YWbMluHSjClD5YXspJr1Hi4dNAk0GoOKewQqts0vYW
TCsxOWnCrfIezxlOP5QL9bSWJz63A6fPa1cb/hmxQ+RGlXFj7IjwUlC4wG0tWprs
0tHMV0XY/YtXoj/GtA5+223ER7geZh9rAd2gtMCWTUKYGgOGbmoeu2cL1zg82g+C
leiGdERCiE6R9QJLazQtefi3oWmZOfjXbu4YHnC19v8tHoavXSr0HsOhdoW2mNVk
wQOvkjiLbpOHvvFz0laWGf8aSTL+5urS2Kzf1RwiAddCH5qldX3MpB8W8HnhAaDe
quTYRHs3da5Rcw157fXMxBfMqsRCcmpIpOR3bm54oXFeuMdvu/qiFEXDr1jbPA2e
r+1ZKeH/gnaMVyiQjmhxwvxYtYKBiM27P0082w+S0u5RcDRQlihuJc8JlgwCIo9m
y0VsTa/HrK+HFfFgwn2coiN9J09S1Mr+dm7ZSLa+Eqb6oZZrJJOjEFq7YklUhELu
sEfbDEBbLOcedHvNGcAi8o0bqKGuLeFjP+jjs70i+qMpSUZp+K5yTKc94ZJ2QTjc
E3tuhd6/jt1ycWV4s9xlJlHa3eFa9J8UAjsKDb5VyUiURt2/uXpfrvs2eVKKhjtz
/qIkvDqXYI/6YEsbjSZWBDu0390QpPNpmzw8mxry5aikrZZ7QsV4b9YzlAMj/TAt
QBxxIz6PiEMh7FuWnGHPSA+1zZPEo2u9C9wNTVmV8dMC3sCdu4QTg8+xtSPd0umR
Qu0tcdDynyjGp33D1tLKp/ZTEtD9NhjLJRfgt2+taYynxSmSxh6rJQvlO/9BZLv3
T5m49xDHJhbKShLyrriJpMr9aYzyKr5Ln/05GDuqZUASRWazJCNBRNjrr5VFuXW3
qMRzBqWV3pl7+3p6Ut+ssrWeU5aZcOjCuIaL1cRTflsuXvmVU4u3icipwXZV2SQA
efFBwdpzmFIkRxmwZKkBN9GbR92LMIvUeFDuvFamxPVwi/wOm6lNx5NX3p8ZJh84
uqabuvtpqZqujNvjKMfXzotxYnWZPeTtCJEzrKIHuFf0jaPSLevde40PtUCUZ9bf
XTbZ64XQsJqJJWYP0nEfCEOJB56PY8vCKvU6cJz2SMncfCEa17YpdDnRfbyvnGKA
cJ9uDcVKlQg7CgHW38Tel3DM31JobQ51jQ9ulTTEGUVN4eOqlP/FXQ93FVvF8uWO
7JH/e/n5nDNZMVLS2H1IAs9ZTzG5itkFgSsY+pBBlK+FCSWRYxAWigP2EURh0bBP
Gfd9pV6xB00EqchNpx4HGoQS2OJ+w/dCrnZ+CGpKe+ACZL8vXEO3L2JEQ5N7p2Nh
1n8dfQsWVAXgDllpaCQzr7LtViK06Byb/AHxXlthzfw=
`pragma protect end_protected
