// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:34 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NtFMHsqtm/wa/ZM0uNsgzgVoEy+/mDdTXjmuxmJx/xbOw/0eNS4/Pe7zAaZLK+ml
R7FLnOXpv1BZxwbZOPcWrq6+t5GLCCGH3FdqOMr/twp8KLLDiYf6KpGRkiG8W/NT
Z0/ylB2DQG3NhMmSbXxaXfFS2O1IF//BPdB8eK7CYC8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5216)
qEbTd1z6TO7tkhtvgTzGhb5/JlIAuoZNE3JhvPTwEyp5HOt/uxkMoKNsbdm/fz3b
tl483Cd9Tp3Ywzn7jFcMAYwO5BZ4e3qLC9jjX+pxU7JM76IUo7L9hZgEGHHNkDry
yBMUe2rjiNCuywz8hM5zpx5mjO+0LLz1f/yTCfGjiw530eFiHCWDGycpxg9kv85J
ruQpNPEK6B9QF3sMJe/gquo2uawlA4myFLVKVZ55tqQXeJV16L4oTuDlxoSSORia
76tCkz6UexoUCpr531jqMMjkwfOZ7UyUTeyTv5wELGv7jgFeeFTjC3Y2XJ8nZD69
kmLSTm9XdgiBgu6pXoaO3UUHYqSfPVEARY0+U6aWbwY9KNRsYDolSjGTiTW7yAIN
1AR7yGGRW12FMXP/qIqTOhq2XgDA6ELO1kNPdI71cqdEqZrpV+SikwsNnFijupEW
ua2XW9G300tTBW77MPjWxSN9K9S0SvReciBpyEMkeS4wUiR+dCJZAev7ABqGAhdG
3uAZ1rqGWNTlTDjdMgfcFpsBDInHjk06qRo9RxUqVZIAcPhecmfbBDpsx/jqcvki
zi8VkCZWoC9sjsRNt0Sqq7ad+njxPZ/DX4p7AdRbNdpbiTxHP9C8p2uluBqj73Ob
QWijv1B5Uu3XA3clyWxg42eWM08j8KHcgQ9spkpljcjeowP8maA4TvlIJSjO9USK
ubGafyqn9ktf6UabMgLnPnDO/wpnHrxxz1FB0spOn/NYF74plMzxAMkeAHcD95WQ
6Uv6kqBBp+ncrVLWZ4r2/c2PoaJRrDpgfxSLpmFJdbduhuhdBcPCh+d+MC2nV1N8
MzVDvHAUSWADII3EB7PrtOPOSy9rXLjEj3fV1K9hzW93hMEWfdSXjC4H4oqn4ilY
fwtLQpIiRnJuT9uxJD6LjRjboLYLVvCQ7zB7uGLFXq9lcGNgu12zdpeNbMkHl5o1
ZTVChCpV0ZtXhPYu8QoNsJSmjLoNQZMmXoMj/6DrSPY/4jX5KL90Ffsm/2A8GkYV
IGuUmGyUgTARSFxAm95HFzTYQ0GUbyWkred3SFzr4G8X1PDC4fWARsfZd3QC/mmB
l2lQ42ZeWBqR/C32iAFXUKjKiYATh7mmH+F6mS2QC34U5gv/vp0Cx19gtiuEseUl
IcEqKbks9yjuHVLKRlk09jmMx5yL6ULLG3QPpQ1i8t2CQSFtrE5NuGtmh394m+mw
Vc0GwynkQTwCp03aW/km8HShQ+WhtiyaPW++7Ya+0m2diS8OAwhkoDV+gPDFHbhq
kCTASsDHIMj3GR024Ob6hVDJWPgDTq3f6YX610Ryooo3V7FgbUBUGTSO4MCFrZIF
KN7jSMgoK33mCBIbImY4ozOWcKFDfFprBmvbBIuL5VxQxs6ZI/GOH1lS/KwEzjA1
Iftegm7ekBNcC7xyyQu66DLRJV9Pz+MZZES7ReOhstpKfu1OMOcWGq36P4oc835h
Fjfa726geoiZekWbkpJ/9Zad5FpKan/n6pT7r20tnlYYWiiDYYNraSE4hE3OddlN
vZR15dzLvd+NjYRuLmijIPRNskMPcNp+cYLqEEeg2L10j9G1fOI8BMbrMv8KSUI2
vAX0gHxshLnmgPiYwJoBupPn2w6MI+SBOTafzsLDUHqxZo1gHNme6g8X28+1VEwg
xfybJDThxqUS7Lfi4yFCwu40LxO387dWjgpYdjN+4cHTcva7woVoundLGlnPhGMf
msCFo26D6r4DWT8H7pkj6qHFLhTdJb1gFBi7D50R6AhIEbv0eJotSh6Vt1VKbSEO
Fpe2TbhRZIq9OzlkwlxUfaD3HfZj5SDtzGx8FBbcFweHbTPVUkPek55lykZEMvI1
fM5K/LkBN9W12Ruv/22Z1dtrr4aLGmJfe2HI+zIGet1+qgM3JO2Z5XMi+0We1Ty2
XJZqJlXtL4gOXP99CSRQx8aXmefrfvBVTeZPTzsKB2K4aGqWWZK0yj17C+bfuJzH
2HraUhg9d/mXm/MnVOeBrvkOCLJ3oYLPbvwPkI9GBxrc1ynCCwNUm1s5IetnVorY
48VKTef3u59FCbWDt0FG37Pul8XrMaMhfB9ANfZR/Z9WNyXG0jljt4jDTSjDiZMG
fe6c+neo59EfKBgQ2PmNr43jvZPzVCTNXb0tna4CJ87O3Nr7OKAvEwbLhVDJ2iNH
nJwaath/dYx0ditzCbmeWvEROFA0Km0PuB+qBFDLEkJ8eDjeadZ9D92nv5bUNQte
icS0U2eaK0kL1f80rm1u3FmihhjqaRfkOVbegiAUbBKtcC7JxLqn0Z8mi2TIV3ug
OL9IKavegMmbeX5GYHAKSlveyn2Hp98Rt3kQlxDo+vP9iY4SqcEm0FA065FHq0yy
Mg76SSg7bDRm+fKMxou8UX1KZki2fN2IvLoSHw2s/NgNG4Jgp2Jhy8Evg9DnDYWn
Y/fgEVQuPoeWAMNAdwVvDop9x+XfCGi4R2y6A0qSxes9j3Sw80GLxuuawgiFGokV
uTjUki31iT37wQI8xWIgcsJBWJd4cNh066ZOFHiuToyH0t6m4V/HMcO3DvNdXcTR
vnst7e705HIlcH4Fv0PIv07O/8weKECW2GYr/FmO9LMkN/fZjn0u6A07XJN1wEo+
MpMK3ioM2LgIhYlToq4XujcSSgNY3oBcOq5fihpWZQ6UGl8j/VB3Eucj1u51vG+w
rmuXuvSyCFyOS1th/4rLaV5orvozPF9j/U4DMiBR292u5WjQw+x1Kv+uBpdsDZ+p
66GUFW3dWJhzVPI+f8n58ma2YGebLmZHfrQ7Z7mQYCTYYrcQ14t55QB0fqhlYg5Y
mDYfjMrPKHjV4exTS76jbENtaBxggZob6Hwfad6A6kdbhVlf0oG1BhPa3Fu+y0o0
qxg0E46cRxVPRWKZx5PtEY73oCzfPMXl0HwafQy6C+x3ktCDWUvfeBKq8f01Wfq6
VLZHY81jKp8e1CDbG6ud4lgSDCY04DsTLCvM7dGPMdjEH3d6tkBfJHtsyYdsB/R6
41kiCoQ+DRZGoFbWUaE++j621Qyaw2/eN9ndOmh5zTaSL3KeenPETpK9VDM8o5fj
awWEOT39dEGuok2ry6ktC7YJazp3yRv72hjLlPeLbfYLirFhL1CNwLH8azT/Zbwf
/MuR3JE4YMGg1Q6gk63KpqPs8qgw+radGCnp+tI5Q1DFtTo8cesisBp1qgrmPbTL
BkT/LU85SGLaYNkeVR/pI0uEPUcsxM3XkjY728YsnfkQvGne67sN86eJperZBL9E
XrLoFUoLASfiwj9mJtYpZDbbHOS2u1khfcdz0VFi/Cj9eWQITtctgKC07eUA89iX
Cuq2X/iHIEiyHOh+Ur8n9/zm4ucsAipoFn4bjt7qNXjSn59aLHYwbDE3Qe2fcZNx
TeOoDH8dsE06gsVjWhnhyWgtX7GLrOGp1kWE6ndxQVkvKNay3N2mdQ55wEoso7xz
hleumQ/BZETovQgyicUcUiJ6e02iLppsOw5hXpbI4wQKlRAg0N+tPKivEtUamMWN
YN5KPFfGX5Djwdmrmq6tJURgMXBuzcpQNzAjhW5IzyPHy/gfxcP/WeL4OIQZFnV+
7moznOgT1EBzgn0tb/tT35mycyX0wyEdp74LtuxPkym6cizKrXwgQBIeoT+FFQzA
h1vOmSOLsziD94dxPOnKh3FrYERuIxdc6pYy/92M9TdO9+w5u8jGjA240V1GOOtr
MtwqB9ZZwE6pt5bKr0N7LH7I+tqNBkWqIPwjOI1EeeXzL8j8f0tGq/Y9fuWN+Et5
QcPkuofX7i2f4oNQZSL8t//UBBto691F/2ILnXqs3AMAK0cn5fDEOfLxfq+1jeC+
ujev+8+BoXh2tAUmdom7XsRB4BW1ukTfF8BDxVSpeSu1ECHfzzCpkp+Ozrwoknr0
/h7EYFf4FVJJeLKHTn/SQB7Ip7AmQ1S3JgJdWssc3tTm89NMUzHdzDeKKdR6q6+H
X72BuP41uPS5KlqVT/WeRVbZ/aHQ/zRJIZoDI1OWR1wixmYwd3QfWkekd46yMC5Y
NoIBC3W3bbqN525D3IH33ivS80NY7yh3pSbb6crjvCDg9UGWIunm1OyQ0tdpsh9f
+PK9GGFtkhLd7VpIzkmgM0JAXejVt9+4BZLC/ZIzZXZmfgOFMw8me1ucvrriflWW
eCgqtBNpZy5CLVC8Gbc+lyc7I+YSlkt4XWqjfrRPlRnzdX79p4e60nNOjSqHi2wd
rSa3mYi/cEXGc9WPo3Ruam5pzzOsaA5pFmFK6Y0AvOkCj/+VdOhPFSxnQqJwXgtV
5BnOOUlqu0jEZQ9IHSHdv2lzgkLBIQkP0H/+FlLiTuyb7YkdiiHDe6CboadKbamD
ORKSXFCWHpgBh9dxIse6etTOolO5DOP8ojvl6Eq3iMzOntlY7Dcr0MN9nj24Vj9O
JrxRscvu59GylGmWWTPMwCxr8cMyCGIFQE0gc55PD86R1hlQHlLt1/tMmJZ3qfUQ
FPJUEVpJcruwh+2v83ouoSlW2wu0L2YwVoNNJ1mT8t9Atsy0fuhZXIYlZEQcQH8w
FJAJOiQaYr1Xh0BpiTZqytC18fM+pHEckuBEB+zx1q9JfWUXVdVPIXkgHoCfgeEk
zZ9TWMjwPZxibTNzhGzs0CnmubEdeB4JTagqR+GpmhNezlNuGhAZXP3l7CIFqDX7
AxNYaNeMWK5JKWjT3JtG0Roeb5vD0BABtwaj2LwyF7HOXYkgvfP/GEBifHwTqM5d
H2J/vzDVmtOLubSkZdqWgUaCXoeO0lnjm2ptVm/lY4DB1j/bw0yThtqCaKMkVsjh
3y5x0ZhyUK8peAQFxgHDklFAcbsO9fRP1HcnWM6fTZp+Ce5Wx7sI9bcdguZKA+MR
omDswqAjEyk+wJHgvS8BxAXyo9iphWRGubzER7Ujv4SEyoMf2nz4Wsmg7AdKQHgK
AzepuJjx4Q4BK8+4kXawNy61nc053UrNkVxZISCx13eNRYnIRGAwDEH+HeH9l5Dj
ylmQ53e7DoEfU1ar4o/ZZ1GkmctGfwbD0C1jXIVVl/Xbfn+sAq2kQvS151Gj7nEn
K1g7ISGaoYIp/0i7lTYoCDLl4INH/fG9HxFeXM2H5KTrmhyzIWsFmHKZkDkdWb0J
WuXmi/i62zLZ//4c+g/Udu9VrOqBXzO/kR4lLrEHd6W6kV+JFttMJmJL2naGPlRV
hH8fJQ+IrRfzxFhhaH9XHBwjFnxUvhoSBEt+3PSVPa/hbL06yGI/93q1tWZRODjM
5LMWcOSZwW39wUlzP1+afc5RvQPF7k0e6YvNZyRJSAAUeU2r45Jiil3j/SIC4Ub8
pQNHtUABUZhyB9a4LHyzZJSBRnqrmnb5JaNACJpNM8A5CFUfYqrHCTpWHgE+iEEB
cWlK4VNjzblHPADX1lmhqdCdRkVCIxDXs13m6yfsFGX5mXxMdh+tjJipTKGZVtCy
NXtbdD+A/ZHfgXKkxkFlXrS61DhMwZ44RIUsy3i511Uvvdbg1IBmuOo/mGCFPAaA
+f/PGsvDeLXldxehnDkJ89+sO60H3T6SeIHOpAoOW7mX/7IIQkqyDlCbLH+ESikw
gGDB3oh2vVRgtOnboBuHSk8bIoqMPRegwmy0xsT6CUjA/j8B20Byllvvln68PR2Q
LNguJRn7XK2EaQUiVM+tGs4aVPpJVy2KuKreQrtQK8K+fTHq3n/wfQnTz+I7UNmA
12gTPQF5+UImdKU5Tn5xxN67E7Qb9frIkgaYzJN2H+zd6oylJRcRDU7YO8r+anVT
5ZNBS5aV40dmKFCmm8ph5QpJ1AvDhB4zF4uRsOE+3W6CWao8ZmPfMM+4CHw72T6P
HmFSeNE6e9lTbtBmpJURSPPxV/jV8tUUzt9wV4aAPxDFTmcQsX8FRRL7lilthEnp
LFMelU5yt0a5WMtkIKvBU0nKCrY0Kq+04g/TcuYXvzvEzM5fa7+idQTKQJYlPKxr
RSfoElIBtm2tz6FMgIArVx7lKvJ2GsDi5A27xfI+MkQpFXdAlBqvjPVnDVU+wgvi
Lq7MA8hXFr1dgiZmgC8z4w4N4v31y7T9ujlAvrj2LsaRCOYap63J9Coz9ur8thef
voQzmhyzYgMYIhVwreWdCYsyxr8kULc6vRGfft+RdDh2/7NoxprRW+m2p4MKkLmh
OOijMMgeBtdNQ3Lm3XwgVcN19YeaTgq7riVMYhdfQAomDdIF9h/rvJxCkBrCjb+e
YZS4lqnhBk0K5xdx2M8Zn1cdDsmnniXfw+1Af1KXmOG9cPAsIbur4zYQqYwmiWYN
62qmDt/xOoeAXWwzfvyRdqLCHWr4HkNDxbX8XfHoMMXcXDvtwkqp3NqxyVIdDen3
edxDTkpRK7CYO3Nxb/SFxbFLw6dFaaP4hOAIYjir4KhZwX2fdo3qZpmCi+RzqwZ2
2Fc/nh5EKd/+yz5lokku4lRju1SSm3FZE7vj7pklKL0vdB4dVUu6XCksQTAbltSa
WhMdps5K1MSezimu1quOGFs0cGkeC4eC2d0GOMsQDeQI6RVGfbG7eJYwRWiGy+53
fZgvqf610wq/5bvtE0whXbbmjahUmlOzXa0surE1y0/3MkaMdPivZxw8yAcG3iiZ
PZyff46jSP1JvJRkoo2lBlOzNB8Dium+CQTi7Kfxp/5BMk55xL1Z6RdlOT1ac7ie
OlX/5AP6aces2Xj/6swDaifM09sIRm8QjavAzdlMucnN7q98rMo3qqtHXVjPnVaO
yf9eZt16P1f7j69ONHZ2fCSA/J9bZGzz/DXNhXbLOEZqIwk4i7Tziu8kkMxndkCq
X2BZmdFpGOem6c2o/ujiNsixmRJLqcKU+BRbFPv6SEFTf74rGRE6lffahC+a9/OM
TuNS3Z+vqqxoJypA3xP46DVdnJSQhgetNPieeAiUyQnFZT5fl3SkNG4Cd0A1pvkv
uMzYMwwqa4TFxIkul7GfNhd40N2nZ7ycxHVVhUYP4PE=
`pragma protect end_protected
