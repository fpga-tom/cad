// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rbfw8NtG4mRZoBnKFpcozmQcaqQMU6EkDMkVpQvi4k/fGJvK6DkgcewzPL07wiKB
24QKP6Y0F9RxN9/wpUTW8IlwWDZ+15BQglIArrvWqH0ZRGo3XqF7v2t4Pb8/WeHY
O8xodLrL4QaXl206UBcFQM1eLh5gQY8Jkejjxy2uH1M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4800)
RrYISlk6MfdOROn37DaL4brs7LeGMPnp11KDSDitTc+QuMoukkb2yyT2dI23o7eq
7MNCvnRal5m+zJefUnXahqDmVpu9GpgboRwIwlMjRbYbqkGy7tqlAsiCo1hulK6l
dl/+3LQ3iRIns4cM404VnwVVBU0LBWYTtGMH8ZfYw5WeCvBWijcFlgHhC/DWfASS
RiOFZPHUUn5rNkCTiq/UNZbv/4rvX9M+AckGt0OjL3i3o3jjc3nfmX83z9j5IPmj
QczKJKosBKFCYaz9Gtj+nZSTWvEWsB+BfRuOwEFVe3s6Id8EeUuxICqdDTXaB5Lx
zYAnXPIixyHiCqHcxBITFezIxZwhTEkbudBUNtnETRR9ek4UvvLtmNRls/iXRZNP
S14+zS1drWaGGdxukWQoHyQYdKdLmbICP0JT1sbwaTJBRfk8TNng+nsRekuaAiLE
wBhYKWajys5gb6K9KM0Ro0L9D6uD484GBhNEWPsuFQRFyV5+EwhHW8K5TTRM0nHo
UjdueSPzW1I7RY5YsAH5hvkXonAU6L8SvAqxvZbADNF3VeT73WHs51pWGehIrCj3
4MGWN+N4bifLqStKnUdiQbpmok5bHt8LNWT0N+Q7GfT3v9V4C3QZ430z6ndf06s4
/UvaWpp8lGM0+Mwy4gOPGK1qq4wLLHYofjIp4WIh/IC2X6DOXLgZtuefWvVX0HEG
alsKKhy8L0OjXPX+d7+VPV3JOc6Xo3RibEVWig6PiJFgjTBQAuHUl6jo9ccIRjoM
Ds4Mj+o33jmq904rVEC7ZZw9BUSQM7q+eJ4fALh2er2IPwRTM84eIMslMshRK/r0
NKSyeAyr62nEvzsiuSqL5eK1abWcysbF9TYO6Z3V7WMfjFWuG7gWqjjuuMRe7/TQ
x3hmJUS9XVTRXelq3qxH8x6nFsVK/QupimQoaa83JX7iiqtQJkmiS3oEAyrHbjFn
0c+pKsfGliaQ2PdFNsc8Sx2TzqOLEAcno98AglCwFZdEgicMbrol4tjrTCZQgJrq
XLtRMsL9216a5CwTIlAK2gUI2g3js9MoFYy7gHeJG73VCqz8PKChy4/VQljvsDdT
i8vDm+RuiKJBKkqhqIYnh0bcpLd7J7Xl1WiJUO0IRZzeyb3Dzyh9MJPlcjj1XDML
U8K67JoByvxkRVlT2CHuTIKUO34Thx42GWfGd1iwtXbfS6+y6r3K7b1ewtGSG7o+
gbtVAxa/DsJ6ITvXYR36CMsNN9MeOJG6J9j/7faBVzkIXM1HqYLpE1h3sKyWacM1
mQBa1m0vDqnH3t5WD4l/TizgoslpnCKOKZSUGlJP9atD9eeDjUjMTLqwgFR/aRBl
g5gyTfO/Ko99KrJnreAbTqH8PUr9/fPRbTiAm0p+LgpaIaXLZ5a7DJmPx9odDQmw
yLUSAFjPitpFbcUdyFm12pNaCEe1EQQwt5HgCwgTU/iSrZx2m1M8AIwO3G13HNxl
GoWUv5WQl2WIV7KO0Lj5ZB9lEflztRSukWp9RBMnAbWkkUmxl3zHODe8h0h29DUx
D+Z469shRZm64+klw8hr/OKAyw3zPlBKQyuU8ZVHZocBG2og5WieYeJ80vjcya+V
InQpFhfRYZs2GIKWt4ikJk6wbIoDeurV3mUk3KqBnRBw6ny10AJ3L8qA9zCjpI41
OCDU7VIag6wj4ORHejVdJpT4Hgh8EnRwuG5oPqp1ZDlguqsbdVjeHzoD4RqoZfUA
NR6hKiUOJ7MJFLlIlR7/OcPRkxA8omR+N+3EtyflCv7L2LGvi70DvjaxUS6eTcmg
j4huAYWURnCs8KQdg7uljTZyAapjwC5G+aUrDXD9H7D1r5VqdvY6TgNmnUNTaWWH
lnbBMsy1CCTP6H7ZL7kj9ck1i0JfqfRZ/jwI3tZNfd5mSe+ZZ56BLCnKYYqsc5y8
fQTtjKy+nmn5wWrR0Ef6qLLwCrHHIIMF9kUZ2fDQ2Jmt7uJmYtEvwufNqgTM482u
On6cp7o9ZjQBsxW/3OblG2jbJgw0FunpCpH/5bnO+wc4MyfwvImA0UAE65J+OjWq
/PPQAkBVXOoQuIjiP3I+eMX4vQs6oXnlNRU4nOlp0CZIkPsRzcTF4fcLWcnB9QY8
NkjHozlEssiDsiKAOQ0JXhIJ2kyqJfocOkOamBH/AzTkR19VPieMs2+iRSdXY/fi
NGOc76u1Y4YzyrdrC4YmAK81DL1m7JqeTjEbvJhPx0UX7q9FDyCcdgo/JnWoUGek
RFiyQXC5vHdckJfdpS68A/OeBFrpneBLHfXsAj2ap+GNjFWRdhTmO72779C/Jed0
urSTihnnRcSZiXgJ7gzHFsF+zV3E/UszaipInM+yRBmks62YE7xobFGmE9XAHs0P
5UXNb1Dcc4QzzcXbzFLAKKJO8qglNN3aVczQ+olfcRCmBJryss4GDVw+HJlTyHB0
S37obOjRS90t62z9Q1qSz8SipeTogvprXjbQJatz9xW7lJTLKiHqaZQdrBLk3thD
22mipIs/9Ku1J3mPcAkSm5MDYqeUgesOSMWfhqVIAh0ITaJEyo/f73DYtKFDnVwz
BwUZs5Tvpdont3G0EFOwH+pCJZqDv4AKdgxXj9ZjZDIbw6jj7nKMEZg7b0rIPQgV
KQx4Ra5afdv+ODXNEnJejgntl7XOpTEeghLEVgRoTdagXRGBep3Hcx7xsdpBew9+
+AuDgeElHtH/pVDCtcBziZ7TTyC0aOUQvAvjF3Q/ao9H8eFwnsIgb2/imd4XR9Bw
V32ujGYHKu8CnQyqhm5ujHIIp8O0M0WR7XiK5ivdZvCkZjVEaDs+d4oVznbeShkV
n+P/SYE/bAnNEvKcUyIjAP8rEE5k/tUuXD2XbBqLS0XNJCZ2yTOcPInD8yOs+0Rg
gR2PLwYwDl3ZLzD08mpbwdNLNOmkkumIsL2Y4hiX6lgd9/2eCtuNW3LjO0NKy0ca
w1jRo1vZOuZU4crsaitcM0YvNdtTWGKF/7uv6aheNXriXuCL2DJs9ltoddD/4PE2
BP+5VcXVibhJ/rJpK4FaITRNKMnQ7yWmhNm0BaXGTicj92zLd0NZwN0FxgI548zm
37LCJYfzAbsPYaY2Ch7vgoFE9zNHn70iJ1fHlzXtSZea0QjYozjmyd0ksIGG6keB
aFBpXJKTaOqkloeCKpxWaPWWFwgdicNnZEDHf++6Sx3IW4vf7ea5jZtZhGxlebWZ
/sGNtawm47hdPNHLWXGD310ZyEygqPEgzF1p0XTw6e4IqUj2AR6QgGb5hYZ/eh2+
T9EBYjjIkTC29qOUjg7XP6TDm5wTpByoffPGWZ83oW0l8V0tcnk/bWO+eZwDum9q
N7Nj8rVSq9xAbChwhg7PyuTItUmADLO7gd9FG6p7EzovnjiKj1CZo/8dC7z6WG2f
1R+MLB4doCcABfHA6gzIKIy6E6ckeo4Sfpp0jC8FsARdXsGk33dfgxTbpZQsY1LJ
HzoViMIpFkrVH1l9aVZG8d1F6PGPst68p1YP0lYjTVbiSYYS36XyEK0I1MVe1lcb
9dyT6VHNbGlEXOCEpVTkRAMX2C2r1/2s2zihWXuzVYiQTlPY0WJT40gNnakBcWrL
gYqU2IQ4Wk39eNlcT8rKB5I8leVBxt91a7leXXSYSK5zX5gnFJB0+XKKMLPUn+xS
/r9He6vwGsrbAfzOcIujZouuRklgI2jKyvOBCeHAjWeF15skkWOlhdaxGoARYVrd
MkcrhfhrU8HpKsD0YuE0enoY13zOossNvbyjyB7zZR46uQcayTi2VgookNU4SwtC
AGqC5MTg3Rb/5MF9B7xzQlTLbZo58UFEMH0gByGNfPoI7ugZNY0YXdqJR2tekkv7
du2GRlT6m8zVzdt1rO7C+q0y6GOjVe1mXwTjE4HTFAFw8FuPNKVu7J7EhHm6b8AN
LgR+n9WWTaZJ1TCSnSc/5mYqGtxiSHAkejCCmgh99qPv+e34YrmVWxb4F9TPvp31
tAl4oDdJjm3wnemdx87VFBeIYfRUpaJg4wm5yllgVcKgF7rMknhxuIqh6VGPkVVe
XyR2mOvxoQzUQoU5VUOfkw+sSKMbnQRZ7jMibi8igQVz/5jNaUNQbS/DhcBtbCdE
gqCfUyAiExD7gzU3sOx7m1MjB5QaTAiq6/e7bkqPWx601SFi9Np7VYLcZG2fdNwo
QxCI+wkuFHr9LXNAKeVr9cPVSplfdVKeU9xl02eq0mWTtHz8/UjtGcYHSSPlck1S
6diFbo5V799fT/4qycTwzxUwwXHa5e4q+k5u3uzhsTyA0pZaPo5cryoGLl1KWwo5
xV9VxfY/pOZcypW3kfLg2ZEE63IKB1UthPYT0oGZS9foAoySPr7mVFpD1uRYsKs7
ipWk1yIHNhqjz1KeNTVjgeYJmfI++OF2X7Hw8M3CwqLQyn7WRD1HPxJYK/wMbF3V
OCmxKu76A/wNmgAd+zNbnrzTTRQ16UJLkeF0WF1HlZg2bg+kewhd0McJ43uzYKql
+2yH1ka9tI1RIVbLKHN9f6NhW76ekoh0JcGj7CXwQXO0+yBOLkA9Y766HckvxvXs
nQD8pK1TrU+WrcpWgNdSrH+uuss2/07kQUMpPDgayDp8K1WO6f7shkFfGX7/sriz
A1rp39LzFowGZEs/71SUgpwdY8XaMHBCXIhxXLpooRLPeooNtrACsruOmqtFQ6c2
6we18IVKsZyNEMnMKmmaWui8PWp+GesJ1VuozHTPZguGzfP7Y1OhvTvkusERM/w5
Qnu7c9sR2252F42PmJB78Hf6pEluGSvBy4N26t33dk4DfS0qLIOks1o0EbdYZGps
jffQTij83ZHvCS2RZ22SCsaujdYb09vS0VueTutUCwS9Zxb3ZbZbbz/peGxaibvo
5eJYZeGTWedHl2jXPOjmPgfLylQTF+EWSTsT513iiMSaFznjBw1JN4YU2zIqaP0i
J3crYd13PqtU5HxF/q6xtXF5fgPVr/R0Ad9RbN1FiAGh/nhdczLnxDnvf4GEBBS9
NXC5fX0+DiVkboMfVqG0Cnpcmd8Ohx7fj0O08+CTkZtHIN59fpivt5QuW6PEa40a
wEHPbEnoRyD9BDUXXSBqYyiz6rjsB5VoGmxz0/0yiHF2jL2tOh15HdC06KRMzzNp
+0bvVTPpedXU7Yxxgin8qqPpyBYUMn8ENtwh6k1S+kjcpJpdOoait/Bw+EUzOoWB
4wpX6aTfvL7XR2R7qPfNLm4oeN5Ru+O8LE40e03FJ4ctMZOHNPVuav0utHrxU7QQ
Iz5wvCCsQmnPmPR8QSv3fTW5oOt2xCCYY3Nyd3EfaYOtUnma5ZrVkigZWVwoPI0w
LyvdpbppPDfTBQvfCL6w3iAUxOqNrPR28dnowQme3Dxbl/pjuQk2hrk+ESdz6Lgt
FnSoGtYMLNomtxftXdKjosBOMGLCoT1PNha4zoySASYBtDM9udmUJrAuUqXKRB+L
VR0HqaztEMcGRGUx73pZ7I8Xy1k3JXn0a+1KIdzeXBgJKBeJCVGdQxkJteM6Y9u9
q+9yFJsX+/ttmX95Yt41+GBVwHIdhf+dfccLpq5XJ9vYNGSuHjrZkiLCR90oX2jK
ytQNXDHVIvmnK1CZhFbTJ3f9TJG6eqiD4Wtc9QE95OpUF7ktWHWCX8WzBdqkoT9/
EEIRRSYYM+d6WS3s0Lh6y2Z6BqLzJhIrD8IxGBZP6NcLSS8fNcw+q/JRQWJVLQM2
m2l26vt7vpWD8hKKg++ecI/hqrBpK0YhbMjoS4rWbI5iHh5LLQHn1LQbS5bamp2b
fp+vXgJU5GLo8SJIsZEetM5plrSgEG8h97XOdNRBztiCF7GXXvHBUL2gTXknazOX
bMEBKLi7hzPLeigv3DEDfzk35IfJA8/wfwE5iAole+IcEQm7UpFGwUU5hD2RVVrI
zsfty8DXE1dM8Zg4ZcSsR5vZzVPj6s95mcJ8/UHBz/sV+JgO6pttKUa9Qpf9rwv3
qU9Yyy78VUuT0beYJ0vBNApn6Aat6d5zXh7ylBK55a2kOegs1MuURCyNJcZM71GV
4tQxMx/EgTV1jnYhBFmygFpm1n0dpbQs/aRfqBz51OoRMSXFySBSkyvaeFSgCiKA
jZNDHrD40WXtE14p6Z4ZBvbYIcgF00zR7ICNRpFwxdJM8dPqAKG9GqEKpSJFvBDw
mGZeJthWkQZ1Ze7CZOPjyWm4rZo58TkHoCfgwW8vIcTC2ot/+Y7Umvb9Tu5YkPW/
bNIdUZYyjRnoJoMEQzLjp3UOYSe8d7go3F5NJYvGKQZy+qhjbHLiQHLaIvSI/Iz/
mNcIlM1nFOI6dipWFgIGUrxeF0uUjZOFe2PisvX4LnWmdx1ebNXj1Hkm5Ed0lYVu
/yEQHrCES0G0bA8su8Cc1AKx7E+CWgYdVZK2Hj+oLJtyiCk/tRdj9tjW0A2WWjPZ
`pragma protect end_protected
