// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MIpQlwp50dY7pM74S8GUTKp1p/Vs16Dyz9XMZ1tBGtJo1v5dmwNXeIL9Afhp3R/E
doEa+l0GKHWw/T1q4dmd/SMTsN0IEUB8hqaMJLP2hGPV5Z3GV3f83bE5z9tPPqNt
egrw9c+Kw37Da4RJNpmw6oyud6gOeH9/H+SGUGsWSII=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5632)
nfn6kbf9HJfO/PkCqtJhyAuxHouZdoCN0KwzkHWg3MR17T6brHYGw4b7tUZYyXxH
ZrITCAdtKot4ZPuPhikA9wQ7zwwqYu0H6TvznzIcQqTF3U4a2A14zuAs8XuFIIOT
0snflH2vkfuADWpVbQlR5ARoVu1OZaA5bJlvs8nViJJyIuq+BDv6CRsSYvbBQ8hU
1yqE57LtG3qDtSvLHzHrNIP8a7Ja+BdmdxwDAQQzcQyzWyWLHO8FUafN1sXk6VHi
k4QXYGN2Vy35hPCX/ddqG490jfanH6PzGwqgrSxH6enqNdPX5lECgT3gC095CrZZ
cPMWO0M1vsuRdU3ODLjNAiTEk3tkk9mjUO9Zp1yzpbCmqvOmiSl7S7EaQ2Dk/vN3
2nmwiGAvdcLp3tMYSlgelsqh8rc4mi6/DmAw9JME97CoT6Gh5NlyRerZ1K53QZhM
r2lOCTFRo3luqTK8QsY3MVzavm2w5A3OimpgwPyts/5W+GlP6/kKvfr17080Ac8h
Mm5H289WlbKIgoRzaglFsUr6x2rKzbSa6qVZUxRF3bEkXbbz9Jr0yM00hxk5nekj
1KRthzg0//bRUDYN1Ln2M+ky1ZVK/Km8PXiRoR3iUHdMj/WM+3yfUzPWEDHqB2Nw
6nPOxnfPk9FAGDqmPw2X9jgRI2dE/x8ESSQijjiXPPXhHmJI2kDu15XPe3gpaCPW
9miRXpMdjNn3+IVqR7puZL4IEu6LoWlaR97TjAPz5cu9iRoZVWAtXSjlBYfx8RFF
O/33vAASco30gfIJrsACjAYgjjU295TKaX8nlidklNtp0FSOuOf9Og3x9GSOLLAx
ghjTJAsOxczfQUskgMezSwWqP9+GGcv7zA6TkJdgmOY+8gB+lRvfEtiV8n2gzann
dLbMmkpvUMqtvNMAFn7mms64SbTZixAYfV7gCI6PdY+Nwb83QTq/xVcH4woKrflz
eAOElJvsPkTtZm35bkuQJ5Whb6ucXbjfFw34XPjRzzfRgPwGszF6HotY08TYHP5d
Fn9T6MmA7Cf0sAPmtll/GgM5gBkM2FzvJgqQ6IDtiBwVPJ631yJDPCcx59ofobbW
ptYfyApusZOZEAwT+vgQ/lwqIas1foqyFvrBrx5l4O9tEdOF8uz+hutRNSyiwhos
mBkftO/8cD87kc0ZM+45chqUufzqYdWyl2mBkCRPdkxN55rp9xgwT9XLo967f509
zMrXm/sChZ9zI48H3fZvtAhWEbUACkuqcGipUFlaJqZ59ffsGzHR4gi4Wnp3bZLv
+eUEDMp16j42trmvz6RSge6rNtMUPtOycbyeALQq9RZ2RJGdOvPeIAvibVbVaJ0M
VURZjjiMFqHZbu2Jo5eEUnHWl72iZR/cZ2vyUtuYIcClCye9ZOKL3vEZ+OWIbog6
TvahsIT8iJGz4gmwHB5FAEE8w0caOQ6dRFMH1gVIDdBsCcvgDHwASOAB77LgyKBs
OWNzeMn/CxvFzDH7vFmGQhSywfgU5OGJouieSsRcfAqOmX628DChy1300hszwqbb
50Arz8dEcALSDEoB0fygAB/mzPg0gldxdM7XI5A49zDZObM5c7L5xNpzq5dRiMBB
53rB97A0cKiHECwfAXymh00j/hPTu/C+ZSwCahFQL2QyeuBCow3isfa1utmse1FU
9sFN50G+E6Jr+9F+VXtqoBsB2YcsiDl3ZXy6+jy5PmLW1gPCM+zx1v0pwtFClJW3
B7AM6m8xrqc0ssTuTtWX4AiQKXU6l7Xo/TQEGNVGuS7t4KcoCsh9RTbVexDDiQPB
OeEMZ8I1ykLcG0rJubhei93wQ3gHC7lsRLhbKnuSNYLzvnDxvn/qa0dWawsbQY/+
rYzOLZuKLWawglEp5XifmjVheQLZboCd8htBQg0CNxin/57ZW469HfgFBFjVc2Ns
BCHiFsb3JhYiEhSiKtkNoFhEg1Nee39pJ8K3dILcAg+cWlEYYb82Rfry4dBirpp3
eblBY0BVwQAtbnG4OAvajgMV0QqfCO0wzzI3KA0/1U+uWYg3Ar38EMIthejdB0OM
07JjSWRf462yWNC3oaaq6viFGVKi+Aowzcl4Vy8We9RiuwmP5iQ8XKltGtRPUnP4
wx/EIzOzKG68D+dKCpQBD41nqu92Jgzt1tdSHUZltml1UUcHt89wvjhD0WMkRz+7
ABwNN6UApK28jUzs0tEUZxFT63ZbGsPh6Q6qfOzQDHI/6ZIV963jzfHS7tvlmw9I
wEIQKpgmDBhB36ruB3OfnPrrPPJfEp+PTPSAbVxfq2ZyIE2cfFRnPmzPt81en6Mq
E4oKOoBIASO8oLQYLQQS3FpHfPx2aJ/1O966SRo69A7ixj5UEmBa+Jwx2hd/F9lv
xnZdffVtq8IaRQuE2IBqHycHGTzMRICIR18yOD4YwcuRU0UWazFuhtQioFoHKtaE
227iNzzYaIn7n3w+v6BV/WAimkOQdNqnOUxN+F4Mtu0aXGTCRUAaWrrj4fXPWC8O
CCv+Vu7pKbExjrkUz/vv15g2Kb61n2mgzEbQbLf6DQltyChRaG9+0Vz1ry0k7Kom
GchgJixvWt41+D1i7KcF0Larn8VS/fs2q0XWofV1vr1Lsk8vEiJXf2AEzHJiR02B
XNbiNlO99KmHeezGQUFlzQjX9NqbE6tHSxX5Qf/58ywHJ4oSYQWvt4tj0VAQFzt2
Aqc1G8PPSsRJ9us3QQh4h8MHshw35AeOcdBVNhX/bgdAQ+VBUayEmErDgVKnsBp8
ZsbTzoMgJSRLB2M1C6FqQAcyYALyfeRmOTkE0H9azZTXjhBCgPP51kViM+U4+kTp
Wv0sE/74YIwdF5QjmFKXlj6gcrV0RExmpoCaeT3R77WMgX1QnH7cgm5NDSNUeCKl
SmI/ZJtCVA2xDC9zk7SoyRegWAEAUwCMvTKllT+8nzQC2Puitd8nrZqF+/MR/Lpt
7hEekXC2pu0hnN5FVAUXqN5PlO1qDBJvhltqwxb7Bllh64X5udzGpDkjBfb43XVh
Nbg4gLYrxTm/dsKApIqO1vcCZSJLPoYTl8xeUu+5uU1t8ZgmJ9Yji2wmLxZVROwf
uAdI0FIzhMZNJUuNh5BHVsh1MuUXlQG9Xpm0cWVTmvW8qVlyWtn3VLOfnewtl3o/
gQ/uqiMGPxFTBkzInSXMbtpAi7v51f3FIq+scG/MwbdpfK5F3TwaV0JtzbasN7e/
UrKG4sMxy6pnW6HoDFu5ffX2ZKF1dIfM+k3K7G22UskiHX/cCEEk+esJIInaLHF2
fFYkYQP/laqXJOcxF0DWbi33B0bLn5TzA/uzWJJxrCCx3q+7xYJpprgAT1QLbA+L
zkKFhjJKT9SRprwOe7bIXO262QVPhiu8QQNyDtnjQefUnMsQDqRHxXIwVkUX0OPM
rW548o6N+B7uSCm+vbR1zxx5tb+6vvg3WfoNpNpJtxdBPS0GtCIDfFjCkg/XB13B
AvJBHbFA1peBJL02U94ddtVBneAFU82Yb8+vIewNHC95MwT3/mWhAULRMpP0+YxG
O3UgksSDvi2ehQtxiJkVW7N+BOv0tgP7yxQxdOScGzcrO8jUqBCQzi5NUHNSHfzS
YDQCnyT1+dtwmMrkVk7UWMKHpHh19sJceSitWXaJ0klSYzmNvLhDx5hJFzLXBt8N
bQx4BKQAGDPYahtFY6GvJxJLpkuwiWih45X8zH9N6GObvubYNMgWNcfqwikgL4Gd
PaE/O039134F5FD7TOJA++Oia450g1JuL8RbOxwcejMAn+MsbCSq206wpx3bFD+f
Zy//5XeslGZ31KLwoFyxPexT0+LGNFob43tn2gAiL8QOWJXiq4Ywangjfvgm7mdq
zKXgr8j1Z8tnyYgnS3J5Ketb8hN+d5nz6Ria0u1AUrRo6xedN63PZ5mD+gWlhY3k
kFIp+J963Nrn1Tf+JmVmFe8RKq492YXtJFkDX6YWCbsdh2sHBfbHaj7nsw4yONdA
IVbyCGZCdzY1aD8RaATGP7Bc/pJ5ZzOlH0ynBUsi31gn0cC8CHUjSkBxygAThkCB
1KJXwkbxrtwtTzsWQsG7B29NtGFuUBYPa5GTMEsu45rzgtLZ6GAmXLCExxeECfu9
3Z7n3K1h/HZFGZ3e5RXMX0igSowPG2w3da+FeCQgFUg9bhtqaQX93AB9NffJBshb
fPPgIzoMFNYNYcHyf/hNVZkvzwhPY7qf0TWKa8SgEmIo+7lpGHRQoCJxKhw0+8Sn
WS6rqorSUHJYqT2PaRuFIhzEAVZscpaPNpGjoHJ87C6RhQ4ah+fGBIVW3YetJ7Sh
H+hW1FOrqrEj3PfdmEQgOEbifubdvXq2E478IZB9NY5MR49297qqknp75wPrXfFV
fxv7XCXb1hSCk71RiQ/2FeIOoMv8p4mYmjmbioSG+IdyhSEP78VwxVtbgGd6P70a
Fez6ra3TKx79AJv2VuuyHXMHGxvmnIReE6Qq7CILsAk+DBVZmsa1dj4tXF2EHBd+
8aKLMARnA592SeHO4UCp6GfAEYIbPpphBI2Vex5He9YR9u2dgfQkbnY8vMzhfhrq
LTHYotuZTvKYAoNbSf72r7pWQ6fuEwS/lFUCKHlDgplEhVB86G8Z7Q4TXK9NkPU0
racaGQDEPsBxK93NTcXOaweEQC/X1gmPhslSwCZCrki/KluXGkzHhQcsX57tdZJs
+PvxW09T+K9SpiSexosQP2/q5m0fwQpUEpEiVNl4AMqO1Yrat1NbhmtewLpqCDQh
hDRytJxIx6uSUUEJonZfsu5JOCgoAlQXt9Qsu/1X8fQqnSrutd5RqFG2A3twn+J/
KveZcNL/TbGLbbUc0VTWzZoQqq8SAD6sY5aNOExo/Lbj+39QiaGyT4U6Ecx2qo8d
Vpr1s5RA5KeRr3TtcKqMmAqEOUlhrclGssB1yCnSr3GwxJwKbTXtxxwE+nvJIPlO
x0NKsHGfyENmW6R8nnl34ZhB9PuRbFPu153FrGoIgeYGvXjMgTVqOpwVkrux+xhT
R/lZEbfIhw5upTD20y+opnXLpdmBo4WGgA0Wbv5Nm73Dg+OisZCnJcOyX75+vhE6
RATjMtI/h4vHe5yBqpIkFlmISLQ0qscPT0U/YOZOuxzg883gpNTXBxo89/PYw8YT
km4cOTLogWyiZTf0+WZoLblOvra+r0XkPyIm7r9EpUgZvso08agUwM1iPfvvUd2U
tsrD56lcikGjsm1ftp6YC2cPRxjZBZYIMlaVQOMo2kVLWT6xBM2ba0Ei0FjwpKYs
k0MGd0UbE8uJUtFJw39qFZ4WvaNpfw0HGMKLvHj0PE6Zr0rNzfwRPXtdqcfth19A
YKk4vIWd/891nBquXcMKG1pJyuzoheftKotIQFRYkk28hJmMu26/Va1dNIl2UnIL
/vqUsNZnZb+L6ZN7nCfbrQ6/NeRVaVL7yL5eXlcgYt946yUCIpmlUw5LD/pT9Fwe
6v3lVagjElhFg67r2eeBfNd5DhVDFQic94bKI4PY2NwHXqgfQEb2omNmjduHa6Rp
ZN9nIp10/BwChFmXkXKj5OiWzdD4aZmHnbXm6dUlA6GYAQ1pyzt/XCq6TwHN02B+
oQJRc0sit3HDGXJFijmy39VCRFHjd/jONiuAZtPklAEIrEoUgWtcXq62YT2lHjOi
foLX/In9jO26SI/pA0q7uSPQPUU52fDxH2h7LfkW3v5+geE2cB6JbD+HQIutbYNo
eZxohacvXF3lPNP02bifO70XOiUEevuA8kvX9ryV3sE4pwJ68BARTzUFqO+c65/S
X2yj1aoxMw2KFxvM4icr6WoE4zvmFuqrJmSm8q/+gh1OC58MiUNKQtc53hv/lGz6
r1mdSs5Rh0A0QHEJmPAXQf4yDjcy/n2i+EGvc2sem2FoBV1mD5b3zrFpmnBR7v0L
wrQVDvqLYN416VS5WjRChzIQbItNRnHlBH6Yo/Ld0vzBQ6bCJTqAsvz1e0mCnBvc
iZiWnGqa/6mqFwAN/9g79QSxc5yWNh6qJdJFrKwHt6cDcy23PlS/CPdEZv+Eujro
7/Yugsy0Ci3RSyPb3YlyIyyBcB40/uv7yFrQkeOx/wqq08MkVQ8/J7fH0PiPap/6
aOC6nXx8cLc4IFlpGQ8eXD0H4BmVZ4bg9IFX1XTkXvJzBbppCjVjHGzHKISwNW7j
k4QFxRXcuoOihiDevOkgxlVoS0+ujNjjUd90JJXvsC4yVXnB6CfLPaAhhkOKne3k
OKagKArQmR3LQL3l5UqOxWvOUtunRlzP96ePXceqSHiIlF1gBsE/+C9RVpt+7cmP
KW62v4XShk1+8s+ktBo2JE5eH9BHbBSezxO97so55+LNWTt0IfoSLLDIcLT1IWtc
I/eEkrY+ntVnjL9JqMRin3Xf95J6NqbkMsH9kifLqWn++tgRVPxOu9lRDbj+S07p
Dn873N4IFHhL7QRuUfyE5ZKYvXvhmbzxA19tgJahvvquUMHAihwYXlqOGDGADH42
GLeqje5BZo6eWnXLiCUgMIkUIgBJb+VAvqw/tmoh1koeA4O1+QHbt7a8hEvfgjFn
uin1puhZ3W+qaxj2zVWy0UkgySbpsD+cnr7+iL2yJdO5BU4WA4KM08WyBIpRDhF3
8cXkpyGmDRbhXYE2i4VwX5pkWAR4Vd2IOkK4ZN7BToJMax/1B96PkwsxaEFLHGP0
MtW5T2laTwYwo/cF8qNZdeJTbs4Xp86Hm3aSeQmpmmKHLjYil3eqqv9tQ+tEg5TQ
YLNs74WwTrvP223LlfFrwOfmUYEe/1zsPJjoexDL8I0ygBRyqWZG0uhm2iiuGCpd
10hkjwuFNfQ3SU+VCUWHaclufyCgoQ2X/trmnL/nD3pNeJwu1HJAH32ya6KG1v6i
HGQODntKidXt3Nd3gazywN3gY3Ku+hWQlm4sdaHIpPgMqYW4IqWabZ+xMhQeShzX
xMT8DjRQT2urss3tSSebeR+sIrxA4XUcYecDqlKe4ZTtRplDR4aX86PGYTtFORIs
HUrLoAugwbg4s3RFz5KuG9ceK2GLTpOdD+B0wHTjIsAFtTvzce7NcEz14hgnE2hB
ffCvZlcxpudDqWHqP8WfXKZHGjpRvWBm5AocaY+N/af3bu/vjOAm4ZZpHVbdbToS
cuYw1dylf/ekoiDT276Db+DIqLq9sLTKzqjTO3ras7+GLhEm9K4usn3/DLgjCGcl
NCYg0pn+JeMQnJ6XtSaVbOXx52A9YSJxr4V70xL5lApcbj7YzrMSDjhevqOMSV2c
+AjAXgJrr8NM+FxITJrUk1rB50GrNKdvM3WIqq15tPYPeCOUR1SHD5mga4hAmh3Q
ajxoMUY6D9v5Ko9f+Vt3sAxzm82UrTmQS7c0oj3RCycFBwS9/M/MCnJhLEbIXftU
Rq0zNSzoGebndq5l6C9ePbNLu7woKCG/zudSFIVkOMbWS2w3L6bztW3AtDp1la+o
A837nbm6tEMbCiHXiixDmgywuvNUPtfFNUQrkxbbuemMSv0DkIXYVar3XkJyNyKK
Dr9pZB7E/VUmqInpxTIVyg==
`pragma protect end_protected
