// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:49 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IAnEN1M/kindTuMSZk4FVuOB7tlarMqGXlT4qF0XZ+YPqopdyTHhEd0/6h1qD+J0
ztGVDCOLS18+7Wxhxzn0TwWmVxjQvFJfab1sTdZtRjNL+sJV7zqUUvdh0p/gceaD
rBqbfNTULETMecWlx4+iIr7UDgGW4rdwlt1mRfRw9fs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7712)
VUvkzbuzV6gE9Wym1TOhS1HrSHjS+Tlk+dkued/fGf/wYt1c1Uk+2CgqXDOKUqMr
BenzroWFZ2ZRJGR4cpvUh691ak0afXPL4KWMQ2z5uwfEvXb4xIoNgIzuiy3nE7UE
DZNIvi2/YTgy2Y/rea/NhLPdU29dMMFlca1T+PTOfcXQ7b5roM0mWOoKMCzH3Sru
Ch4VhnQZ1rCUsgSsLG6glJ1urZzpHtidC3ySCQM9pxdCgIv72O32xiDLEWKfaNSU
MfWONzkYDRWCtwdRnxZWBVKvnKjeqTC3oEIwLPpbCXAUYZrfJeugL+8h6bM+J//6
nfe98k8QPRts6KEAEUjjtroueGAWGTONw+Zdb6dwjuswyNFhD9xSFXDz2itKDMZ7
Q9fu6pv4pui2Pl6cINuNSxNXaV2lSyv6caqHvQQvhkF1/4zOotzemHkuxvaC+Ik/
5/eImeI8wJyqlzyQolrgiluVelx6n9942bux8eZJ90EABJfsPdvtqz+ACz1mL5co
zSoSTqjleT1zOexyY+Hhh7d3whYDq0r/VljWr8V4rPSQ7w3xaj7qiG0o089JbDTJ
a3EDI+2HLsXBcKHa93KgRuDWBa6g6nkV8SZzHtFyNQZgoUYAuJPdKuEwyRu5KDvy
VnkrJX/Tkoxq/qpssrVUZIdjIoXWrYp62Xu3JzocmNjBU5A/f7cnISNc2rxA9ZaR
pAw/zb8jZ1AT6pLBbU1oBjCmvWSeeakV5Ne+xJlTMlBalBFCLsQGl/zUat0QK2s0
vAUo0ubSvhJaTWlGrfHsPlbttKqCqrAYrEIAs9SBLp/k6FWXfkZiYxxLJIexl2KQ
frVRw1565SCWPgH7Vm2ExvmrmupLxGg2Ma4N6wCxl008G9lQ2KgJG43LL1HvnVDT
ThF5GHPMNjOJBcmlCtVaWkh2NJ0/EQsicDFDY6pysspSwNi7UKOw99SaKG8pkdoV
infw55v6iUdwM3u40uXHFHNr7Mf+m1pcwvvU5uql+nxU7hLtTDvmQl+VQLbn7X+D
SByd1d/1V2UrjczrcymAigBzZnw3aDAWeTElOahUHp83KhFnjtopoYXW9Iismvs3
D1vvwLhI6bQwqbQ8FDZAcaxPMqLak3Ls2swbmSLxuKVm/fSCvFdXTNZwn7X63AZX
AT1G90PQBdZUtxdocV4UFPLx1NQJzoTJQtybx/N/aVPIRkOoOPHx63eS3Vp2EiM8
CDmFol2Qz9zijsAuS+pvmsbSZIbDsMIac/GBsabrCcGFuFz53RKhrVJ8/lwfkfL/
/mILXT4JZ3azO9blke8awq+ui1vc19kjPlay6Tbayj3BIuaVaLxz6RLMEAyF2HWp
hqENsXWW/3R/DoofWOV1UTJIfA2UF7Z4fuX25J5LXhX9k4M0zd/3YJzvUnlidjGM
5Vn8Dl1CXHuUz+uO50hbhR8XSz9hlJHRRda+ZsPCNyfY1x1Xr+0632F5GDARyoUC
HdXQddAs2JtC6CvHjTQcvTJ8ekyuDI7+9VyLLShz17on/4OsR9yDeChFNaU4kxXR
Uot9y1cNcfNgzGRLSyK54hcFNKCPVSpohlWYUxE9+IzTO7b6gzuJo9k35xnfAFP4
tlDSVHpFYC7dNcF4hpTGKbqMV1fHvOS/cyud39vinyRBuBfSF8Yi5mURZ8hHAvxi
O0YoUmlhablG9W3/FTeR846qnhrag0xLBwRs+eqahmiGZRU/+7VXvY4+BrVLNxtx
Xlx2jGYHDoaWhnvgSJLzDvzT95wPxl8cDPUYmRanCDUN5YaGie8QPyfuxn58hHnE
RzRxrdCF9X8qenAcYMJPMoPdpsmTweiw8PutaZhjPayW6GqGN8idLW+/A2Ks1G5/
MaRO6RDdNKZJbDLFpeJltxNtQTi+nAwhoLehwoqClDKr0ln0qt1IGlLT33JfljFy
OHOIMV0ZxJ8EEFc10IMWUa+BHrVdW4cndUr8PudOKIVlhhJZLYQOqBHSVxmbpThl
1oJDy+5gFyIzy4cWT66i8JGvb0QObV0wixC/W14rtIAUWuD5LDDN6cLSaeuPh8rQ
F9BfNQ2fE3aF+Ylj93164Uqhsw9PzNSrDoOpLJO3CC1e+d+VhbK7Gacew0o4xMhO
SdwEYH++JEkaQl9RPieuJutOPwdvRPEqCCH++LiYN9ipZWetx01yway2BFhl4IqW
5CXDlkjPS0ZYauyBFBajOmeuP3J+un/04/nj9JfqIJQJAZDnuSfDZYMYJ7OIE1Jc
SYdQ5efVI7p7M6ReGw8EcWi4auZtOVcwzooFBzADMyD3XPFPuvPNZU9ogukkm3rw
C5YkKTRGAjEQs7thfK/Q4+jPurv2DI4rHyDo8qr5u643zpa3kJJiO/xuN3Vvdo4e
txhnlcCf7xiC9NagdTjUKvdf9t/kVJVduFAwvv+RlzlbnQLUn0LhZLZTbOwxRcc2
RVoauL99y+ZYWzBzjEq3pPcUeR694L0V73ZoK81S+3LxQ2r/OG45Iiwwb+l17a+D
jG1j+cLdvTDPI9n49DXJr18Jclt8jlyrmGow7TPrzXdjmeqhOk0eB877+WG08uaC
KvHpIfXFvHearu8F0ZMPJQ4z5134wkjdUN4sYZMKD5ymwMlxVpvVvu0pQejHiVK+
IBSKUZRFxOgl6mQAYaRkv0hdpluCGITMartoTdA+SOF/QNLCHwV+eGPDiM6iZSNa
UQ6nHIMV5JoaG1DvgYHnmeW4KaLGOSuZi3QbJt8srXTx3/T7gNp/LIU30O/lNsCH
k9F05EnzpjdoT/9bdLq1IGFsHjnOgAXaHimqDDVxKNl2K0CCiC/7qblagWYcbeWp
b0f+04W11hebzWtBoHaSikTxPWELjNSHMpoGUYRx9MQajLqCqP3F/ae4ltcjyRAw
TYL2vVWeWRGNP6HUfV3CiCCCZcTnNe5dr56qn5DQ7rca4vC9X2oAfAnTm7ctkDzu
3zUplQdzb3NdgABqXrkZ2rwkJG+0G5vHtcNJPtqffGs7SqIxo4WOrjZrbmCviJHP
XWdT9WcKLLhH/cOqil6qfSRV/bvStONFnQ4WjCYGnVSmoyX8bVQhHpOnBDuv6o+Q
mGof2N6ffV7AN8OBnOy/owPNb10NOmGdQJy5jQW1ejFmSJ0Rc3bwJM+aZxFe4LWx
ueiCK7mvugI1NeK0Xks6x+o/2wNIljIcQ79A9T7MAwyLWkD207ym38/HUMyHBdeP
i0n0rwyDZ7h/JGz0EwbOEFr5y+WPpqBOW9FpSKImaLvTo8YQddMRU6zVOxTC1o4j
7LAG+o4A5zLzkzsLi/HNEEUpTOP/lCdc4DNklueh/ZN8EkEMqQtqElLX/AL+mWA9
5KwVHEwOA2vNga4ni0jWe5cf5Lg7gVTFEZUV632FlPcX2hx1jrkPfohmIa8gnBSh
y/uIYS1eRWGe6P6CHIDGa6kl2RfYGToDQj20poljd6jur6e2PiWLahoVu8swa0XD
Sukf/s84xI7R+CmjLW92kgVdcxA8Sl0mdzwoxz7SoWLbBj0RRwPTdZ1J7ii4ABdH
S2lj2hvvkA0zZI+Y+e/5hvvspLHPrraeonnoYcwmgbINkkjAnj0qKyEIbF0deY/M
n/WSIExnjFH+9zRCH2s1LQTfLErHiAGrnxjTmwjkg02GC08xuaHxkj9mdgishwPo
I6fPVGwjktUy39G51SaTV3UZ6+k8OkXh1icBGByAN0L+bqQ78A6utWjr0plZVySx
H0eLef7L1+gIE1Xj2YmAvw2wJa0j4NSlRx/vAOayooSa+HXEdJ/tpwyQ/zQcRnkI
P7m2dm7kj6hCYPApgmrkLDIgzj6FYAvkmZ3awa+kPyA7tpEEEG5Cp0nuZSwlP7RV
bNvtAhxVqCyX85FBBMtdVoqgjItu3/JAJMdsAq6Vj4dcqXOnZ7CuzBljnG8FuMEk
h8dIxJ/IiqegEGm1IxbL/XemBpHOGwgqdnNUH+Fbz6dBJPx/FfICNzj6IsYBThh6
SuqwwxmUzy7klHqAd6INCLQHj095CsScce9jVFoUI9Bto2obI4MfIsmQo0QmqXf0
WyL9gQ3c4c7aWc0WP8rsnnj9kJd7mcK6fIED7+odjsj6GVdorncoE/eABXobJvLm
kyrcoEZTM/vkcYayH1g8j5ppu1qdTWqd7lG0pijua2XtHsHQ38GsHqAnPtzMFAyM
WXDtdiGL91EJ0SIAVg8LXfPWr++nyZuFt+7GHg0uk/4hFhN21pVcb2FXtWDbuk8J
qWSIl2eF2TxSm6IftlVyHsdqp+3ogmiFhozpRqGv88YtLPNO+l7R0ZLJhF+Mee64
/m8ok88veXUo2Uw7nZoE3iTBNxp9XepfdVhVycbOd4FvMbJ4Wa7uofO1TBkACDfL
VO/90HMoYTForUsgMJvY4YFIOdkNbbLQJuY3uQuhEqsUGCSBvoMjKlY7xoTP4Caj
oPA4zczkVOHk5vnmUoXaPUtA+CUhPZWN7cxpXFCR+lBXrCknTPR6DRNID1puqwvg
U7TLslozto59+ZbpkmlSi2R7/G5Wt7FDrgiVIgEdBwBRxWmn9OL8M3rti7nji5Kg
3TA2fhjUULL01/2LLkFSVEFg5R8nH4sCd7vmpggpxEwHa3AvlsOLT/zVIPZx8Zy2
X+zr/GxmsTmrk6PacmeIS4tPG1qLsQC7mtPndtj/oXL75ixKgsZqhDxa1hDkQXZL
WSP2+02YH2fZXsFP5cOgOKxuRmb6SPJHa+vRkV18vxA52cuUsOA31IqRgGsphwKr
ySikRL4GjtkB6YMP7iH+OUKz01YRwD8NajMQCeTi8lxTe7NGwGVEGfnP0Ld7h3FL
TdphjlhNrlZSwOkehYET/5B4KeiY6h8Y42UvwoHn3ppsCGFS4OgC7qhuWJihTkG9
cnOS3EjGUNGERThU5AFuI2PmPOOe73PpIbivhyetH7mLJqyrF7JmrzmQPxrFQHWn
1M2s7k4Kg3iYDUcjI+9xmWa2eslTjpmMcEHd4De7NBiIf+0NeuQ7Z+HeOCCUStlV
7VuGoVGkDGpCAHRRJkVmHdyJIWnB2uaMm26QyDqaP7cgd6xwfhLIyb4zj42sJmzG
iSe3SJz++Os0Me8CrbK1HAyhJmM24+mlvVI7J8GA8ZDThTUhyWLhbOztuLOYHGK6
5cSbdXRn3+OuzQUOAR11NC121/vbBuIRhJmX1hkfZDpj1SuJK+1gjvl//9e8aB/1
l0Xy0eT8so6x7JJglplqRRU8Y749CZDXdwWZ/ANHxcSBWTa5YLYUlSsEzi8+RD5K
17Q/FK2w8ckf4ZUEqJBMyySJtLeuLZ7Sv8CWyYn6U0ZRkxgFnarh8CRn7n5TAfQD
rBgu98xakG3YpegBhidawuB5CGbdsC61GIghmdaCyIrT4atSt5Qf97+LjKM192gg
cZTSNWAWfxK2K6BHRObDrE6G1x//h6YbTAKDTjwIwXDwgcDgbxCyyNLL6M/2BbKG
I78Co3u/noFV3gtwjji9KGfP0P8Sz/PHP0Su943Ht23k+h8/c9BEvhaR7OAvgVA1
y18xwlHK/x3EVYs/jhSJnYKDszaBF1oFG3W1rNmc3lOOaU23V0Jv2Y9m47F05Iu4
xKzCo6j/+RiHj5si8QaOrIlVPc2qnXrpiteKKsBUuW0O/ZYVhmarRC2950wqiKKJ
lan1UW4sesCPPQfmeTpz3d0LheW/pGsnez+hvpxgNYomALnMcFaZ5nRIbFH7Yksb
MKKSfeJZLybiCzWVP2UrVijJhxJ0UgY2o4U/pYIBfvqrn5ydLzysJzqSbE3/o4Gr
rQ129pXiUpJRHlsTlI2+0odKgUk6IA10+nP2jZ1sfvqqTP+k3FOv6z/tEFnWBkzT
ABIr0mTQP7WovTD6IQM9hzZLsqeeniGhbBwMSU0YIvj58gaYII+xXBuiWihuHR31
3qUiN6gb9+5f3qbQPiHEA3NKxxCXG0DTmSIzsaDOTF6Q3OOJhcDQ2PLB5Oy+s6uJ
8odwhpq2QQVAKubsVItBPC+VczBxnIMhw+OqQgaJjIuYHBndb4iY2yLZxs/DDdzT
z+l3y3EdPAYi8SHSUqScEU0Ufz4lInpwGalixflFidPWQAib2cJt/IhQKDrCtKPC
YLuvVlp+O80C9vg3pI1Hb+75zRXiWXnEfmoSfcdmyWgOmpl5JFlmDUiA+8C6u8Y8
Tfb3+Wkg89aIArov9r55QasitsacPxoyqf7nqWARQeNsDJmD4VsH7khJGYenRjWY
muGmiDSIDem48VNmqeBrppJBDzjdwjKNAaQahcTFjPbnByijqk2y/Mq2UA2cI1Mr
Wy5jkhF9+zc2ZE+GgyGZRrW5H3YbBOc1TmLdpxT38ZqcBFlAjPSvGi4rcJQSPKU2
JHarFuzIn11Pt2PLTLuSwwCcPq8UPLGkoq8ha8bBBJHiAI8TbNkrRLewnvinN8J4
nnMVNsu6krepGLuLO9bvkGFBTIWM/28atcEmpS57GcuzKX8yIPDBFYVuq/GHnNl8
s6YJ+4RgJq7WjjzjNXtlAjCGBtfouDzNJcav1Z7BxH9rZq+MNqFbRXpkyUbHwsXs
WHvOV4IojHE6NcJw37cH+4C3kr48QoLzBW03ISMg1XIBqZu3z+UoiRC6ZPBPk2QJ
OD0HWzt+256w07oLFVA0lV3/fU8087hEyq9tevWFCmmgqV6l4+6tWjmmlEJMMxod
WM9qRU2AeiniOGZI8/C+1GRKLVjEb7XNAfqNUvxMo9GA4C8Jk8vUgCQ2JAl2m8fN
1WrlnQrkYLl/a9+dWByeWbQPerL8DRdprpTx4EirIsS2SiCg5wc62DbIe+3hzMgT
jPb/0avkvoroqDhoFM+QjGQVcZGEmxxWSD4BFbptxKO6gXd+OLljeFOo24o1nDBQ
/4YNJyJn8Q8Bmcgs8XCgW/xaySch0npRjnRcfPqUEzJdX3UaeBqw60DsJdbvyJxS
Pikl2Su27lKOYh+jmCWBcmraJ2AiSbLAXOSPMIl6vVb9e2U3NRvio3PhhiN/2L9y
nMnQIBgWN7/EKcc0E4bdx2HscWF3U9WAJdyEfofCrX7q56jVLcJIjLJg6tSZYZRQ
k2KXutXqtkmFyaX9cPpMYGWHUNH0Z+lS+Blbe63BEaexAkw6xLlDz/U2rvk9Es7p
uVMoKjyoxpSJqj9DP6o0uy9SmUVGC1YXcW1TrTwfE9u1o6C/Y8SdQwVuP/z7/GVN
SurgMz0qAcjd0woiNh11X/WFNN9GZ3M6RaRGMgvp3YeYpNVLHJBe8IeK/tGuUTQK
rHNZl0K61biKkhm4oXfiKHZp7WAu+jazLhjHSW80QqOMlbrUrser0IRpE+6bdOev
cZkaZUfNO2PBerLRKWPgOjucx3kP8Yw8LUW3PlWuv6KWmun5GeXy9uyb3yhOs0rq
weScEKfu0xlnL8FXpz4YzuzfLdwgpJk54PkDvyujpz91cC4CiiGDYzi4mcT6L/zL
FYCIAoNtvgetwk+Hq1EFQMLUzbK536PVRQpAw0A3+0pR1VTmD6Yata7miHgaDOmH
2SEfzIJmDdFxOmCulngpbNKR3BS5Gsfw5yEB/aCYPFDNh1qOkUZClnGWh63fSYTb
wzt+Oiw4sI30Ocb15rbM4YyQMGbg7iy9VcqOOmyDs9BdDzKR1aa+YxBT7EUrdKcN
dDy8Ebr5HpHEaK9T+990aU+K5IMrgUmQMN7+WkVG4rIKWEjwukVU/lKs48b+mhtQ
3XzKqjcugcv8iK9fV64VnBrzUbKYaKyWeJ/5I455NOvjyVJr1lhY8tjJSdkZCkdJ
lGSDeEDBpNeW2naDMNFhy69R0JP/L6rKLg/57Sg1ISsCaPTzInCq2+Xqz38obfzJ
VuoQ1ehjDVe1+muyC1o9cm8gN3zx6gFOqgFKG57x1GfNquNwExHQb75PB86TkhOY
WtPywQpEB74ghPMB+dpdGPTw1uZTTQqgtgoqFftS7vOq86vz1A2n1Kfly02OyK+3
y3TX/QlgVDGHpDHoXXl8pOAgI7f9S75KohUYJaHL17+KpE7GSHirtCooWE6V9iJz
contWlnkj0StCEmOn5buhHXN+pnRjiw+EdGgSd6m+yOdkxH4eX8eGLT+uitIdD7M
4BWGn2f+Uq3YQCcm1XSeY1wZOUjpfSnRBC0PMd3847mE10HTOHT0T/KjPIyUFKa/
QFilfomYXbjHOdeokv5nhBVv0TVQ1qqseDrrtdIzCswZCqhEazM31Cc4+liMo1Kj
6u5RAmm8OPWtXqVwSbt/fDb07ICG046yHtH9TUMoiwK/d22FdbgobMHXMay7gnM3
V9INqxU/Whd4L3JhAR6sqVnZnifIEnZLvDv6BWxqKYDJeNwbDsJH+I8eeIiH2hcC
b1RwXNSzIHUK9cGU72kFlkms38bfdPjVpReO37F4gqa9hX44yxQ2xWj+LTCK6sUH
gOgYcpftyz9A0pgzgiFOYtmAJpj550a71NcSXiYMFZ55yOOPekbQiJDdNw9WDdSR
gUMLaOCPvnuisSfvGV1a++GwZZstaIQPRkH0wChaywSICD7iVkOyaeVAKSDZFHyq
ApzBhGqY5B/BTW8KEkDtIqYNwa/Lpdut12i3L4HYlYR9unJK056oPCDCD6GiA0Dp
c+habFfP4Dq9vNgwtZ9cFHY+gkNglAx5Kp7Gq289bYBFQIWMEggStulGLQicsr/J
Dw6GDGUx7Jqi4XqenR4qc3GpazvyJiNcYSkHe+cDtaCqdcOIzV0nhRDl8n90WLjM
nJlC34uZrshc+LVbQD73imKNDRBkP/ybryJ6OBNxo66Im4FLEq+Uu9x06Z0AZI9Y
qrMK2eZYDnoXhn2tyhHDh+w2ujdmP+/9nHPAg3viLsrUCGif+MzIN+BRPVpEFgmO
7WoJ0u7QKBAbWot7JLXUZq08+uEcP653kljXHluMeil4rVHCd4y3CLHd/AifHPVI
Y6k0s2SEfjEsX7TcAR1LmAWmErmpI5Z16fR7VDKsTmnxt7sG2BrC3qxpn/sdyD2z
g1busXHai+HfdwSEh3/UoLYTsWAXG5wpzFEpEUM4dQ/vC08Ol55gogAoARYBvc5D
XgYr7/BZV/h/o1iiY83NOlexB377g8wPE/nPSEp7PvCFWOmP+TYkmCJTg1agowTE
JXOKABefvIdk/t7IztPz2efk4a4iO5KkebnZzGl2GkHU4QeAc7FYTrRRIQeu/aFU
xIH5MO5Ed4kyQkFYiKmV3Minn3TKcxISXv5aQO+7Ryibvz1HzmuUTlcp4q0a6UUV
2pGkPsf+V9Oo84kyiUDCM/Y0r/8yeSEcFGlwSEFqczCujT3hZboQI8LrFaJU4Zmv
NVpbU0mNxnv+LNv8JP2ymQTbn6eAVbZdr0e2m44CKOMePDbc8PSZvJW0/1iniAF5
UjPC94a/f7oL75YlR0ZhJ44GIYaAHvs2DXXVM5T2xiwcgdqgEDgGxtxHeo48n5kQ
8GI/Br4b7HwRwK+TrR2saaa/rKk6Px/+dFbfrbFJn4qcZRcA5MjCPgLsCq/Tmd+P
Ndfej+D/S0CG0QoHXPo6mRXoID0J8CPzjCdwkSl59BEkCy/jMvXRgSv0fhK9/ka0
nsE1imPsRETtJSN+OUhBBINyH3NbVrE7M6YEKNIII8QjTc1q/6+JxrPFjmO6vurM
WDNox/iWMOEfsUdbIFF4yWEuw+SQ8gSLUz+Z0j0Hh1Tz4u+GO7uqjWC09NsapNnd
CS9a3S926bqmMAZdeBVM2NDBBzLvRnZqlCI1e2OeajfrOqfdQh50BbbuJzTUGsnn
XD9o+1no/mkWpEUuwQRxI1PV306JigwurV/kfE5BsDPYx7TqWF4geKo1ItiA+Slf
6Nyi3Wej+Lq0s+8vZWpFTbDJ7YbpzDia3x0nooFFi6MprmMzKE9XueVhdjR7GLgn
bXYd8whU9aro/TIU4h9zl7N0pyqrfwliU6LVtNoLPk6JNwa4n6d0mBjUSyitreFm
nvB+nHd+gdXS83Lg6+7awoPijPTIOZYCR9acYD1rIPX/99hlDdRgK+fULr8a57Ie
KpNB5DRlpqkUuJbVQy98Hrt3lE40MbWv3uLhmG68KjTkTNKssVHyu5ES84+EOqWD
NI0M/b9rsKEOPUUd6RIuzU6OZDoFXtQLckoYuYomlHttLbT43EklKCP/TBkTf0L/
fQ0oqY2AGw61NOlifL2SA08EVrBW5KUySR/0APj3qmy+7xH4LV0CDW/p6+u7dj7T
p+NU9ldYGvoeZiLqWUcFEc85Tb4kOCwTl+OpQdb/LzOK8LCARw3PRcADoJqwtEj2
r8XLBQvXIVP1gsAoQ+FkPo/j7uSETNB4E/XgnOiB9eI=
`pragma protect end_protected
