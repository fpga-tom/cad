// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
djAI8hVJ70G7YugN3Pl9/vP2qmmzNua1aiHFaH2qcZ/AboYz1CKKBZ9BRlXg3ny0
vIMrMfyQ8RYTSqOth+tSd3PpxTB9UJ+EBjtEJ+AI50aKV/F2LIW/O8zXZCzvhBZA
rvJPm8jiyiYzFczkq5VWPzEGIcCACl9V0vxmBX8mP0c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11168)
V5J5uw5GZrJrOT5V5MzkB9mRhNLQ/1ensH3YyW0CRpr7jwL8v5yrqbKDOyLN3l4O
4OiIFeuvcfs5bJ6SuOexURNiOAOGKoOIUqxGmRyGNAthvJUC5gtJ5q4sJqEe6Pnq
9+lmnvNP3U75g3vRypojJih/unEDtosKIDJ5udfPJ5vV3c7UOCgYpMa8yO4/IwzY
yVx9B8wlB6GxcDcY/Er3z8OS9yMO8vNCwh0bFniqZC+TEI00B/ujvxeixbXhcAlA
y4TkGCY8JB9GI6bzbvK12PNelyO03rx2p+qLjhA8SvK5AFEmuTWr/8rEL1/8NgqL
Pt+MM2Ei4E/OyWrG8OE5ER9K1lRKPLBDgK0C3F6csp4kviJgNzE+Cv66G1NX5QTO
O6f3ikJFxOp1IJ2UfWqOTAdW82CP8GfOxvpau9ZwIf0fxTw7D8nOvyXcsXjfNlE1
tDJ9YeuSpUMow6pliw4qsmWJPfVanjtWKnFwCw2t90sViIjVbB0UTjP3p6nHoKV0
lkNNaWsRJyvY1b4llWtLSkHulq73+VkFXAGzKdku8i9Z9cUy2jrf9K4qk/AJ3htL
mMap8p+QnuofbmfY+aFrNqZ2vQ+rBjCG2RSTExmA8noWaPeAv/ErXodHyUn/Knqc
oDcY7nIuVdbgDq0ROne5vAbZVw1wJZ9+TOfJHz75MHPPXjE1wPavV0O3Fntn+RAl
wAIDKZnpVwG+cNukUNTPB2lPr9USNiwUbTh8ooZsO7+G2RHbxbVhN/9PMvPgKleL
2aBPk/0cIbMC1wHQUWuWEoJpLtKy5p+Vo01kOi2EpTzkZd6tjbTzQ6r8Xrm+CIm/
rcrs5n1O4WPfPXcaM+gZfX+nHrsUErVWXuC6ZEoB2uPAHF97Ppfs6+CEERU318pV
h1iz1pH/Ebh0UOUArZaWshgN6Rhpz2NaiJqDSZyVyQxekAFDYpWAc+LS6dUswzxg
+tL97wantxPJs9azhkfQSU9xJd8qMwhL/V33h+UNA8r+9ggWPF/ubzrDmFUMkKa5
RsHQQ56JnPgIWIXNO7McI1csUD5sb82ao7AAi7k/j38hoH9nNK4v8uKMCa75Y/bS
k2fbOz3olcIe274kN247nX9p/VHemdiPiBg13q7B7UavpZSC+2bgMljOphG4lTB+
Ff0GhG3C7GlK3tsrsByZQJo8UxOTFT0sOyCz06Ya+D76TU8aOffI4FugZS0zvN7S
6mfo8n9o95y3abOkpcUa312y+PBT/ZiTyzwa1wp7vTWSEiqy0ebBhcnNkJyK2U+p
BEtu1nS5ncqZ6bkNA2utleFhXJwbBX6L7oqkIzfhg8WGv86fO1XMAfy5iNFWjbyv
yE+n3YyixtFTKJgkOOBxPNcYqx0E4K06D16dsxeQ3nv6qcgImIPFglmDvrPjf+je
4nWekfWCW33FonuaEpf0gJAELGXwwXTdeJZJ4jZkkBEzb+3zY5pGH3h01gnie38h
Dceb/Ctu28zZ++U0Ro/Gkv0OVtTV2DOvoyakjwmpxTFIklc/9a6UQnxMoKo0DghQ
vm5fiMH/MXf9Ox1qqap7aLGZgDMG/3CIXxk4s66NWn0PdioiBWo7iZLDLi9MVngx
YL/BZbZRI/RZxN0EQBogQAmpWkI/tFw8SEe791SKYg/NbWcWAj//7mKLvS5Vn7e9
6ChrCjWJRA3dcT25KtOWDdQuK70szPjG4DH9pokYap1mXRtARN+qiAmC7Z7Cj9Vo
r/5dWstLFsxCVGutVL8ML75+/o8bAe3SiS5G/REZg2ZNe2eBUXx7rEI//vri3fl3
xAo5EbsXR6+LPgYSHlTEJmkM/1PcU0o1n12vAHD5DdmcufgpmL1DgM8BK7WSP/yf
cac1/WVAVqkpbfpo9RHk05RILiWftwvI65UEfTyCcXHvkl9mceHYXmjaMTav6HBn
D3jwPEA8Ike5anYEhSf0M6ZTu4vNXUco25TAZcsSkW/QI00tPdwZw4WcH84J6+CE
Tp3zIDQMHHmPJm8EJV+2XnxAs8CcRUS1O7ug1A6Em0Nf3B3WUjsYLOa8h4dV8jtK
cxeKC+EKoRYBuBFuSZQ64FcaCB4YrEa+vwTQfvhbAgaexft0TQEA9BLwktgfr/dR
0RvJzFquF+xWCqBIWoIOwz1AacM4Xm6PcFWSFXR4psaahf6rJUiCUp90dDyQFMcZ
lTXUu4cKJZMe5uvHuU7HedENRiedkupGfgsrjgpn/Kd910hxOo00FhaWIBp9fjca
1NcBKkZTmlIg/xUwcUmRc0gir1csYP/DLkdIlBmTbsrp8uDxhnAZqnKkRa0G3gzR
4o3UcpCldDFnPaMOLwOlp+mi3jJ9XWJ2uVRffMjeYsOr/OH/RJ8kN+NT1WIcMorv
KzmBay2YbIQdvFuHUYYKJa1RPRMXC7QuP5or50BoFVv3hxIam648dVaxFArkhFBh
E97fOL1Fds53XVxkMr63Emvqj01OlNnRp1hKSTwIHAY1wRJ9lGe4kfAze8rNgbAM
t1gFWXojxtCygSDRpNtJPodQ+TYRTSfaBfIpcBBIUkeRHos/Ab9Dq6hNmif09hcV
TFiFWxWIjwXv/OU/GiKGMH2rq+x39bqRQk4f/4wr9e+/jdegELIVMuKm2xLrMJrm
/+XuJTqhK8/ZhgCchr/TxlGcuEoj33Rg+2Avalz0e+G4onFvN4Kb82a5jITuG+IB
GW8hfUh1LW/jBi76g4sxXEDUMP7+Ewy/+e/ySq0PISkUWMLmped0t5ZGEYhDJnXR
b7621YbwkgwpKRFOfL6WorTqL+/y4WzmPauC8/4vjlDNX2EisPvbFpXz3gWSlWc4
sPeVqXdX25B3n7UtD5mV0ZRhlHuH1CBE93XG0BGXhvCOr4R549Z3pp66e4+kPZGG
mHXrmCkkl2JDCaaAvAiVA2CtkwWnbD8tEQjsI3rQlHv4NLuUJ4wFLTB6ahvMXI61
YROwJKoEWdxCx1MowM5dFN4GLRIMD3XbBSm7LTY0hbtubYJCCZR65VbKcPNQ50mN
YkCH4yd0/98/W/DfAEmIzRwUl8FaoqN/OXPIdTv4Co3wuR0LHI8sFkIjlQ0E8jTC
2TmgdLgL/vajGI/sjYgLIxGOKwXAwvgAA08eSbY6QlgIJrsOqUS1ZXKGx6bHSY+g
ME8BfKYKgLdL7aNzJYv8oVa7eSjapEi9Gt3cyZ/1WErrVC/EpWItO6P7j09FzlQX
E9Fymkml/2jebfCvtERa4YXn7lrp1/Kaky11qC2nNFbqCqoZcTLRUbHpKG0SqXN5
qLwwpqmWZ7gkeVHQW7IssKMtTdpAFntVICsQ/x3zyJ/9zB7FS2CKiwIkLr738OG9
uSfkxMlrsplSssRq72/8t/kOK+Sm11A4552NUPJ1bckDfcedCo8FWYQS84CH9DCv
xIIgeO/qncAId4dHFUoSO1SpZzzJms9wjcPEt7yfJyaPqX2bp0B6+g8U1Afw9Riq
LpONZgEcaE7N4oXe8e0EGUh9zfzmB4/AGZtD2G14nk2JG1G+63LtWdIZDBiscMKp
D1uXMtlz1lFn0x/5Fe+RhjSWUr31SPQp2/CydvGNbypfm0OcmXrIwb6Gjy/rigmW
B3muamLxRbHBoaVoBQttwYuwbJJ1aBtjrj+DXuFCRC5gmqoEaKd6BXxX89+T1si1
cF5Nc9rIIs2POO9VrQNojtA2YMObxSU4wLKnbdVQwZx8l3112lx/aTbOnFTp/ya9
PXMwJvxeDBgVoAU92/zHlnpQX6in+NmESOarebFtG9EtRLbwvAFbcT/UZE0/48ix
JDpxmN6hYfQWahZwKmJU7RaDFvVwl7B/1LtSVBHa4dIVc2vTuQhwqbNb5CtLJhJ+
011o/9U8tCTD6ICaccZsU3qbgmkWKdJnwFDfsxuCccbaxehl9mhP6R0iT0FpkvwB
IuaY9YgSfmx+fNhqL64ARSKo/lMnsiR0dpnPSDqPJywENSbj/ESsfiSqhQQuzzUP
pwa3N2B+/7i7M4SnU3JWkxjObvRWzuYmfpttMKC5uFA0f/NS9Kn75ZsYyb4AOq5l
siZH44WogxxKvo7u9cuqrGJA5p1wpdEY/7OneVIpdsItJOzFUZ8sGC99gjbOxADY
F6elhx/PMTN8CrHNxlsnpN6VY3tRA/ikDQJijbflGqDRvA8tmAf+GHwkFZlAE62t
4JUQT0XdBxyWgd0dzbYkodzLLthM++EJuotmvAdmWZJuATRUynWwiFerWp72I4D6
ljCA7J2fkCe+MnIBRABe9QdfdJILkjEJmNffLFJ23/tBbdD+8XMnKhpK1W1/3wvp
Nm1gxWNfufCsmYMuFCzvYNTWZPejjXuD2C0l4PWJNwNyPvVoFO9EbvjfDDKM8mPb
dG/wkyX8uqGuChkaM1OjejO+n/PgbFInJ2p2chi516/Ev0A2XgG6KBWMB4kdW9+I
7FswwI5ZHYOZYQYRDsxTPghW0NCiUIEpI0tlO2Es+K9GrOEWNNWaDYYb4EvIvmRC
udNrWEoUVaRt3C7COfKDMbAKQzFWpAp1m+vAFzCXZj1TdPWV+QwZgwLsddrx/au+
nhldoSfg62XZVM/1ZdkEGtA2kO4QuUyDnVMJnFQaUBSkIXJ7et4eqQHRrx6/gfGl
jdX089OtjFa6H1C82jsLOXj9gWOMn+Etj+/kY/dtk4+6KoGswvHchhcpzBXPlbzS
029rh+VbAwOiAuDySq1jvm4tV9a+HsVK/Dw2djaSUeEwXnFz1GGSH9eehchneELx
t4nlkVFN2qPF7DhWBtrSsDjRuTjaRE1e3TYpj8LXtZkdpBUFI93L9rFkAWnVk+YD
RdaqOSK/FjFIGrRsvbIdfICyJIYu0AKeulPStbBxLGf2q04/okybfeBCcJJazmWe
vgxQ9pnSIBJMZWFAGKExkmAv1DmnMgKb/2RhWFC26YbKa82XhhNGEbtb8w7ZET3f
kDEaBKtOv0ZfHsvtCQZlG+XMJZzCkQHsHi/TCv5M09hAMA+3L+Gi7jpGaKx7awvO
FIhqpDNKl9Q6QHjfqmeT9HzM8M4QS03+gWKXn4r3AtWkiC3dwNCzQzQHt1CexF0/
VTqMgc7Y7Dch1zoloOIwJG4fPCcz9BjRwiYpY+zbewaRPwsN5l0VJ5+2rfG0T3Fg
hsLZO7h12QSuOwBzw1sj2LA3CYXHwPWcAS7g6wr+wjCKjLk6P70waPah1nkF9wve
bukQ+44+owO60yFSr4Y74U365PwKIfT+32qr/X3cwndGPoq0vrCcYyUbLendydJW
Fr3bl+upC1hgtTyHdK7E32xxK7VG07cLozXCAwGUIgARDzf6WMkMXzKVIZraSLpy
rCot4JTEmn9BQE4s3UhEUTzVkio4KsgaKdF16dpkb+V8HSgV2MyqSszz1TGm13Xi
LzO9H/i8Vm/GTLdRnEB551sldNK4yaJsSU5oUNaQ5n56BYGXXaP9T9MRHu7yrlGr
yQw90gqxO7L+EeYpF+HtzNikdBxm3mjrDwN8m50zY6oFaiRIcD2gLelXnzyyLazJ
yFK06g21zfZgdWE5l6w9KSMu+Bet7cr+4YWcFEkklSluICrtS+1uxKHlEWw25IcN
IQJ2G+ynxo5w6c+XPWSmZxrxTVIgE739krwIXHXApk316QXaQEy4yygOLu2ETiAZ
WOEpZThMC2JZqKet1uG9mXkoY69tNOgok1IcwZObCT/aU9+26EmOZVb4prhoDWAb
qrJE+cwrBrQkzCcdeVMzQsBB6M1MXNSL8B7kREFk7uVVZrkynjCo5J5pZM5XswCD
pnip3a3osXRd4DU3M9g55kD/lq+M1Z03gDt3Ot2m24k4REb8vrff0tzkiusLpr0k
nC8XHFOpvY5cRWCMHR9LAvWBEqOYKe17uHoRKvVrZ1qrJsrL0JsUoSPVoEjCr8r7
Y7138ExWB7bt8LSrZ8NF9UFEaru+u5PoYBB2eA/FWAUm2ZolGIr4VLSbNdbHJOPR
j6qsL5sj1OfonHcBEEe4BySLG21yTrMShs/B9ldVg3djksExJQP2uzxllTg3dXDy
WjtfSCFfNcMMGucVEnpTMLh1h5EyDxNCxdyD4+R0YQz8zDxPpUXx2h2EPzzH2Qbz
F2B6U6jxHnhTiaDmNg27wE6akTqaJPMNdwqu1fdVYV3Bt9LqGNVti+t0qjJpKT8H
rWPjizhqdeWphHEgqBh5HLHv+qyI8DT4KOoIn8U++43CBjUlZrxxznWUWp0XiANw
LuJfOYVte7n3lfN+1g0kTtuMjpHAqKIQs4KwAZq+wKNOyV2uqMDhu22xuFdWxcuB
SE/P6rtMxbekoSY/r7fQMp55/NLBcB830dX7Ohh4j7LYVeGH4kAKbNslqn0IhMCk
PVD9S2laFqeq+uRGGXGdZ/8tQ0bEx8pghryupWn/NyBDGSSGNq24NgXlUzF93Tqq
eCLXlFB9xmhbGG3TVt4Ye8o5FfCOIhd8ufvQ6NYa7FUIsqmVg3uoyIAiOLA+Nrxw
iv4ZgDUm7p6ee6FKQS2TbG3OOpZGw1MZqVyWg39spUKIYJleYHgLPZ3B5cDn1X8N
w0Rvf4w8WycHd3SgZw+aSE9650tCNNkxJYWg517at9As2w3pzc8G8vhxzlXoE/8e
Gawhh0mn8OXTJCGLiwTWD8NB2gx7uEeTKY9Ftg20p9Xea2ZdEqZsJc1HVLgSzT51
ouY9sZ+ZrZi2I1y7OHpxzGCqkfFupfQdxlU8sQqIltQE6xCxNrG8pJoFArMyyO4P
Dbh9nBx0TEmGp28sx0fkTVH6uW6DoglqtUX69Ti5XCiq0mR38hnMxvg1+WXzVMLx
UzZL5qR564jv9TrWK6zdf583TbX4IveHapD76pkHLysMz8RSv80sZ/6wmGbTsztg
RGxPuKMB/9PqwIal1FAP1XE7mEwV3ji/9T3MZ43tXICzbSFFUDsWH7+r4/laHL2l
gzhpjrd4TD7yuhE3PBOs9pogL0TjMIlPg3oIQgHUbELywgrxEWVFmj3SNLBrUXtK
yFf7fm9uemwBxRe7XFT2iaalu+8CFjIhvpIWRlrrd2gDOaS6gn05fMhbtY5tH/YS
0fOKmbvsLOY2pcXDCfMXvqkBsItubXWOFBmRK2qc+DhufLR7BE6L7gWOUMDHjx5c
dyVTzgTSFLRRMu5O3A/JcgkIwbpT/oTHxYa3lU1BxHH0WljuJZnYIqk6Si494YxI
qmM2L89IZUfZ+gTwJPo+HioMNL/C99iPlzTJDsPR6FHG+TQQbWXAyT9p81+VRTaG
Ykpax55Jl4I8yuBV4RKNej3/wwbyj7BtvPU7GnuN+Xem723fUkCj8FCzkW2hWj2+
v+2ndsR66oFPsBd67zFbwnWkEQPeYtK+F2Rhds3rduQtbS6wQqbQ1nGmANFNNS4y
OmI/EEfeDjbJx7puE0FtswzRZ60QdIU0X3My6o5YlaHpkG7nRjJZrCDqhjPwwSey
eXyu8uTefs+nz0i5MRvwSVmFr+KIVm/BrdOw78yKBvTsSFz40ZjQdjU0hQsqHsW3
srU5Xeu5cP9W9wFMn0tIgeaBx3hHqXFpC5T6x6mG5tJxmM+S6gvtPRHDzVzcblgg
M9sXBK8MnQanplf2u5Uwx8ovDwNdhAOPchfQR5fpsdTWl+tglJ8uOuF65KoJoUBo
UFwJkEtMd6+9zeOz25zch9ZouEMiFfblp0bjoMBl+lFZ3poxIbYOi5Egpmm0zQLr
+SMkC2vBKF8vAzK5n/yLmtS+K1TQ5q2bKnufLrvGWmuGdnu9IJK3QE4Lb6l95nmS
XTTmy8utxYFF7y7+wj5mPMAMY/7bcHPfzQ6v5oB5tDlC3b+90J0LlQZL+h4WQXvX
FMRwLQIU7VLOiRXk28tx/lB2c4ctA0qIj112RY/Kv1D6EewhMzorYvZbt/71mIkW
CcqLsY0FBXWyM8JTrckNcYJbEFVM+B7urt+KAnE8wSUNLQ4B4hlegjxRLzs61jkd
VgQ2g+f24kppbt2UNpnAdX/hi4QHYJLn2XifSkSf8paiJFhBfkXOuvWWxHktR1cK
oGlzWbFcWtldGrLCrcoBFamBt1/+utaHgZSN13djBmjrqraDglI26VXeiIbEMv16
z7WcoQHsppbwqdGs7ybYP/j62h65wsbGp2XhhP0FGjA0tEXMfaYr74LOP+xLk44l
ruuYgYp1GQnq30HLeeQT/iSLE/c9wGoLA+l+l/Mx+tCxynBAirxCRjB3H0SoJkd0
jozFAQN9tLms3qmVhEAoU19dmyN04xTyFBhlhW2n7wUuVJcEtz7uxkM6gOATLt6n
bwknYYF3damnK+EhXOHj5ca7gssLSU0Zk5w/GWUv/jKKBTDBmVLLTVOyHha8zwDX
I6fu6NcGFdRKnf9YuOqsqKUoQoLq6THotFyBKu27VowhPTiJkPteH7dvIzd9WAB1
Mp+BaE5zyvgz1N7Ag3FGC0QuGW3t5AjbxnLvlYvcEsizfr47s2mxGQlr71x4MV5E
7LJ2k4KUqoNDJYb8dX8uAeFs84mp0yJv5idjmcU4LYY7jYyyH/KiIHVsSTiqm4SC
e90ZHl1Ia31R7Yx1y6EMVngtAd9t9NPIOlc0uTF5DoMcQ7azyWbYBYA1nKsNcfdE
8RCPuEHVBVAsx9hESb7MqLfF8fL19HIx60L5eajGWtz5qFX/uzoJvnjAL2SXEg09
m5Hwp7/wJ5mszP7yM4JsHit3HDjIaXuqUujWUYIJIftCGq1et7Q8CCRr/j84FvLc
QbvmsgtZd+sbTESfRumRX666FbsPNYe0lwHC92l8eE1N8vX58DdCUjNgGuBtB/UJ
3KiqbmxsJhQaxxxKQ0rLNkwwd1pWemp3NoEZXypLZGvKuUteUztNUZEntC58I0R0
AinibMzMgjS6iUYYoij4qBKlv3VMYJEpCwdLiq/aYesfxXLkSa18F3tU2tUtvb2b
tn7CeBbwKf9SFLzf+dxrrVUh0FG8h7CC1VAMK74bsojvdE7PTYv7s2eDVo+fV7oD
4CJ8bQAcC1omE3395NILUkzin2XnPWAI/FZzkF146S9p4N08+yOLpc1CNxIqielo
WaJt4CsA9uZ5ZiyAhLISDy8JznousyJ2F2vVoBGF5mzzr6cXKxuEBL0rJ6nA0t1X
+Sg6Zd53nddSwnXSUbC/5+kmA+VsUfbkmTALn7232KqbHHsuRjKF1ECTJCLge5gi
1jx14PMqlWiLfEWz1kRUUnTUIHLbnZxyGyespmca8Y6yai8oiPUzWobHt4W/f4rI
BofpwD6GitLcGOcLuGROtDDtXCM+/STD766c3MtXq08aFBw/V2sqfqwQSQyKk+Su
ckk/dgcIVhH1nrrMzypFFbiKg6u+Vyi99G41on+gLD/+0At7Uz0a5ZMkbV79kFyf
aMPLhyTE8JeGdMCeASTLcNTM0WaJbdGFtT3mgqnxGH9vYIlu0hL2I8U6Pt8/j7Ui
h+y9AN10Uj/34YWfIolzNJPlcxy+ui2C20VjVQLCXarpHedQwJPdDqNif4p84P3C
XJUJW3TpmZm8tQCScVIMjryvPzcxto/35dJRdlzhaSviDYacdokcUWfaYiTM9xrm
ZONd8qnxev2eBxThjxvuhJ/NLpM408aGp3lE/mNuVEKgZTgYAx49IVunuCDwlCHD
o6mcc3H1SQ8kkp1tKVwcas2jkGMv998ff75AXAxuiv8jW/NI80bp/DlQnbXFVd+h
SbLS+czpMSRtwmari027cXRyeg94mZLwx99pJWpi3pz73WwE2rnT0DFZ4umyz422
l3eXP7QiOBJIDzMXF45CNfYmvyGpANhwd/BMm04pjR/Y10eNaQPXmH0vAIq6zh9F
m7RzmV2ZcHkcEFk/Oulo04TJDWQqXnyC+Rn4IdKm2bK32yuZ+wThlqjIea8Iq+pw
hHR+DFfG2WQ0RIvuyHxcv0GVUN+CEd2jxyX+tlbbdH/CrqxkTwbo12cDeoOW8Yzf
53w3S1tpocUgm4PUqHZv+kEq813Bpm1sQVqaJu87IJSytc0UvPi43nxPFRncvtGw
R5hxFnlLMOvxBWkLEWFbltujjpUIJwCgr39WiM9qWrc3dd0nGqLB2lSf1QiQ8KFq
uyznjo90/oL+buT2OpY7gzm916Kqt1DnyR888mSISGmuGc5x87SIwDzLuEGFpy7S
pjKJjYCue9vF5y/cEzmX5joYt15lILlrJ8PtSDmQNoWr3+Loiz9qNM0bLdI/zqYR
7R0TkEEbSlbC/wSkQ1kSKXBxkRo2W+mPZAIOQE395k+YHVD3EIncLNE0FAI9iyNZ
JyFcMEpKyAqBBR9I9JZ8Rmq8g7XFPRkdfSD7Y1jISSwwfYj4gWkupfWKUtJ8I/6C
Snom6mtLCmuieRc7PDeWhgjsTMKQs2x1hMRTnbNsorTv7AkcQ5L+I/QDg6+tqlW3
6LcUwviBFq+NhS1Ltj4KoEN1oYFH6nF828N62PpOwQlGb3CFcxPAwKpGnQ/dXcpI
UkHOkro+7AgUfFDkvWMux81E0Bb5ELADAB3OgnUoZotJLCZD5skkdvvWjzKesRtr
Og0TtLUItOS1BcMH6kiAMHCTP9LI/9OOIDN4zRNea5a3vohxS15Sp01H0Yg4n2n6
OTIS9xG25NNJH87Y/cdS0828VKEpNamkWpdIZ2w2q9j+m9zkZNAyx+cOdLQjnt+j
5g5vzcq4P70DwVO+54gh5wasgzd2kPqkQwqtOOAHAPrWcjuj81W8W5YY36znFrLK
86flPnGdmyuIwBYf7aCi/Q3EMaAStdmqvOc7dONSkP62VykKhNu937t4/hE/IVfv
iBFaT//gdCbgyf7RajJD/vbWJIUlocelhmbH4Z8sRU1tUrooyTTBcjewOOR7U5Hd
F71h3O868jjvif7s26KRnUsMmEobA+FV2IFo8Od4WUIS5ScX5RATmBjjxZG9/Kl7
XA/aSU50G3DehwnIeFtL5vOE8R6vFPin5oT/h78/BTzmvTGexqnrRcnOL0JHdlz9
MfJDOXNG5GZWxbr9AUmMLmNoMecBgsQL5BW9t/TvQg16xOSiXrA+0jw6dCQwesm9
T4qWw/vOiIVolfAgaNFBPLymd3dBgFFyLRC3s8/3VHSCNgRVm5OUDDnir3kXE8nB
4ajET12cW0Y9Oade4Gc8qin4MLxmjYpLJFKgH2IPwB4juaA/FJkq04HAXWMcIl/f
9CGOe9czBTUBmZOLhb2Gf4n9X94Byi286Sr0XOQ4AtMgYNcc+K9g09YTrRpKWHxy
ajFIs4xSWNgNiMSgTVtkCBCDtfgiNFi5N8VynWEOofkIoNe0x7wE5opuR26SpRj6
xnmsq10mnTC4yZj+22Brs2kpUKuNabtB1AReC3wJezq9EuDlMLHRMIIa7opKzD+X
ZUfyk1dtuPpSka1F1jzPMQopgre8+9YpcXuvYHLit8L58E91hqbpDBJTZTiLsMeE
IxaHbq4FlVM2mzCW6x6fDcJ1nnXDnmq+jLmjEHq1J8PhCgoB1xAPMueBj9FPrn+t
u0EiXVLSGhUdwpgalAk34JgHYDpYhVoFwq7ELgD16i/JbfNI6IKpO8aIQNFbvj63
SJM+hvwwiLkGWfh+oPcPe3LTJlheqGY7lAJ67K2eLHXNlkJwe3uK47qPeFWBwVpU
l8acPZHlPo00LKtjPR+b7nioZomPYtJpSZ8fJABu1Fa3kABwVh6eeMDlJAfYV3Az
XHvqWctUcSOnR7Ox07hk15tNr6Rz3g/So+p7ghXoknw2LU2kD3e2jtAfv+spsGTY
S+M38S/v+ALEL2t/JXMdodJKYZADMnrc8X9tPkMJWnODdTc7EKl855F7nDF4YwgP
DmCQKiqir7HSBjEc9I9BPA++QCU7GF1ky8aU+cyoaXResM8wvUKX3h5uNG/fKLdX
xTT29KDD7BVGBrGK2KKDNA6wVeMQLt8HlT1ANOH2Jzl+pXnWMlkGB07uWBa7JbiI
qh8L+fsp7BCa1GuEY/mj6LGl7HBzqCqgwBPKciKMt07yFoHFTBi84UEqNOovzIEL
JjTjFuBeBzkqwYUZ1XeVHXtoT/35bR7Nyp4Io01L681DcQ4G+YLwaiPCNwGQy824
GATitGRzH2jHhxy0YJweBxzlqbHsRaT1ioNKiW/WN/YjvFEhlNcrtz/9ch7G0psr
aePOfKzk4Bq0eQIrELLxqboFt0s+6qFuk/wtS3RPJukuvPZzPvj+dGGRyybqcpjL
TXHl/BEXaI5albMdnk7q2U+cYEVzwPc3bGD7g2abypFGm4fra8yUjVNk/KCoVUgg
MLvY1C8ZDnODwE0RKD+T8BjgTj7aa8KvWngmw3h+8PN05nyvdAUElsiTrzXUcpBH
N4aAwXLzTKWIAncXJxRsroqD02NS/snT9UtMFVflsD5HObkS3NK0lnvebOadkhM8
UvYWb2qxbHtOQeh8uDDNi34Z4z0hZvUCnO6GCuIMkQ4FOa0l2ij623tb8rjiKhLF
GNNHyqZrqlRk41+MGcxVCozePjEptjlDCagU3bZHlSx6tWTNQGjLj4m6tsr8bvrB
E5gd+jrRIOx/IC6KCDGmj8d03pjY3VLivMRCBg3LlranoKc8NNTlvlxba14p7FFx
G0p1pOuPAcPCf/pa9JTLAV86wZepPq1aZL6zXXAPNkh9N8iSFISC+KdPqwzxemhG
Z+0AEMPGENAb1/JejPULpwF/2j01T7v4nJALdyWhZv0Kn1IxMsYJ1OSf5nnj039H
o2EogVKQniIu5SzsGd3gsbrPg78coBbXGhx9JuDP8UUPaS9I0pee+BMGpxVeYzn3
N/NkOW5gng1BN+H2QC5IzdkfYgam8GAgek6xy+1+aOhnOuzpKFhstQjYq0W/pWnx
1aFYIuco94dpg8iutvvWJSA0lYfu4esvBxSdDQXxe5jYcOSXZk6+daKYnHlY5RxR
DGGOMFK05+TqwF8ennZMGSgSgZ40oG6uWjGZ5gkRD5iOWtsTeYyL1x7pq8CFYnaj
afv8gDP34k1ZGdsnaC3lQNI1k/Ql1iq/IDf1M/xFRutGai3GtEcY8d28lINpI1GB
9o7vPe3bxEuVY18a8fLIVIo0YXlm5CDrQvtk5k/Qu4lOZtORad4At/bf9yVIbvmZ
ZQbrA5i/szbHwVXMd+aDHcrGGmuC4nU6O4D1VFFcPOu9v8r9PTanzK5+0VEcRoIy
kv9gLA/jYWuIr9lqgGJ8314vr9yrR5MtZ6aHc7T6ueiSxJuE8LoTaKpYEkhwHevB
WtKh2zoypSsaBo1M40NyNkN0Gt9Kpvdn19jQy0Kl91JoAwShgN7GztmSmwzcASWY
JAiFL97WRzJ8B+NIlln1oTuQXQamdYB4jD0b3s7uH7D18Zi0BBQZ++2KwCxHLXaT
aMheOmY/Q3ClzfrwB0jZIjK/yK+mDsRNulWMNhfqDqyuTaSwlazUGLOIQTXiV8g2
97eZsOBq9OOAaFa1ak8SG9QSNtKpyIR8Mit+brlq5BlNwmCG3MSU4jc92sDH/GoU
d2W9CYivTrhHvahkSI57H6go2NnPPC+WQ+XLRAKXw3ztCUYjjEpXh9yxhtXtfwB8
gqwvs55uVSUS4dKM/CzdYeYGjXvr/BvD7DlHcTxUM07I9AtznePR/ABC51L9zYvv
O1H/7FQf6T9Xpx6d+xSVzB/SjMJqduwtQmOJigbHC2b0gugR/ZSJp6cBuWU80Pel
RQgi5yQMioU2TnvLsFKBRJ5VE2/MZPNRbeRZ8UTg4Z85fjNrwcjRbhonylXPmgz9
Kl6KZWWVubK8m4KYITGRbxAHPGa3l0FJLOCEdSAtPBjd5gxdE+O8RVrewVfVjkUM
ShhYhaMt2s2R7dnkU4WyPAvCmUwDb8+/w1u9wsFH7W6rRKIz7bA64aGvRkh3QVCe
z0K5AilzhX6rF57jT8tBvltcaJUhqkUoRaieqOIwDf+DV/LP2RZzCKu+emXwbCMx
os2CjvnwrBFo0+VVqpTjGA+mS1zGAgcna+5UwQCsUFlxV7A6MuT7Fnqa7urRno4F
cyhceQJrkpwAXpW/c2EEaW2CIMyZQNfhmuujFfI7NUMnDpho0/JWsnhn00N4xDTJ
lpduMsDQCH9vUR653frPqU8buNVh65gc5d1h3OGciwRCWav50vGROqVczOZhUdE4
7e7htV6FQlTF7m+GfMEz/8VdoNJ/6FK4j3/dA+AkMluj58XO+EoT+ga3H7YTyenx
BVJ75R594vZ1Z8kAKPvUMa/8piExDEsEQTePZldU+SZShmueAr6ZZlToI1NkR+f1
LnzwImxi8msfARH0AXY7YCzXchKB6ccojWvZehNGU3qesvrvsyGlVziA8uO46CHk
ljGevUBOGeFgSctHFGs6rgOFBHR9A8KczdJrq/d1dTE/wWEnVXEI/WMr+nwJudwJ
EmfEYcYYPzWYfBOrK7lRvvSXaYvC2TOHMIaikmaTLmPVqz+HfrP12MjK2K/bhtTR
A1fBPysx/lMIzlAofx88vL74dyz6S5QgiK+no0VKlWJ8QrmA0JV9VW8nfHaZuFE4
EH56v8VzkdjWu1GCOJ2BepJfzxQnx4yd8cib5FXeyhIx5syUJdUkaYgkWkasnTTd
jVPxm6Xda8WEbJ/x/2V0lulWN87udR+o2bDjg831ajBqoSq/WWWlNvTINDMJTmvO
UMPOu+ALuT/64iQmU4t+sAmzqxgEK/ieMlV0eVcufRD8bBtAavXeldChMQvQPMaV
/+8vRWEq4/Ze1LLCrt29DNTGenazU+fw5GKnZqUyA6zJFVxcMYfCYHqJhD6SAtrh
fOG17K7LjkA3z7SJu4Be4Lpzm1hphsjC7MrEE170BZv34I5GqTDDUBgitk+mildl
lovt5GUdF8YYjLleMQmMDYUkmc2kEjhHZfN+FH9qkInC2Bx98J89nvWsXKutqWfY
/ex4963u35yWLGUoLla8od+Bve7vQGNPU/98IVUqc+0=
`pragma protect end_protected
