// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:46 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k/2I8knnXrHSLcPKUp6dsS02GjmsJVkMTOit58yujXAEbuGAQNtwJSI6FOjfOKY+
V3RkYeI46Wxzjfcgm5Ycxll/Npu6tm+y4HyIOqYI1w3HPA+wTBJP8DBeCBdBt+rS
F6aTL9PQArdyGQXfz43kn4T8R13dKfRxHjqIENW6qCs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8416)
6Iq4VsAtnvmh5qJYhMbIXfrgMhuqqKVZq4rYUjL++mI5rF4nqYd6gV5RdGD35rTu
2LmSb675mDPNhF7dqEpwfCa2Emhowyya/f4Ex6wczRO82tHBFpNVuMNRGQOH3yNZ
rFtLxmECOkw3cXqeqRlQwOdJ/vSkNc6rWav+yyReq179a/+y7LTteHeQbAJ71WUT
sT4wiinFBt40alkR50ERoxM/HhgfHJSqjfJoOCFEeJgjq6Dlymc6mKn1E1fynGLi
9DKFgXBiVMTPmvsbArQHA7XqrGWUuG2TGhuq4gF5eGv7MZygRrc5QjsJpkbPJtgO
oOsPS73U2/WCQR2V6xKzNr0Ymfus8+oxv7BKpRx2r0d7CDuef+7KN4LdBWFsvLSf
s/bhHkJWm2FFzVbkU6pLx8N5mrX1P/YotoPhfRUTtIj1yLIOqGfFdKbSnj4u1XZZ
6Po3OLVk+cn0DsU9xetv1+RfbnL5wEaSFWleUVG99WJYmfWixPX1JYsNuLUjIGNb
MkyqkZyxsuRu7qx9CbGhXG50zbUIDH6DNbxyVQIRzjZaQLi+zoqUdQiuIT89zIpS
3MkRH2Gz3Ijm+UdfriCOZNZUTyjbmEPWDoR9iMaUmD+t6f9HRVfyEiONwzpO8754
AvgEvSdKpm8Tx9Z1/nBVDo2kPIqm/LmTeFs5yxN8KBNBJWTZPFkvxpig+7Pf5fMy
IoqVpjSwjNYCRiyc2RZITU2NfhVIa/2HML5/5is6lNw/1/yfNbnn25e+/Mv01mWo
IQ+i70CS4WA46aT2vOkTnLLdZOe/07zbRIjrtzZfhXnhA+qXPCfjHJmaeucLl5VW
lJFhqeiREnFvInYoI5y6O+5hwe4Knzqck+wLbkB3LkDL7Sswg5h8DCNqWUA1RIdR
7xkWHAdVtTos2iQE7OuAsXfhAXv/r20sX4Di8Hu3+lMZVMNzm4jM3p1pyakwHm2w
KEkZTS5LFZ7+F4kMVZQq4J+rmrT36K+6xz9THtkDI2b48/jw8hTP7uPuH1CBJJWk
ePzY0qyKiDThsS0XQDrwgTcWCPzpK0meb4c34NuCQhysfFqraJjdBQdYtvdZ5GT7
MznqcR/NmOFPcuBokE9HbUk68ahpojUPOAyoH+qUVzJ9lk5AxXQeTyf542knNvFe
hQ5gzwODlyqSbM+z+d5oYV1EbqnSsIPOg2CNbwApwA6+IvERU2AnzYGcUZR93J/i
A0DQpZPVuLxEsgUzQFWrH/maGdQN654KkoBl1HZRzQrYbBuWoKiSMxXCeOa4CPAk
PEOmP08SYVBBnCRwfzFXzYr91eVRVWJGYiJRAonfD6o+sD4StrCHXsNvW1W13fZD
iYe7kXMmotS9PCDCSvdUtTOcNngtoVJlZrvMQ3J8H2TfWYq46Efwz1GwBKe0uHG4
4hh4zceB7Wo+IBZ1EwwtOnir8LV3e7GVGOsT97Xh3L95SHfR7FNAXCOGMX0JMFLf
BuRYOOsiAwmnuvYl+AmDPGh2XDCSYdflJKxeW+kcLLKieUidsayoEaz5VQoWq8Q6
OR4vSepsR2sunchFAT2//DOvUHwVsPKSl7k5/tAUBipgeYtvRIclejWcZrUs1ziz
5+RsVhfoKndRRnXjaUCsmHLvdCRbQLE9hsqn5blzxvYI591IQMOChM9eiguqwVFC
UN+NVOFkIrKhayo4I+na+w5hFeFkuQ4P5z4UB2FBJdVZ9ks6DXj20xv/DvmmD2WJ
QJNr21cCBSn4Qw4kwEr7IS1hVuO5wIViD5ZyynUf8J1OBDOj1x+fBQnyeTLaU9xO
hcWK3LYIhahhfMZBX09FaPKjYc+ZxjZD4BVG5o2szY7qnWr8/WDnNiJ65wBwScUQ
uw/umcNoUp8/TdTpKhnPQhmyKPPRD3taSCbDJWe9V+XUzS76qKaRHJj621dg2x6U
wJOZmbMgWpjBknXHZQnvsOQRM74peEo8Yo1s5h7AID6x4cLl9egB+KeKYw1x8Wh6
qNqoFeurCgI1Zca2skdn+BlNpW/5cUcpq/e4UJiwgg2TFLdSZjFfhM9mPZD2UBLP
tKdjNDXfcg4nWknfIUAm494ph7n5RkucSHVAZ95xDal580KOjrfn0IuYt13cn2CS
XzL0iy2aWpDCllYnJ8PGpO3dTnxFLSpGCXvjHV+/+JMSPCbcrxumxCZZkwcnnhnG
b4S4r/wQwe8fCN1kOt8hxC0sLE11GixIcB71FiZ94XZ3YF5KvWyrB46IeIExuriE
HKdolCepHzRRTfjWgJQSwMoQUEWlorovtzxzsc0OYe0uRHuPc9pc0DFVOR708rbL
5rHqxRmJyFNXtkF5pBUPVTSI8GYV9pts4Fo2GQAMpwkw6zk1oCOZhKfTv2nkuSEW
Nc4daGnWcVAWx5M3EqKVYDLLIfJqf5wfAI8hpJo4VKUhoIh9bbBs4pQZ4swkh5Ek
jFbZzmk1Ae6XwRTKBwWg/oevSa4K28GsnKV/JfrcpAERXJc0McJZHMv3T7nWN2v9
ohAGyAfh+72r6N4Z1O/h1SYXMnEV80viQwL94F8FRhDhuOtA4L6q0fORVSN8Fika
tdX/xmXOf5yCYxnAhUm//I/vJERjjEb32LcZB8Nf9RR6PrGiilQA4UtBfll3/WMi
AAYDRmA+951CDtOtQXOMcYM5xeLi8gC9gjdSjbNh8jhDUeKZQrHSnDnxFSjTOzE0
MciA4w8OeIMdFGrkvcDlM0hSKi6kM0KMCpKiDmtCBoiWpNWTzc6fix/7egSqNs9r
1rAajm1AOBnmxBLqF3dwKKTMtPHDWRXUxWcjs0Hewz3gSMrgeBe8cpjrWlrn+eZW
6A62mfjqq1B6MB3Pel4j1mzCfjEBoRGC89/tM1B7449hOd+Hd91B53q8nZ9IXHgg
ijUmm0OmDL38XZkDVEKVqY5u2f0AALwGViQ667xEU45XGHqGlBordu5JZaKN4aG8
OpPwAm48KjJMUIq16t8mH9KisyhQHSK7kJTMkm6rYBs3DlnzaNn75J1rNg2kAZ6J
iIJw8vqy0hiYEThAa/R5x6icLj2zUzEAPpjAY6NUKPAxcP0Bau+bogtqXiXlhT5X
xIaXGrfSuCdU7l3pdZ1SRXn36KRDPiqD7PVyLMzPZDboTf/h/EKn+0RNEPpVWQL7
xad1zqgBAXNDeESfa9wV/SqB59AKwQMs/ghIaMUcdOTqnTFsLvVxxUpJmzyyVxCt
kedjXnjfZvq7h6ezxVpnwGUKWSxedFvwYqxNgEJjxj/YB5Nv3NbhU36bdH/R5d3V
o+0Mbp1bh/Lz3RDjFtQIipQqrybwPFKY40RDgg55VnjH970XJthpf6BYb5o1VgPT
WvwfyJXA+JxtmD7t6PG/2SoJ3ITmF9/DmTbItqAe98l/wKTdRNIK8ytRPrNzkhZw
WAsdBDrSCThbd+1Bnz8yhdsR3yYwLRBUkTlz69P0E+0zEaFhMXqhISb7zEjnO8ZA
94yFxAOZfzcAlBF2al8W1EZVOFJ/4fXGcBy8ck6tOQf9YjEU8TVgrCJkXahY3IM4
Nyf6OffebtaaPgmPxXUMbmuJyjsqvOKeEJ7JIQI3AWi7rR2HxwAoD+9h76Es379r
HN5PoONXDr7t47Zv1dPuwksHJRogOGKuzAt5vNJSwR91mcqOKOpSGVYfWkAYgOVd
RbvN+ZvdqamgjRMStQheFHkpztu581/VBCC8J8Z012i9MNXi29E1ork0k0MjXtOj
HCST6Qx7winwUPHxLrgkJ6X5PLdJAWkh6uWd+MiNwg0dtdCq5LGbHAhN3e1xjzH0
F/uQ53+/U7/9HOL438H4DyR/wwgdW3NBm/DnFD4yEgUR0uZqsgQUhMCmcPuqTl0i
CeOyA6oZrsmGhsHsZJtUIeHvaBmc7DWd8kFf+eKDT2kPXVB+ybu7S/B3RTkU0hab
jqx7tJK/tBeaGfCocaxBXfPneRbPXvZs9yXNUcbj4FFVkos5Xz/JtpCjuaBkll1T
4CmZoBDn8ake4YwKbv2hHcNDbvgJiSRc4QJEmKj5iNLw/zqXhEeFqJOrCLOo+s23
bsYxm2nrhzVcjs3ZS/d1X1TwPwdvQLbqOwsl7jnSxh8uaegDl0+PQs9WG6qIsMBf
Se7sNDqzw4Wywp3qCuq0d4s5L8tJeuCvyFRkcbcL4x9gM5OsspZZOr/ZGOBW0FuW
yIDz7TQSriff6oYtoXvq9vy2SgQqozPvGPvhivWF4EbNTx1UumSaXUb9OEfNqnmG
B+hhP57Ft8YsCxL3j3hvNyFFxu4ED4M2zxHEV0uv6QEiVaQNH42gXJ3sfrKNkjMD
ILHTWLJ8TYCOsMR+B+sJbnlvi076auwqdTqAy0iJ3cuodGj3bn+IgdDLU6l8UoeA
UNaoL926TLavphZ3Z/73+IIo7AHD6GfUoqFJLWLl3pjqyhKPR9RGHlLfnTrtCHr8
1eg7gZWgb1dFlUiUr/GPQWmAWBltqa4rYSAlHPGXSsj6u0RyjsSJiUXZIzHCo8od
yMBOQS0jjcjPtoejz5/NXw7jE2xs/ze13IFSD3OaGbXnWRVyHJuAZnwNs24iUPpY
y/gp3JygLU/dOTv8gNOHdBD8uqUOZNtJTCfe6Edq3AZu/y6Y3ZsHlv+iH46i/o00
fEa8FqxL6ks2FNwLVokMbtSSlAvol9MByDrdR4BvbLy/h2pSLP/ZfJPGOjKXcLDG
7j9la+SCiWl8olBXsTNeqXcCMBa+O4ymiagB27v3j1J/Q5vAbGfDYhy9iebOsDIs
Gs59fFAXhwJb9CdPQcJdPYGmu5d0CVbYTHaZC7nlGrBuZePs5eBPCal87PFQ+IBs
1EZuxpAhizvC2b94v/lueITgCtefa5Wd1MgE8H0RFl/A62pF8XYw7Yp/oP45oCby
xZSQ4R1gy5yyqM6uUZHTi7dJlmBWG3eEnnCXBLSQ/VYrQ1Y4WhamQ0p6xrLP9cQh
vDdHSyAbE9IPHnrPsg8uGBhiu8MQVzB6KW1jlTD7jJgyo8ZpLwkJj1qu/UyDT93X
YEZ614afeJDYDsFDmm/Q+SHbyKmayjPHdU7HR/sNkqyre1tn2Q+EKpLG6HgAvOxy
yxeJXZfLeSTYzkHCK5/tNv2JFROBBXeWiM77Scz1aOc5K006RifbHR6FiYpWwoiB
Wrxr0UDBRJ0qa3LaCVU2wcIQP/4xTJo60NfzHgEs0A3VRzhwNMujBo1jqGP6j03K
Rv1cFKOYc+jZsAccvmkWwIFqKGck0vTGx0cdQ63ZubDZi1timUL3MyfRiEI/ITvq
b2es+f9OhZznuljJqPWBYVA9p5pfQMNZV2xaxqFSbinJiKVd4KAxmOT0TPH68PSO
ckY5qS5VpTrwLl0Z5uzeXtjVehtQBj/RbESGeS5kOaABcp95UkWF8/SptlyqcfP6
CsqVnRJsCfyqGh3KC+N0ttlOPPDY05hQSDIpVZkVkMSCHo+1IastEFIHUrfr/Tay
5e3QSFmCoB6Rje/WEhJGRb/bSTZnAtAnkWNbHcs95/RmchD8yKhvSiDbBng0oQX9
huYhCcuUTus9dCJWcc0rW7uT8/tqWlS45kVIIn5OelOr9k147e/3XgquNPjDnauQ
HdA+cuebbh4ru25eG9PBKwAGcWFV33CmS0wCG0Ys3PmSkl6iu4vOB7A6x3ZyteZT
QdUGZ45W4Exe+LJXXpBshJmpbPqAVOZKcTFxmfPYoe7YjQKh8I2TxOAks46hLl+b
yytQG8vqymNXAzIP9nroMHKw/Ow2WDsU8tVsKfUA6G/SiitXE3nH2TyPuxDBIptF
GDjvHXzHgTA5QDNRi2P1DFGwCDKjEuGY6uejzEIHKbADnwrSoIlut8/GhTHkCgHw
TF8eFVDErbkM0CVVDURi1Ah5LX1d2G+PgzNjIWEnYlVzzA19HhpNSEnlM4LtJnNQ
cJLkw+FYdgHqIKC5OW2RBIO9jawm+1W8XXFYCiGQDHHzwFGFB1ILwoaF7eO7yFsO
cQVf6hcFqQZdNIGwF0rwpBD4E36sXUFNwgSmMvEoS48nyg/GCOCnhtmQ4DVRrxIk
zAc6H1Tx2XZaetVbcuCXMiyTSr5VuevOpuygoYYspWF3sN0RNo40d2zKsqaq6CIO
ntOCjIpqV8nrUSJ7ZLhLCZJPOapdWa8rjorYzjaPsi8otIU2PPZeu3n8GT2pc6cz
5H0tnjYS2z96p5/nIP4Pp5hW/6CzOm9gLqcStztoWh+9/7F7HXepN+NLQ2ZnLIrF
4Hb5/q6yQ4aRepTOJqn3fBZ/TLkIW5LLNif4EOUxPFprWAfct0DM5dWxirvXM6O+
9iPDFul9gVmOrhCsYrwZ5zNMNC3aO8b+EuwYiy+qTkNG4DorVXVwL3fZxy2D9hNY
LUdX+UowtdsuSLpyCEbwY95vNKMu2McgQMf4yeb6wP9MXKNDZNUmBWDINQHm2ZOP
HC1sPRHpQYSe+1WuJ6E/cilvFjRlbcea3of6QJg650eFVzCy22Av0R9FM+GZLR1q
N72QF1mn/tR3P1yez5vfB5TSPR8ClFj6KH5cfeHI1p+x7WZ0yG2UhhHaARnfvIPW
vty83PbLiwntKH7R1MRF5px0ISzZfTgeZN2IRiTZ4z1N+zapsF/SA5rSv4QaF0HZ
qFL0N4K7ZRRkEwir6EBaobELgE5nuP0QfuvPm9n2ue9mKc48WpmDtzJtFb6xiUqO
Kmb5v81DM9Jcq24imuGVqEVTQbCTSyVwTsC3DA3PhcCPwYCtki3mTlO8GT3SMaKk
D1lgCFZozrYfeW8GRFOX/EQlyYJY3dNp/R7fzsysl3YS7cJmKhBvBYJ92Eg1y0uB
JPBL31AYADACV02oznWaAknmVkC6AAv5+oxkIBS0L6AWJy/QC/XCr5FK0bP+7xM2
KUZHd5aC0g8vCBnvLOUhUc22bFw+ABqw1ht4/JCRm8MQRMqMNC2F4SyleDKgmKmL
P0qwHBLNX4fygkWzT+KuepPr3OEN5nCDt7AkVMuf7XJLqvq9OYLfONoMaQqNvP6a
UVs1hNc9tHEXQ6Pps9ZH6jv53fd1drFEG9tDsw2wjByY5lhGkwxHjqCZtdnvBFi4
YRcCM4IMfb37gMF8uSSyZ25E3bHzhhoNLcBU8XBGjvyi6t+TipIbVSqD9Rao6Xav
msUyg4PnmEYOm77buR8xCiqdSJNC4Y0eyOKDWjOE/aQSbvPGFsEw0SXGZDxaE5oV
DomHSA4f6vurQ6/YIXIh4J5y04zebMpbjrgRFYUQZb8MgKgU7E37bllK+Tv1hmnj
eD/sEAdNq5WY1erPR0IzmPTfj/Zws0LHLANgSJkYaKQF4jthBg8kx9xO+XyKtpmi
gTwBtFsO4lV/y/praca4TehXZJ5GgBfcHKvKW37Fb3ega8I9UeW+efO93cD7TMMe
JdacjG92cCgAEie65KsHJUWWvP2Y2CtBB2fQcuJSqpiaIRuLlgrCI5P4l89GpAjc
F6NqaGLt+rkBKEyhyfqAO7RdMrOmtfy7u4N/5stoMjGe9tRxISxfRKhZ5StzMoNY
6yONaRSnmkECWdcnU1+LdqyqFnqqLGA9rrOBR0M4lpZa+Aqk4H2+I+crvqhhru7w
bm7g3BN0B5hbgLzwxaKDspZP+C9YtnFVTianoz7MnsCHnFn2j6zk5akZst2ulqTB
61oN0CBcClYSCJSAdARXP2VXr5abdgNwih8CZQjdAg+YY9D/xH5e5OFft4puL9Gr
rM1Stx5BU94lSvpw3OM9YKDJ63FSJanJB5jEPhK6iY7+IiAXlC5JPyWJcoUmusNF
ExPe+gc/7Rr4D4QKALwoT984lvR+NJgkQL5lZtw0n4LMoa43bJVOg38a9Lj/TgD9
+9HmwBgusAAGZt3CbcCNnZxylpY+EabMzdehVAtFR5TKbfMoGm3DnCcrFVDzEZKr
sDay30xqlluMWWPo6bPYlKhSKw3SqsL9Q46C7s9PzGi1vDVDh3Eog1Gh0Oe2rnKX
hTsJNTUBtus4OFnEk8B2Qwlg3Djxcf4fA7BrZE0/qckIskVQEbysd0xNZCs2P0Sa
6WbWICv2mC729Ee2XXFKY2kIojpZZ3JPGmLpG5H2lbmx5SN85qa3s3RBJTl8BWcZ
ippBWrsR3uxBVxj1Cuw8OO2c5UkEPiEJUBTp+FPkbM3oSkQ/Tfr9pksHuiQQtGUK
3wS0HrNuV4hktU8VXZmJo6DTwZCi/pHx1xCiR54sVBvIRbcYZwRqo0KtOVig17Bk
qiuX/pvfFCXv1stxsKZtKNDTrIDU6hKrGtOB0dqaTzPB14o7fxKuB/lJ4h7rE9Rl
mOMLk6b6u02R+Oc8IyUAjrQREpL609f2R1mddz+aIOAD0ssOnnMDH2RaQse5u6+6
JDdk1ussQhrFT4gdcKba5ic1bJuutTrQWrKitVdMsve/AYxrBskV1a/HsX7me4E+
SN9vLvVTP1tXzoe8CY6NyfP8biVD/7t6F4vE2mCfqT0GwnBM4K2XMWJQwmizKxa2
Ghe3jI1urjTvrZbDgrMvMMpM1lyU3gjTnJLETw7c8IbjcWlU2SellXls9p3Rgiqk
WGrGHwJK1UhHW66IvmSF9Z76ntwQPulwCon3tZjVceX3h3oIw650BpC1j+SFtbTL
zrU6Db6M8+5Zin8yUtKeSmkB7WRwrNdhqzw+xMf3YW3V18pABa+1JdyEQdYD3V7x
lfQpp6flF4+6DbMWSdiSCIdJnz3EfatuDhN+muNrCorvMIHQQZLSFmljsRc2qmyH
t1FsuOc8GAHQr+wRHKbbH1gshKCr2DZD+6+Ech3Cp7dQoskKKDqPdcSBbwNe0laD
kmXzlO9AQWR6peT21YHhOyCgGHLsXbiAkImjlccsJx3KbTMBVGarODmzSsgCmHCQ
6ZKQhrpf/R0asXmRtgRnJBrDmYdRN4nPZeJokfXhv0Uz+YyHNhp4uQA0Chwsk9Zs
ZTKYuRijv8ACT1IquxWzXDTebcwK+n3X75QRjzYmax0w8wCkCXJkgAxsAXRW4sFq
whChv/q+9zZsesQ2jf+hW3+8Iar8qrHxphotrti9sH7Su/4A3AbSqjEnM+o1r1Rd
ZhvybypmdxLTHM9dl6VWvrPPWxMtufVjf7y9Lg2CYwEempUkn07K4l/m1hxoBzbU
80ql0TTpe5fHqzdIN5v0UYY8+8Gm//fBxVX1qyyQ2WFF8v3VJodZzQsObqjvJWaE
PM5vxaoP4rGJRjs5020CpUzklZReSvw23o1oVwXuNySeDoATtbxpqGHbjYzDv6CV
vtkIYYJ96IbgJCj1xtoHwvO6/MVlByKTgm3MnCNTH3it40LYPxLcwEQN4biNl2S9
vOodvOYpKDaqjpHL1L9GekUi+G8cYTtQylhM7kbAUuivnaQXiLc+A/bfpQCK/pT2
Jf+wa4N2/PYR64o5L/Tmon/csGH1tv+x0ym7Yfr4VvO/2uJiXL6NsLyPBeEkuB9u
mBZyCF+Kb/TmAtLoVYe29rsZzLJ1xnuWQsmkG81oIXiYTe0BIyBvOvg79vv0ojMn
jvNkKFk9w2HO1H+Y8KPVhvcDOmJ8goGgZk5YkpdHkzurRSgfdMj8N4vXrICeiWf7
vdCblIWoy0yh5KTxnr+qhdEFDBLcoev0sh/4Db3jH95248VEdUSXZg4OnwwUCpvy
bJW1XlzwPJ6TU1qECyQi6s/CMj9k90wFcoP4Ga/Z9/B5VEdfm+2TqQP2FlaqUaem
RbkwIrrJMLIONWjeJLZca7OaJAfUyNS8B307T9TgCVd1lfOG9fVyu504X50ULV9g
I//hk8fqG+NALEu9Wl8Ban+Onue/PpeuK7X7q/WxS7QgxNhFFB4LaiPg8sxyhWuA
FtpAtLUDtHO+Q9KSe7kpKA6PIvXBaQncUyHvZMfFtnV71AOhC8ByaDMw8V32wOzU
mSSxDTIpTQjs/tzJxSIlYuH2cPCNV2ogKGwIPM0PlHk0gpg57hf0mJE2IMkMotLr
FDuLcQPVrvA/76XFDz7xsjDonZFec5ZKeVdK55X/sS3QFxKzjbCxeX4Dv38ED72Y
S5X5nyoigs7TBycy2DKJnFrNP9au4J4csZKrzkkwNYvc3NE3PT2FeqBbAjcnSkZF
nbGpRq9bqoX8iwELR2iuDWgHuU5OuCr4+kJJJKWowKHFkcH52GcruyeAgmO1NKN5
KBnDf7djNwianp5dTOfzM8CEvwChbhTSqmoqVIhFfvWqjbXTdV9Ho2ywsg1Dwcu8
sKgP+dRFZBqEEfWX6oU0JsszWsFc7ha0pXnXJdskdLKJoYTdO42NiYl+K9TdT++Z
5ugtmY5MmlbQRLX+Hp1sNYCttnPvpTolRF1xmqZj8jSvnRqiHcyh6nxSZwiGMxfm
5NnTH5GJiuiocnKpIHybMb8kvLypRJDJxqM9hYI2atAnB3VK3pQ2szBIB1CJUNzP
o82sczFnvjqAgHsk+914NC4bqPJ2yF+g3D5+90CaSG/cqfC22VUEfY6yrQxBNNpx
gphB3Ureel43mWcL/t3fynPvEk9oyFmW4PFUKYZhblmI97GI9X7h80+PZ1sIZenW
qnQjCmL8gkIqy94ssBZ4Dom5Ukei30QbB9IzGrRVQVyfBjYCE7OojdomIGmx4cqW
GGtBjBUM6t9u6hCwwA88vagPvl9FLTkHSeP2f3UnebZrZvjow1Yt9iMCN6TSQged
XFegEgc+8JLTRGSR8pxTYHPNZJ4tNjtU9zDluzN4o6LSMJQGjBw5wBRsNvYNV3DR
3dml2hFAWtpTz05AS/rysaAoBAD+RdAbUHhZYCggJWh5jTZG1BB/Hl/Id6MqN4YU
oMHYhNpMPqRowCLYF3r2P7bWicRhaU9BuQ9Rs33swoJ51Vrd4E0ewFiiotY457ef
rX4iiXUfothRC6h6g+JnW8crO3fbRJ+X719v6pd9/WfBzkX9RfDMwY/26WQCwC0Y
2UHkq2AoSLl5lucHmnKz+niun6v0dWNFCDQmg+iB/43ZqylJbPJJbQfVSRhTY4Eo
53rZVxdFRvKWVDg+14p4k4wQ1bMTh/GT6ST6tRkxEOwq0dH9eUnAbvToM3hrYvJt
w0WfnKxZjS7WmFkvF6tTB8V4RneSmG0yhrq4XqXR9K6uztobwMcLcAG8rXxMaMhZ
pMICfwUPmdMgMqv3erJc99v5JOsbYuBPJGAq9MEudK4WihNPdXy9ECxbI+HMums9
zzDd22ebSe3mg9Il0IWx8frdCXHFWPUg1LVhR4EH8YkiGrbk9PnNQ0FhnLnhR6TF
MOPzCC5+ZppKdWCZSZMo+g==
`pragma protect end_protected
