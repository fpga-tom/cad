// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lshcs3XwlBjzegdPvMamuKgiQnuZuTQf4EGqNje7ENjEiVbY0eAec/6zvVSaHjbZ
a+ngf1ybD07TNDPL0ls8giguF4eJdtKeSazHFfsRbePX0MCG6pW8a52OKIUb9U39
REj7frOoItSniFk+G5rvYJ4wyehLEHYAKZZ3lT2pj48=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22160)
wZ4jx28tSHY4HBHUU/R9imcKA6HKaxa4kzhTWM0NtOG9+yps8mqtdmMR+vcZRfYS
pfZSfXvajaGARmfqzE8J9mAhLY1Zo4K1Mw9eZpktl6qv1R2ke9qBJSO5Xn7XlGHD
elbqfnxg6AGqzkIU2viYAzFiFrH6Y8yJHEQNpY8V+NhIvJRympPZB1FA+m6JqSP3
1v0iIw+/QSTW9KcvKZ185txvzmaonIyraiLzEIquvgXJSvIT2VXjG2z6mWI8B3q4
lkxFz9bQheasoe5VgLrkBOQCrUISt2Xsc99u9pmPTKn/42BMc4+NjSIeMSZ7Pdd+
0ZNAUrnnNGlk8lw1JEo5q4NaWvzllqusTpGunvSN2fGZo0EeP3tI459lRKhbb1Tj
vEauZVozhCyutC6BU/bKY5QDCuRLodSsVqwVNfRWxob30UAtXK+q4hyjRiRzLhqf
+ePMVFqjpMy2RVrvfURedUPqO7td1onywIFskbe+PP5HLBhRyhRaHq7Efi8egPkW
3e6lKikIjyFfLeJi/jZxwvogONFNrAkgiToVkgAT16wTEd8XPTKmHVEkf7thqoPW
bRzzMBqe7I2xEHY/xRwBauWi3mXgvFvm08zvCO38qBr9yW+vkWdKH1yUfCKflF5q
K3X2WajBDoaYyEUP/wIrNxdGjZODu5bA5XNCjirpavA3+wI+qqcV9vo/yyvLQhsF
eTWQXsuzQfObMjWc0k/aJ8lsgqDa8T/OM8E4tpnUfeWzHLl+f6P9gzm6hd3OZwwK
IVv7Z+W4h6FS3rsU1G3DWYQXW1CK5l3z+dJ/QmdVaFC9Q93hp2iffUcw2wb1iLpW
Lo1kYb+xw4s11yqdOLpawZHXWxRh6AbGyqvQulKWvl0Oq88ladpUhkBMY+eZNZXU
Dt8Ar0hmGZTqnFoRRcdAvv4D0JcbCmPz0ghRQLBTkH3f4Csfp0nlT2kpzZb3Lg/4
RW7bBNbEbviaxcQUy0SJ/r13opVPXJj/TEin8GAXsfolyrZYnJUKbIxOlQtF5EDP
2JN0AEYPA3uHTcfihXueIooeAF7Da/GmU9XfuBChjhnk3ZbccINVRWADng9ep3Wa
2HoFLftbIADzNcouMHj70fYzSUeg1PYKqx0liI7f7kJFnp5/DnpzwG+Gl8uFAv71
WhCWkZxQuBAd2eWCYUOF4iPL5zIKRuiTQAQXHvBG2pgYApFdD1VRqMOLOuYXuvz+
TCVrUJGbEtDFkgOWo3g7UubSqN1lKz0Blb/ixjLRVsTvCklkjunWJ21qbXSgUCt6
cuk7Op/E8oMnEwn4xCBQOPOI/zwOEasnmdClYQDyeoH1OOLIfEiTN/NwvNSp+O/O
85TGY8kRwprpqQl9gi1sNB0JXIKg/kzTiO62y4+10PWogFDbajn2BcYtvWJZVLIr
3x0b2/Q5ppnGbrwAALxs+bpuEWBn/TJe8QdTAolybxkOI8uZk5b0NnVxourikpPb
VIG/wdtNqPg2BRueiSSs3Uv6eee94m/n4PtugglXpAO612GXf4Yh8iAi9fX7rjFk
RcBkJTNwAvYgljBvdpXbaAsgMcJ6kbYsZxvJVqpTaksWseu22rtsxAa8L4Ol/L91
HGm+VrdUi7PuSAd6q+IYslgqBVji/sUEakifgrwtDgM4DenK/f1BioQ9yNlnlP0W
tQs+0GZAkZLJncOI+pFRxA/dUytS4bMGhZGcwkB4vnnShXTX2+diJ/jK8PlQ8ytP
zxPyXKXBQiwTTxiCo2U9uUs03rJCn3uQlLPjGXMU2WJWH0zef8r2jIcJ48nh+BG/
gQgyR1IBSYJIdZKUcJASXw3dP6s90MOYdzW3QGDaQuPrZs8mzlt0RNu/ebjurmg7
Z33IFsfB7+DLj4dgw7KSlNJZ7MAUSPD9hdg9K5hir2srAaEI4e/ldaUbwkg5wov6
szVK0QBOMYd07Tu2aBvLvf3STaXKgdl72SEuPYwl1QZpAAAy0//HwEed4atvVhv0
VI+kIMGIFn8kfMy3jEon0ETCBQGqdF1N2D8+pgAGoQHZrGvW8VdboK3vk0O9TL7S
DH7dAKgCn4hkDbdvJXMIppMtZVx5GXgLpxGXRrrT0WkdrYie7B9kGe346566ci5q
E9imO5WQmB1gKAAeC9aWp0gxyO3t5XvHfPmkPoIX2uN3flHmT1bYM1J3vaTCep9l
5LgZ9iUIdBInwPXIi322ETBHta+SZvC7gzR6JmXH71S6o5qELKCKbHMlizqeIxzs
et4NRG4jTyrUa91Xwpu0laIPiZhjSg2Vp9e5Zcj5lKL8ZHU0NJi75rsbQmw0GOGi
Mw80uURxMR8q8dBgXWZ2LD+ix1MO/XgtkJGZwMnUIGFK0Qc4jIaNhZm7xXGgNik8
iqSiapehUKtZYb3KZ7GR/a/oDSP3WET/RnyPWXid/pQLgjwSUKdN73aWr7V5eCuS
qmRXXP4NBsFqtd5qPYMVa1cCneIgq4MgxTFT8bpLV3kcQgR6Ff/OJAzqDYA+RlFW
SSGD3Wr5sS95enpxsm7jSpMOrgKCsJzUA0H9+joCppzJVhBeG4W/LEvtOTeyZ9Uu
kWNmjawmSFYOtRimAUwuWTzxoAU8vHWn3NMOEwC4Qui9eRsR0fpbZciH+YEYXLmX
ya5VACPRMTUJaUoH79ozqXuCLuz1I72yo9tRiFvC8DQPCgvuKFryNHLzVAgu7ujM
yc6z8Tc+7uKht2nt7+5JjixccIlD7c1IVdOhWoeE0Nzo9A6jRQ0OdkUjir+7xZYo
khBlw0PJq33vHaXq4+//V7/v26GTYBs1onmL9KaFOr2+gONGk69uol2i7lyCv9Gy
j5kMC4097IR2H+3wC23V4LbtlOTJYLxwSaR5Skn59PB+T8WLTgU4nHFiMfjOJSif
M2MxjsKZ9MLXMSxMWd/K4Ed0GdfnPgaphZCFumMI6it11s2u/gOqY+KroCKX2ctw
ho2GSiSahX5NvmjQeRdPt/pX09QXJja8ywi6GUukdXm6PCb11j85UT63VS1fZbw4
MAFFyRUx1tMk/XQ+SYqjnU3pNWSFnHzb2C9wRA4HGDxe3ZyTCM41ngmKV92LhMGm
2FDRW2gZh0CgACqNUOq21/iI66bZcwo9m+ASO50xp0sHEZ1LKonMzeXTH9QTF8vO
1DOxDaf5Kofar07IEvtvnd0kZf/Z9TIjxvLk5r9ly4w0VK0EDXXF8BActmy4nOIc
s4Gb1hfIUWf26HvRQ40xIuBpbFSF0TSTFJK7tEtcaN4e+00j2HcMdlqjivzfSvam
ogYB0cQMXiHwQfYGX1s64aQrWK4vCRHCte3VwfrwYkpbBQ1v6n6VzEYpOZL0ZFWy
3eVaAOYV97+73tXSQmdYgm8VSwcSQ4RjkKgpSELcu3YimLR9ehEBuONdujGq+9gS
OzBoTlN3JYgSd7YWAbEP3fGNeNbSsKUtDpdn+f8rVu3NrWwQCrFcLDUaERgstnOg
28CBUdoYyToDwuE+GJQgKEq590H/nBihMEJCSZd/4Qi0yTkuN3FnFOELHJacaKCZ
hZr2y19rWOSt0WOwEmBaxnMr4egxvr9XC+GKc1Ltq+cfrA/93zAaWxgbafx5D7sF
9zcD/QJCtM+MsJqDf0Hx5Jkv0V+d8aG9xDiFixWftvvXgnQRO+WdIau29wRcT8Hz
wTNE9BHHVNu9mj0Nvqgw4SSiVDha+iOOC9gY/B7XVwS6sVdfBXOnnwNnul+2yM6q
1EPV496Q2Gosc0HIJwS+u9FViRXQ1/Oq646LYky5K0m4J8sQOZJ9IYtI/OY+oTac
t1/OX2W+L9Y98DkiBlEYdolzInjrfb6j/5c1BJdOOZUl4KShFgAnbNgeR6/pJvDk
Y7QXWPh9fSg8h5dzqC7aX/aI0Psp/Rb6/Lu8gOk6vP2cWRGQ8WCUbkXGV+ufcWNs
x0ksu+zJafiv9O7BpiczCE1RIQcW8UP7htZjLCgIiVnRGsf+lZM4exTHWZRYgaIX
nit+af9nqNPGiGzKpVPMDnZFRsKOaCq4TLBT289D3fnfwfRbTgjwdznu8drf376e
+Oc0pzcz4+AB4Dk2bqoFv1UrGDqT6W02XB4rio/qAYMEifnK9ZkdxU4Chn+8QG5l
20ubWcwlBqQkwIQa+K8Aqd6tXz0gOWtHkYQSaIrOkew7/JPD7RaCsecSwJpZiRw3
9OPsu6qrkmbB/UQQxko6BgydyVTx9phK/SmH/a5p1Cqds+VfzZ9fOZvub9nqrC0E
jPiFffMW6wbbrFsHADJMkHy11d0zLu5vms0aVlUKP9vWymxhGe1sGPxrrAMxUvPD
2xDbdBMNtl1RYCKEvr8UD9nf3VDmaFLeNo0jJeBc3TZdtNgQ8DpFe9yzb4n3GelZ
XGPbrer0AFbTdkXyEPeKaPDThQDdRkNZsUBhnOjvox9TPBpg9jkgYeKdq4dRfX47
Y7OcabwEZ19kUwnVIvXxLggtnpDOzIUdVZ5B6kptDzoWfBwB0JFmybtaoxmy/ZVY
nTmqIwRzx2O4Y1xP7UMXcTEoQSxHv7099om3mKKy7CYPjG8kqVVd7HZjeh+UDKxj
07DQaSFw91FU5jzIc89yzLnp5XDeRT1cE7nXxjVL3RXBT0iXcjokihgDYZdCi5Ut
cjQS17YEaj7auDnyxNh1fxAw5fAzCx07prYKNFmpoQJ3tPq6mofFYv1NsXIRbH3B
WZ7lX9zKL59dJSe4yc4jS7flwxFX5VqE+Ra1K5BTXiXdnzl7GyC2ZlW2jxxgPoRg
NCWIvQLeWOCUWbPKVQouQXhSTP4sSk1A9S3iy3B7mg7+XH2SV3AA2oDu6j89a0Pt
GAOsvVB9CP4Atu0JaS4aol7nw0yrU1TCrdIvgQDHaKFUapSPKGJw16/9KOfa9T85
aCT6XJrQ93eqCrXhF+YjFEQUFWA6JLlBpVGG1gznWLQxzDYR6fs9UpDAXe+cHAf2
ns8C2vABz+6h0xGWvmqLCB6jyZqkpnXdY+tt5VlSVUHg3m2/E758dMVc619aHe0D
mfHRhHgDcYLJHXO6cuzC9BQ3qw+Wq+gNa3Z4avAMb13N+LEFSFcqwsdRUQGo5fz7
O26B+PFd8+Dt8a5qd9qE5xk/WodTkKv+tgHUkezBMNIEpZyeSuUhJsBqyBUZUHQN
FC/LiSr7e4qvWYjz36ocNGfB8ant0S/iEcXOCgmoJs4zS9WM/PHUpcJJOJLuUKno
7JhLD2qu3n2AiP+Q4eNh1cndtwwm0KXqCpGOOBzuLPZfP06MCl55J2zbTraKGp22
8G/naIR8hgdWX+eVQvefteybUcxhNkfQi7pBoYR51OX45bYA1UCmWxcnEBRnZtli
ePwaGl6OuqPp0zDy7y5N461MGfKRHWK59u3Jv3PQBuu8V7nydiDDHaiBDeX/aYsA
TQV4tKkvb00KpDuvq2nrPt2od54q5GRK2TC+f0Bf19N/W2p389B/qnM0OId1kKJN
KG0THqdbTOZBg3cV0X9gLABV8uMAPDb0kdRfUg4vdSh1Vn2ewKx+W4vD1csltJ39
1IT6wCF8mOc+AEqEgR+LFkEQbAeVSHcJM9znyiSaLSG4xU2j4FH6MtuQz9u2DrJc
QIWDB8fbDZd/cXDw/C+BgTuAbC5P5rb0G2n0l9v662IJ8nL9xPEGYAXWO+LG0Lev
otk5IN+PxfvnM0zHpDq9aXV6sThJTp8UWDTApTEP+fHRO54orAtG8hDckTyA90rk
RuFrvvNQTodYjtwIHdhX9GldR1PIMS7f2cxw2yOWwuYpXL9ZFZe4R/VKIDtT8+RH
EI350mSrBHMynjcKl0ZuzbDmF136jIwMYDa22L4FfpCxIwgYUVDYuWKjZ3AxsKg/
WD6T8zuspI/YPT4Nvt8t/QQbCjYTroRrefUAbKmtEGpMBuT1KoM+VVSkf0brylnH
Q86wpdoryvTd4/EApA8naSLcKFngk3SMIZ+57F0kVKu6b9xE1WE4U9E7MTLyHSWk
NBBHXT/VyfsjjPQK1dXvU0aZSO9SqQdveVYSzSM0assN4Mz8y+QqkgpTKNPEo/JD
4Wx9Vacdy9uZNzYYQVqtninpctEFvYsprtJ46vKp1YgzBdYCqq30gOER3Tn0fXRz
dP1wCyCGfP9Dg3Y/P4AHr0tsH5+IzY0Tlb9pVD7wYeqfcwomV6S8YvN4xS4+60U+
k4E4immrwM0OWnzhwCLEvLipDAWCnkYtlDfPWLf+45ME7FZWwDpXpjqsuKiG62af
OB2wkeSkZqeR1po9mTZpZ9cYef/OLEFiHYnmBEJHs40fOrNCJN4dShRM3XhRA9yf
f/5XJU9eubzMV7BPIOY2knr26ps/MjOHsoWlIg4rsi/Vhepw//QZyFfIImJRPSTP
MWlIFGHj6mGQCQ80vUVXR9DkX642dSJ9FlcQ/LynGKHAslfbpAVValhMn+5RoVlF
1I/S2eqhemAxhgWUU2/BD5JJI34sBZPpeYfjyJ4Q9wSU7pKNv8syY8J4Cyjg3uki
rTJpSDGeCvIbs/uNQUWa8Yvqd1OfwHF6g2cEPZ/hAy8jxhqLdPlWOLtC65v6K8Je
dcnzaQIQaB4dOu+tJBZfjLlxThhgGKY403DrnUPpbUdfL7uMoRJ+HIBKt1NVQJt7
q2lX0XQVUCGOnu/Q/KT2SO+9kMyoUiHonp+6sKV8OGaRG3Jv4d/5vt2s9SMC7lc0
drSzgM+MCqog0oajOH8/eczG8+aSClxeRcYMZWEg8bDnDF29fjDCxKimvTtebwCu
KaEiBhjPJHXxon711/NrPxRm4Vt5al8xqsvQ3CrjpHO3v3LNh6NaKu1M3b9pUW3H
RfUHjL33tEWUsE4NmOqTNoVWDDGMv2Vju1fffRrh3MSTYqQRgCJnSZ1j3bl2BKmH
mAPlS3Ok3+iyN0XqGuFr/ljJphz/0lZHtwdJqLLTlT0kzsiQpbK5dEcxhZPwTN07
DzQ+i3L1NbpncwesW1xiQJrU1R7Bm4RnrhJDfYGntxE4EVQMJ0Q7Aaxn1HtJ9eYD
35CFxRmwxa8dHoKDYvuE10bfwlyQYZKAbz+DTQWkDR+Pfd1ud57gsxaY1SmDrz6r
hlskGGrfG0Zk0ORyKkFEeP2iJqOtHaXzDCZ+YrVs7oHbn+rGQgiLTW1M1r2NGVkf
pKfoNaLINl+rx4Aw+17/16UHQ+9sOpGYV0kIKHS5GjHnxglGXLse98dnZ4nW2/9y
JvrFdvbZbW/xeuIiOMHzYQ0k0vDPkfrSFY9llqUCc7J7jVXugO0t5DJ5A6eOIfJk
e2EPR3i1XUjDuE87T4J/JpNz3Mm62xe0ERWqSrlr69j0puIBmOKF9YYDNOLYyrRg
4GfckjPaZgQp6SIbGGe0rof9Ar6eKdw7XNDfngTIY5pSXQeSgz4xeoUq4lTOJBtx
gYx/7SkehrE7qq764YL6TFos0/wEF3anjLwfZDtRHIvy1bpfpWPHYL4WcT2x2a3A
OGm8Nq4pQop9MjhU5SyzGzGM4qkRRr1G2/ymz4Sa7D9U3m7yveqkBpvfPfZS+6SN
m0qtadAV5z92nCM8ckhW3Cy03gsZsTrupWrJ5WUbXeOhhU6iBfaN36IVd7viBq+C
T+tWzGqX0wQSXuzzyA9Fta9Up76ej6RiUaEpLr8q/Lt4E+NL/3QXO4yvrc7Eibl0
jigdPvy1tkmCJ3waRPi0Su9k4ucc/Phz2kFnv1ZLazIuJoTZDI+rKW31SI5JcDWq
tZIatIbDYDm9c1rB0az/RrrYgZAAcfcLEgPGbo5e0TKFwbIB9z/gtqasn8ZHs7jq
1UT6ZQ/77rbT0VJ0wHjR58hvnQRqgsYw0F0F/A9x/YLUvKT+mbeMZ0bSCkCzS7v4
kpd7XLeNEjQXDWImBbj2OYxfw2jsq5dl9UJKMvmq7WdGAXGgbhvMUSaJlhDEV+C4
uXai+t3GXuhwVDJN01wdLNFtfYtKAidN7FJneKjgLx5a8AWoaez7VTq3ZUPniZv0
mgWxrhqpBFvXq/dHuDVij/zUrv0vWVCX7jC1b2TJHvqBIyRHB7UgYh7dDaUdxVXl
opKvIaUZz/jKKXcBTBmptX5sBRX0ltEcCEshHed3Y5FOBnXPRuDHKs5JO5cTL2bx
dIL9XjdwKBFqNMdX3+Igo9lgBRKaQitd/IGNZg00tRoz8iB4GAVAyB61UQ9to6M9
LpCP/goL5ZE+JQvxAtx5ISIGj+FseQDmc1NuyOHz/Ww67GuN/oWOf0+SUVWYD2dL
rhqLFoqNLXrMiz0DGVNLe60xMfqBEwkxpnm+UhvTFOFhPE5EpDGMmlVqMo15x6Pp
vRwuXp4qklB6TR8DGdtylT6E9fjWN8wD6H2rdkr/stcDGb3rIpKi3yKzHd9Mbg2c
uKVSwMn8O22gmObn3lpr9NH0hlO/AZJAZTBi/f7MGUsjS29K8D4sZA6X2FLAzgGh
tvJAO4p45wgPDV5l4+6+KcPSovZZtq1jMPSYCu1nbjy/D7wC0QTDRSkyGFXSUWyg
XWTkpRn+SgKnavzjaSSQ47Aw3Ywu0GVftXmVvJfZ52b9CKKsjfISXaGy+kBbGVTP
CRgtCxUiOwIdqYyvJzk+SQ29/ldsSKdqR/B8TS5LJVspUChbPnMcdbx7W78ZEQgO
1mcEIR9lyKHsRJBhks6vI1reGZBldlxRqw6vlhBNqJ53TE8kcE1E/b+26RmIH/yF
LTnJEDN5qzGrEDdysE09/UXQSKNot1ZD4BPkXJSL/9j1JlajJNwg2Q366wHP25XW
yHSuNN4TifQLF5u3gqbQfDO0vRE9wAYR3JMh31SOxnYWNvNbXMgYZv5XMI+lU+iR
GcDIXR00tWtWV+Oqjbt9dddjjmcP7e1ChU9MWr2sGeawl9H1zYwOBZAIciQ7jJXa
uriaRkcL9XJVLTjfuW1U9WAHjGsonXU0I6qaOXM00O4cZrpEpVTVhaiOUFzQR2pb
fzPrlH8pCx4cClYA1DYQuIFxfOI/gof6JdQZnZGqpUMXuuCv5dR0EwSddNjxZ/EQ
e70zudPWnShuTG9zTiQJN4qagryoGm0Gn2BeXM9j4T8jCof/KExxUQiW7MdXbPA7
IQ3iVKTq6koKkmJLgfM70jX506T53qiDG/pg6mgl8OBEqw6N0Kb75fZqftb0Rd6b
dvAvG/w7O9l/AE4D63bF2SpIWfQzZuilndP69K3s0LBOEikTMZ2Qp8nsJ0Rkkiqh
PxERAIJ5a9h4TgUu3TehnncWXZfX/d4BEkXoP2KLYaCMl2P29ZBElv0ItUoXL2ms
RO+OhvAlY2KBmyNQIUh4QHd/2b4E0W6ucuReIJEIY+LAkqBSfOxVg3dt4P9pkrt+
u631dnOVyTWEf8eubJnLeAQcYG5VWYdfyxtii5J7svpLtbRH9fzYxyyHNt9CjUYi
B7jUC1WKdZg9WA80UJj5tcOSnP6f6p8dlCfoR/KbwieLu7QiBaJkoQOPAhp9y6LP
dCR7UOep56lw0OMBchvE6sXLehBIUbRwXJY9YyO46ay/UDm9gyBDHSuZ9uYdG36v
V0Uo/jV2cb4W8eiVheXOfAKtCYL3ALbGylQUxp+M+ADQ7If+tUmpiuj3fxihhkUN
JQwME3pEf8ZrP3Q3cVuU+t7GVUBWU5Pr9YEOypcpqFzyUp34/eIHBZkI9LpxdYm7
3+T80VtXpPfsWK4plzJSWBuzWnRaHWqU+xdK/wYzIppN0O5SY9d3mnManpylYCqH
4AGkUhXvJPUkQMHEpC/XtS2zY4daNB3lOzCors2ClbJtFrOEmrEzINR10+XjnEj5
e3Oqk4exWYlMNNBqiT54aTuF6zywnlePyyhj8l/CaY4JghBDoSpk9zHAH0PEBsfn
n7jTjYzH/D19xohoo+9TvsHS5lTeXyUSv1eSqT/ldyZ/UZixU3/zLAdJQGZ8q13Y
ZvCEFIAHuHbz+0MT1yl1hdWJdlNsgHPPXW5+IVl6Dfg4APqvrb9jmogyx878lcWT
qsjj/aSl+IXDleWjrkdrHkgTlyGaiimACSEpZ2XCS3/N9rWsIDTtLpCNNARrn5Ea
FQktg4m+ecoZCTa6ub6WByQIa224+bNP1uvxOM+SSMnu3uUe2uTkdZuys2/N3ZRR
z5LgQRuOzEQiMQjTUlezP49+jP+toFYURM3oo8kOl0IMe3A/EWmtNgZQJaqhdVvl
FRNRXiNoXZYqf6ujdAG90tYXQrAmh3FbvR6geVGjLR2JkjOMh7nKauyopVPT9iY8
IIEpnamSqQrAGgc+6AxOXtAERj4kihJvqaSIpOZe0oJxB9VPlsX3U4WhDiereU6g
MHB62p89GBUBKXgqj0waEJNgH4IgXyg9R3U9GmCZKCzY9Eac7FyHs+oxeNJ95npr
CkL4EYQ8wC3LsvjHxVNxhHze7TGyuErGADZlwPKFIy1hUtPr7Dz/RQafegRDV/qi
g/FtQrFMNn98pe6SD33oQwJrOH4/lHwuGwLsmq80xPt3/4N0Kpop9/GfdxjNgs1A
2pgNn/oYTGhU/zO/HkdQsSYb8KTGuSgivn0Dwgj3+nMu05+BwEDQ3mj8P+cOzWfG
4nWLox1A2BrNimmbRKOMjJxCFe1UPSUrQE7CGZkCfEOmwpD5Sies6RjUav1aLYMs
3VFDip7j83oKoajU+vwV5rFAuA7IE8eklsUtkQy1Exx3XrxvS7CAD46tSE+0WBqi
5gqM1xXybiYCWNlZjrdgdmx4UOkfMF+4TfCMWeiTQtIaMrnSt7IEb/81UVYpAo34
geY4TZIVCoLf8MIAwmhpd2Zze+id18KPdQCun4h4G+ASaOk3NMxcpFfinoS2EspG
BpIKdutHaSq1jFqNApw1imq9sQIfNNSl7948zF0vU/d5e6IxHJMxy5xuRpZvuDEr
tE2othlJNJrj4xUz/fq8+D3byplYpyShoP44sBgzRyORizDwAvwIYZ/nGBqeI190
WN+++qsd3FCRf/jEgIi4MrBhQ7vWByWqOXJ3H9bkso6yz0AXl4+b7zcPVRIOUI7r
Pfdq2ohI2n1BM82a6PUinkrkW9TUdcJ5Hkjvg7Vbkp1BgEJ6olafURmCwzww50Pw
TejvxMYs3O4rG1Eeh1rbtF8DfhBe+wdyS6IV/QwLGAp88REgPSq0D9pmH5gRQC+1
ldHhUef7lJIzDJwvKZRALlvloNzB0fVND59tdGVNozaUSdf7XnXmFYoVOJCtx88D
E+4yi+zuKPCLsaBjcmX5IECWfS2wWHfGA2AAkiU1s+TzeMEqKYZ8/UHWghtOqfqB
doUlGx3SNpW9ThKOyt60fWwcidG08VEU+PZm6kQqM1rHLa4iNxjgE0KU5JVDBHLc
ddhhbUUj9KjyVkye81QMFAIErm4h1sUz9o8UbvmA2zPRZfJLrBI9UIAb2acbhtBn
aCDfdUwoDDxyzfvtVRZI6IC+52aMCd8BLTP9y7IWmImwV3Gv4cNebZv8dfXG1sSk
B1mYA2vWmjsDCq5p7FkFGi7uxmu9jkv0KJzuOvef0zEh8m8lsOKIhaolNcxs4GcD
CIAjREl4415R6nv3OjprRUB/9cHqAqHXjd/l+DUOG5gyYuB7pnhxc2hvfhI9qsLr
TDZeORPCDr4lZpbCG2UlHllPkM0vtbLuAc+ES783OfDLxcgXo4DSy8tq09Yc6hlN
MN24Ss1HZ/teJQzwWPsjvxm1ClP5DGe7fTg1vg/xsPG2z/AmQ/IlpBwg1P6JiEzo
fEx3JzEgEdvToAtLEw/IODIq1tHJ1gpjhgxfFeWm1EQICNweXHOxMRhFEAQN+jg5
LfgkTSU0BB/j6lwQEM9ab+82dXWX0R2Cjkp7TAuTCIeyIrINMHeCRwY+RyptIBUN
9/kkmvT3cXX1yio7vSb5a8xa+NxIKSne6Y+40ezz4MEe/kSdxe/oi5oQoerPp6+L
BGkCTFb9TWwy40Q73Et1fCqCT3202mlmMzvF4gBpmTsVzI0Xtk34IXfF0Sg3RQVy
7yHSLX1GCVJGZvUGayBy5GeKzm6OqqZ91wGhHoBzb/XSf/Xcc8xzylDpowpQk46j
fFHgBjzMgbWSd7W4VhpZrT9Un2cyij53rAyGcVqSgJr9UHMAAryszPgye/pRj0O2
vi6k7cTsSLvmhdDqK0v/TbimUM3tsYBM6vswZD/at+ICHBSxXYQHZ6B2gwZhwXB5
tBGI8uAPaWFmD/JWlnjmMj/P2ZzgXs/z/u2vxw1qwv7D/xJoRIxDfyECeSESh7BY
wf/UE9uQAqcDEr40Om0eKzQwxlGrSWxgvnVCKni1HIIL8v08tHAa4DKlH+SdE8VB
5qRCgep7JIId9XIRXHd61FDk+t2EcnBYWX3huTJLPhIYejycryRjXZ8GAZKjQqEy
nLdvxraWPZ8aCKgYa7NhX4jdBA77uZfzX9k1cMdRTbw7aStPixZQ/ZrDeoJrop3l
c+p6MvCyicYDo/buVwxyYuXB5SDT59c15AgE/ERL2I9gIXQXIDKBZRNOmyAjvQg8
6b5mQa2aTMK64JK5SK5sibj2phjxOg5CAtJeJbvWo6Byjx1LvaE5foGaWcT22jR6
2Wgu4f/PbOw8QZrcGKLc8B6TDpQpbgRb91fR52ObPEKjoyDYCgm2RMAeGhlIEibg
3y/1er6aETXVAtg2tJsMXp9TseDZI7Gsgnjmbwql1QppHvoQsA6U0IM/DAI+YK98
ZZe8F1akBGgjzlawrLGYAkeXpKLMW+hKlGOiG0CcDUu9WCOA9FBU3K97wxmkL+cV
gyFCtFOGFK9TIs2LDTr/zpXQu87iBGk9jaskjWibS5LirZLSZ0ti7cLNqu8rk+RW
j9Q0tHjiMZv6OhyMIPmQUL0MuXog4QyPAQLNrdspGrHpne0Ijiv1336JYoZwoObX
NGP75FGl4H8E1cZeSmUSQME7ixrt/Odm5DNoKg2JZd6ovW68F6VZyVeBwyUOvFY0
QK86r3NZyE4BTjT5MmFqkFxXWF1NSKZ0bp1s9a693KVi/nOu/YL5FkOWnI5aLNH7
WzJBIKmzXcyXnWBnwbBKK77uWvv+wthMxWvBKi9z/vdeltRikgGJN15r1nylXLoP
8p9pKiAIFpLsgGcswWTHzZkafuWWHzvy42UPz+MVVH7SJJ1Ba0JLvjZd018j9Rgi
FHkO92a8eWypw8vlIRCTkCDOs9vfIwGmvor7yIsWIXXqYo1YiMhH6mFxs2ah89Xv
IklZuNnM/TNK1CucNU4WleIXLPrEtYeDy+qcjVi7oSEq37f0Qg8CsXPmypvLgeBJ
WtEvFaFyTppthHprOorDXizUISDsckfEMTfGReAMVuPbo4cPD8HtCdbMlRqOe6N7
VCu0rOPp5tqFMFvVXOmZ/l0oZxretOgnRf2zSCS3M7BxX9Y2yKFDZq3rgT6wwoRh
qEdcNHVmGTU9cYLRfG51I2L0R/jgZlbz0wWJDJfoDYIobcRXmaf8MG9QSJaE/Toi
DT/dvi6ZqcQyToo+33Bgsw2vtxApkkntGdGg/RfdoyB4lLYuwGt/JsujtqBFSVtg
ld3v2n51QNxQsnObLEnpWN8eJna6KWbx9FI3qKyEsRQqeABc7XWy4U7bxM7YLKNX
Kn99s3wXCuwEzvM+W6AOSxP0Srqgc6uukQba/0xw0yEVhgJowoUiIDyOvmpQRRuG
5Y+Ln0pugSHNGcy1buMg8+8LhNIxYZeNNZR5LgjwEosybjsLfeKjXf5Cwea4pEKo
EIzXszW6I45ycJvd+Lpud7EliL3BYIInJqXO6BdD+JIAV9ablzxDmD8mbKulbvkb
nS4YUWtBT2NV7eGB7h23XhaHSITiRYDOWqT4NvWPZnLqEzo4o/Z5qbrbpT2joKE4
rc20OCR+5EqfiyewpxOBA0Vy68wWJeKgUZRDSBEgm9BED2PLrZf8XloeU0mWdkmS
3ZKPnkL5+q1RRJfnm+d6FE6RJ8sctMGxstRxoK97alA5xipq957NPjaHK1dHloIS
dC2qI9gld28UUC8WmmPiact1ueEtCybXkm83m9J2UnGMfcmIbZv1lbzee2xFXBts
BAYf+CCzuZo1uOMOkhXgiwLQHetV2IWfzt67V4kptdxksSSKUdAbMZ7QPc0S+5hV
uafp0TBTczs0GbJJ+SDKDT/HZfV+dk01yWruY8JvVmzsy8tNLQddXlUpxE/9Q1GQ
sqH+VFW6c6xmAMLJ+mccfgWM3EUPNAmztrBupMlj5JAeXLHnkS1SfRA4aI0f+h5r
+k+7VWr4LOI5fZtuUSVp4TiR8TQAnOElYM6OGTB4TJdxGg82nXCnlTFI+NOzbbcN
+yGQB8AV1tBuhsLWPoBBxm6yoxdvSiQ8TMZYsre/SCqkP2+uVcDJEpCm4jFZHsIM
0i8Lku8HMz+IUaG5oJyGR2vAxyezGXzxEOfOwqeFDeVHIb+FML9aRgD7W33H3i4y
0MOSX+6kQK+BVJHevEZSY/GYhOCa7Q4PH7GlAcVwZ9Cu/GLWC/VH0vFGOqdwv2mB
vbD+PcmuT3fbL5MI7VCmdpvVv67Gn0DQ/J3g+RUSYQR4AK5jbtkj/4HhoM2wgVo2
RGDuivV0A27Gwxif2549trKIy+AyUM6ZwEq/MLKb0X5ZYuWc+/y8Ij0jJbmmpmXf
Rt99/Jq7JoKcrtwGvDwb2mTmPoArUCf0gr/QGMrzWaAfbTTyZAYGJyH0O6/A/XhX
zizyRteaYm1+jJmMOL9IjAHGLbngSdC0aQdWY/jww+/Ph3bGNXCvSvQjgy2YTEac
ScUdT4cQb16o9k1zadND+a+N2FhrKCr+IOHEfJ20QCuoI24RfWOsq7OW+ZVzLTkX
BuMdEHNY34iERQwAu2eWYFsbvzHnoSbFHxHVQANyG+eZAWobykhYqRsSBZl+kcrQ
fj0S+q+WaRhurJrc+p6TMeSTKsngWhnItlwBd7TxP2afk4KwEKUdEDa5VlVW6QBp
VoOT7TiMCGmHBZ3GoM6RVOL0c30gBdq80DKrjoj7/Q5YqGaYv+ozvW7QgF6j13n0
Dd+vUKdwNoY6B+/+jBTQMwSvEeoZxjz0K74KprkmDKRaC0lrlYw1lTFotaNC79BB
jLyg39d4mTd656J0Fbtll+pihOnrd46HudQAXkYgJ/I/1oWNexLLLWgxpYDIXs2P
wSkq50JqZ8C/HKROjZR83xklcdM5QjS7iRPrtuLQGgaONXTiaTeC9/otVY5XQqBN
41JljbFDqIK5PG6RljaRdspwL1zfaiNIjkW72Bq32CEpNGnH514UGHZJEkXa5zfm
Wo1qDmd+/TfoxMjGJTSAapFF9Cez5gbS3myFfgbOY7DVO842fuYEhjsG2S2Huhf/
LvW6EpxftUY2Cb+pQd6iu/oXog6PR1veTkLXWbpXWmWvzSjUEQVpfQ31mojTHGvF
Q44QMqI6hQaIpnw2lGvafUt9HBIP/ArBg9LgCgjM4JoZ3dR0cSOdgh7HWm/LE4Ih
K6MyY83DUFZpyWKf38qdeIfI9NZSKD1IC9yE+TeCyPoqPyy1ZvHyUJPOBsBuyvwl
KPy1Oakc3hI3N3yXSmjZJYOa7i8nbDQ17VB3rwX4upbScpk+/kHwNtEfy0M46Rmb
L1fC/2EOBr7LZ+150cE7xWrpTw8EkpRpwgTvBTGRzLlmWTk6rLbJY0s33Z2kC6lY
jB9Xzvs82h4QUIzN8m+JuEEI95SmNyL5P+Fm0+/1n1s69Y3VlrjIEl4wWnBZ1F4G
YTyZnpAdzOp2UXl79ii4Jw7w0XzsAkwfxirnul2Ep4c0OWDtL0sFyVBWiI3vftKY
iwkdMtLvCHkEbN9b1HCOv3/CZm87vT8L0pi8Bu2SDDxJnYV3oF5CoiE/DA2uy5Gg
5WxGjAc46ZkREG+r8CClc3K7nHZmmzL4l9i98cBpLxVVu/iKNhoQD6AEbY1gyAA+
7VPd8JqPaec1iBX9v4EGTr+Q1DFPhjc//LYZx7zueaVPOKI4rgLbd1ei51+ojdzJ
shkhpBMOEqRWOBgtQOP33wnYefUbiWJfGQ7J9TArvKL1kqqVBo/tzJ3ZTwFjowjo
5+QHr1A8FdFtPIK9OTlhq8IvhCr7SIxlKDWPs8pq7kci+DhR/Aiw+GbB7iGgOSUG
YDRJBKWpkjCKMdNNX2fbP38P1BJxJHNYZ2/t5n3rTKHn7ffU5sDQkkSB7c29EZf0
ga3ZGNTZ7c60xI1S66Jjy7SsEXII411HaD6moVAIuCsB3eVYwdAdtwIyjAso/Ufy
uC/k7PlUv/9jzX02TVP8AnzfBkwhQJka2spopUNmiLfr6+KqTion4fF2k+Dq/V3s
2ddR+eCiAVqro+X+bPAQzsfNza/FA3wbXjz+9R3kFq81zKbDVXpeM7oTjhP6pME+
LzIgENLVWvKfI5oNRiz7U2vJzXP/M+q8pYuLKDLmloKNXjOCy5SraLcqqmfjRn69
rDbuwozzbjxBmbH8Pwjn0avn8UPD18z1tYyHTWRvQ5SD/b97ClUzhMGnvYE2Wjzb
DlJauCbx+K8IdY3LRpRMx/0KkyuUYiIjszbswDAq2Q3ElNbrCYMQywpUM0puly3B
LpVY0TrL8K2PiHEZDUOGBBcRQi8i/rqLFdb46vQc8mI9NjnIPfkA+3SuHX7msgkm
vSB5PRMum/UE4g+FxXbOeTJ920oG4stL6mbH2HBv5s5NrNQx3pwLwFrRcN+8pUKJ
j5hfB2NMYDZO1o/Jle+MCCaXhwWivAYAAkrcH8frvQOg6RU/Bd0FLkVI9bx6EJnh
vjDLXHcFAV8RWipkQQ0MFZYYs/27cwDijT8v72yM9Cq+/Ic4Sc7ycEo/V7DNfqxq
/sklEx9lxTrwq9Is9Y6zwLWHRT8OiGoR4xXxG0VtWAvExnI4LvzgqkWqBIaNOOKd
wa64tv1gTjOp14nEExkhgVjx6GVF/kgwyuGDCMbJV8Thwucf11028EsV/GGfpfkZ
drRPOJlUoOhHwAYoNwHM1ewXoVVCqZO7joKNfSsOGyAjOro1NjnzJRMguWYjoWxo
ji5f4AsdyJ+iOGm3H+nBL8Z/O2In7nT15lhEmjgMEO5qxBYunoKF2B1wGrIimIS1
vlsaPu5svNfa8Z80n7Si93cj+lDf5MBv6NiYNgChU8r4j96UZMlKYEXfj+nIV5iR
CNsky65O6RAC9xO/o1ZfdpXgtZL6UCatRQxecYSMjaZw4+E1V1RT8fdMImWYTYDo
9IQ/T6qTFxRfNRAcKLbOfV3pCRpicoLlfZX25FLJfWyYsVFKAEmDNQOgpT+6nMcK
XC2LvAOAXNhKA3Bqr2+94lfWaPzm17NTck+p/COIIui+jwBbOE1bYGo8wzXz/r2n
uXAOi1/yEMKYxcNANC5nKWvTxDYtNC/7Mjpwmw21yfVOV2r9hn2pITKIN4HKKRp2
4kBJiZyJMTcWn0ygzZ0p3wpXZ6CbQS/ctack+ywYQRMMjmhzWkFBEwaCP0yOBagr
YeWF/RcztvPt01zhQOg87HigkIlFmVcm1GxkDNs8M0H30fxMq00kgUqDRc2CskRD
YX41cgUbvuN6Sk0CNA0ES9J6vlZaDKVHUwXk7fugCC9f8bW9QpOuMlznj6cFV97S
0qWqEkQxvD49Z9aDitAUagTv5AI01scZ9Y6DniXUy3dKEATMY7+xbDK2wIH3MaDu
WF+2pELnXwH7x1O+i5VEKSdt2kkyUpkKSwWQdzUzjQfbbRz3Zc4lNlN8QNN0r5JP
d3tJsAzvrDeOgx7Hgd1Qburvp1UjaDNavSIh1AT43Mq9/I1cYEzTFNOzi1x5JDbw
bdWB0OTievo6Ym7Od+EFThQZ3fuxMOPNfBse1Jd34jBX5qPWB9hmnuaAeYiqCJWx
CsdKw29PHFcwyqTtrL1rKCvdEcon4Jqq9nyVNfmbHc34UuA8Q1+smQVXqz7+lT5x
+BXgeRMGBroBI3LAXCwMYXmLWbnaTPlwHqhkYy+ctdwPSrr5QMaLTHcjr/6RZVjF
Z7hv9KA18nugnuP02OaxBXUrrQ9jaVPXhRcJ24Y+IazYq0aY04KmqbgOXUyRmR+v
WyaQNh55i7kOXYQrwNZkVIFM0RiXpk7/i3ZWdud31H1HlXZ4YZPNXS1YqK9V2qn2
7mJumyF3KB3EVCMNu0ypQ4oSlIqrnBPjSs6pj2alw/bhMR/coklj7y27qip44Lf/
jQppO4V51yxJYI1CNiZXUHbMvlbKuPogDHyi9glqtCZQIGu8Nt5a2o/IK9do1DkY
xVv9k5UVvqJ22XPyhxnAM+x1NE8ovsB4TWmKOUbc3Yz9yrRl0W6wXSq/K+m5EH9F
smGOq7/PmTN5sPHBu//QHTuxZx90kLz50D8D31cq1sAn7eiVc+WbnjYVaIMri+Ri
Qa7ImU0NFyPrL1t287y9pKKAP6xvLC1VAbIgFPfr6XZIyGBfFDTKa+78nFZmvJWr
ERNDdwQ+zzT1dtIheDhyGOjUExrogi7IMOqYKvrDvriJ3jGGPESB80vUgOgXNiQp
XNFbW42fLbjQIVkKmRPIgIZnDxrfSja8khPxtcVXFhbpYDmi4HWm7FUdLtBzQZbd
8dvUiSDXR7JVsNziITKRnmyUqgwlojsXp02da/UBu3QFeSNWefpneNjCTCOa6Vu9
PGjFmBFZlWw//olqRNtXg2QARzR8uKM/s3kn5ekGTMSD0/NUS6WWM+nEvJJq2NMO
s7vq3m8HIE7yjST1hKbCHLCYsEu2FCO+t9Y6gZ8n3jW9AfyxVa3U++tllWCuvqR8
RUchHZWoDJM1I+qX3BB4REogJF+18jR8WdtD7d0A3+0HGURlUSOOH0ksrSLHU8EP
fdlkYArxb2S6H7dWk6/wuUJelHOOUfrbO7IHig6cejDJqVgT62YRy/XXRbep2z4X
dL8QEHEpt5zOqMJADCdrkhaG5e9ftHtGDDzD5RFJo8Nhy/qxTmLs3cmOTvYFfBie
wpU8xWZLujS76xDPSW5jD1Fx/gUkEV+iW8mY9HqEiylmH1j8gdyyDIpbz42JOaAE
Fe21wIMfsfCWqOhkQ0gCNWYYkxfjBFHAOvVH1sz+uoUim3RWI2gBtXkegplS0d/r
o+wpgJN1c86FHrTNE3uHVpkjFTJEKv0Wh5QZzn5gQhSHtFJPM/fNVl/DspCmYUDS
an2rNgfzeBk33InJnJ6BDBxU1LR2CCayE/AYoYyd2Ncws5aPOlJOuHNxLChmEhYj
8lzLatvwZxoeUZG/c2ssABwiEDe20ltKSDk7dcBB8OOKypY8/eSyUzAq1exiXU5j
fJO/fz4Imtx6L+0Ll7bguRFKeEeApUZcK/9qMC8Vi7tBFi1how5Gi3y1VFVUtxQW
EMqBpP7aYnBnwJOvAmlJ5MfH1L2a4uUCH3j+Lx74XE1klXeKRqGWZYe5y9e3A5T/
vrF21Fnv7GRikjdD4J0FJOxiOSZRT6K4TfQMVL9wwlR3D/v2nCocHkyeQ6Cnd4RK
I2t22Slxyr2k+PeMQavZkPuYpJH+0cy9nswfmmf3bRUZPuFuk1+WygRF1hLDaZGb
YtN3A5MNr8uDP7el4zQXCTCHK+zpe+Y+MPRB/qptbPYnHjNlAOOClZqdrxS3IcfG
4isOa2fMRQzm4xVnxdzhOEOEP5MGjLpzw/FVZQrS5cgr8X5O5H+0VJf8W0/GGBRg
GNPT7VLKxaTvxvEu1uL3NdCFKrMmyCLaxBkr1s2Y0w9eRdNgzhmoSt497jvfjwaV
V91qfBOe9QyNDHvjuM62z9ZXB9gZ7GGFjaRIshgkCdSPy7XzbX5rJEE+/Qxf7k5O
vY2kNmKFAHn5zmHa64IMaC5S9FN9eWhMRIXRCP7RtlvOTJV7xFRdCpZI1KnIeUxN
Fa3wJ3q1lrk2aJ6luBS8/QB9up9l+kFhtXEpXiK3N2Gg+r/2TamfEPVwMVxg1sby
o4aEWfs9+CW5d21j/nk88P+GZhLOCu5DNSG05lTe+70i/7vBFJXJjzurSUj2LzG3
gbS832pcT82JEOEhtXSdeecV7rHiFj2DarP81F0P1PnSCdFdzB23R07Lyfl7Xq6a
1Vd5LpuFl0756XDC2medqML1L5mbmPt0/PYt7r3KgQiSf7UfzYtUm+KjZMvdGFeS
Iu/hrqxIAra5bFi02c9s28jGMESTHXMvnKqL5erRMp6y7XTJ+ozutPbpNhXVA7hr
JEqyOk1nKY3/o8LcUwnkoFbZT9d9fk3t16zDHDB6JiasSS9z2vaEv0c/KiWK0mID
ta8HYKOM+0+PCAsvPYmBN9AQuWFQj0OYriv4NxGMnfkZIe7onMvW76mA8/lETqMk
CRgGD1OrNMsridfqh79j1givTojOGM0CYu+IIMb9zjjvcHeSdX60UHm1BJKT+v2J
xd1LhEBZNhZEbbQMyvak3LVaAWUGQ5UtmzRrUPHvn4r3fCYunvcz9w073k23K4S4
o/+DPtptyeJu+or1kkI/RURp6kK+XNx3aLq5jDYWViIfX83N/TcApZLrj2Tp/wN3
KLnYwQaDp8CPVC+lYh5ZAU1j+plEGZdYY8+I+QefIjdJgAk3ln0MNfj6hKTUuIvV
BnRCahVgXpinU3Uw1mWFpNztb6PAnpCqxdLvXJTSFl+zcRk3OnQR3Wc8OLJZd4OO
j1TKb7erPtDDgF77GJYoF6vGUwfQkcYNhROdHYRFkCgBxaQyQQLDmDblfOLVvgiA
ciVdEM58Sl8Oqdubp2Jpzr5C5//5Cn2i0UjHnGlUK8Fp2KaPiMFNdQzUOuaqTS+4
N7mvBYzNK0pvDoePNuZMm872eyYZgPORuXcEF+iR1xRxD+AqPmkRMreVEErV01Ao
mfM5AsnONMHH8XuXZlcBWlznCgjDqKvGmrypHILoqlZsTj5sgnH36vjkMpFcCvcY
Bjq2ovZlEiSyHiCFaLAy0q1UkJsYCLcVncUyxZUEEuNyDjSfn/r0xDBmsReJZ07T
546sQeaF09ZWBZzNtKOPuWu15ysce/IeM66uZ2yF/r5Rx2PQdxwKuKvXcLsflSrW
9ksRKOPdmC2NwXCK5kc7nu768WTgYRbauWRcxUZzj1BkklkfL8F8+u8sX3/3WhAt
0KeGx+94lFvC3m7pR29cpETR1t302B6qS0Z2P0yORfIZmkeLBs3EjSOHKFshZ7lm
+L2RE2ev8vyWJpcTGuAN0e5KDBvzqP77Galszp1FkeNWszyhUgQVRJJn2Az+r2e9
3J5yPFDCXzAFznSFAiLTVTmug3rWzvBWXuSD0/wCJ7glLouo2bNDLQ3yhmK3WAZw
45EPSgXdudUYFtnsZ8K6nbQmheVyzAPEYOm/pIgHPPI53YstAnrHrBoLWb1di+VQ
YQvl67XP00d7ex98+Ip+sSR2uSUZ5wUHnBLI01mCbJEZ8SStjGhrgP1y01NwD1GC
KgeYQoDyx97d4J97rIlM/LEpgsodBd8GhwueWpSAeQc3oa4hpYxm9pfU+3ICH+Ir
lJ7AaUD0aIW3R+5yWhyf5+HLDoB+HVEtJIK9vgsOQHPuPZrkdrWCfgg40KCW6ALs
H4GnWz4V5wqnNVywF13hXX0YFUO1q6LnyOUoxF73sN/f25SqHvmOJ+vBt94avThE
lMaPJz4PK3aWvKsVHfFM4oGlMiq2WxUXKVQ2GXXpbRaY5vLtXZquRctl17EiUyj7
dg3Q32w/+h7c0pIIWeXc7zHLYdmhNAopQrv+z02R8Dxmz3maeh4w+05niIiu8MMI
0VDrLhVDfhbnK5zAc6HFu+kQK0BQzTOdMmWD6XznhuSjfTKzzKvcE2QlJyckZRnz
0OWEPx4WmUHF2peJt7z7pfKmtvC0SCeSFKcSF31GS0Sf0azLJaC7M011dunNgspI
o2yHyc7QI7xcmbjHYIjfL3EfmZXSW+1/vUIeARaB90agyLiUkrDzl835aUien7Tz
ebwmVVYrYWAHLPrzRzwHWltOmBnRJQiMOwRUyX7zN0UXDdRKPf7P/FcYsVVh1IJY
6lMZJKy7d/6ViVSjKtLZgGWgAelvlTSFdnOTpJ4035d275TIWKDgWvfcHGYxxu5P
d0Exh79EztYxGFmgJZSA+w1vwUGRgR8AAhMy75JPhzpM84OoLUFXyq/dK76jSJcG
afLcbqY1AAHKm7WOYnG7bV0KcY+bxxbGAxEOkoqDgVrohPLq4t/Ez27wHH9d+v+E
Ab6qZxSh8FxLHDNYJ191JL9868r9YgS7bSJWEpxbRFFzgWV/QlojI4GhoxIN34zV
9rNCh4DWFm0vBOhLmdsR/hK1h+rxdx7VE45XKHAOyViAzKvKsgbo5aCT4JTu5+wJ
svcD0s7Y5pHqX9M2CbtmPMtOKdjKOicgqT1TYCvC1PjgEuIYq2ACR0SBLqMNx3o2
s3hw+8r1zR2moabL58wlsmvarkrDdg8XMlcLNfjYUEvrnUeTZedBIx5ksxkfMnul
OiwnPLaD19JsCRHjiZrTYEpQlJd0bnV5xZh6nrmPQayYg8bG6+6nuZafcY3nWgy3
R4+airJRXLMBB8xhSRW8mv6rt5q2OGkoHgpfhMPHixmnEvzKMfPgxXGqwXvVwJPR
F9FeizsrrCbjCa+Sr6fDEVa+AlmYX2v34W5XujYEsAh2dptXDA+z3k056e2cpyob
hV2kwByQl/+SbTVy/ErWLdp1d4BitR9vRZMQLW1cwYXU0qXr1++e1efYg1ILCxlu
TVOUbstyG+V5kpUDjLAobRW9LGxteB96/zGo/UqQNDcaKex0sABa/MzRL/HMwMMA
q6DPCXt/SL+XwHGB1aMqawMf35CZ2W4dt37zFDuEs7SjUsPXiv5sCth7uVL1DjGL
xKgVxPQP9exHzoEFPKRf4DK+FxMdoMmMQNH4PVDxsP4wnHRD+muUZ/AX5ZZpcLBj
0DfOdI4uQ02yOp2QwoVwnR78RqBWKhVKzmIM9+yWPAb9KjOAUw/ShKFmwtNcQGXe
vf5kuTBrPyTEo38n8QWsdbh4yo6zVWNf1mgfRWbU0UhxPltL7qR6xN374Da1G9jN
U377bCRoMPg/jmQFXyPxWXpqbwPkZoosnQ/EF+8WylcWkYCl5Ja6087T+U3/oi/y
UjMrmIdnHB5AZs+kRkdrvlSxaJyHQaJWK7OhLSDBdPsMtZQyGsyFSXLSGGE8RNLP
EXYJB8peTPUnpcYUzo4HFVEsceiUHGdBf48JJ7DzIigEnh/u2p/IfdJcoYLtneEJ
RzTOjZOKlbSesPsuvLwYZt7ofnxW4n7lTEX4RdJxkMwgO+yaFfsHR1O2yjle1M//
2Z8YQo09KlOgo/P3igyk7iW6MnVMIOAa/BQvh17dcjUPN5288Ol/EeHe4mppVpvz
P+i8I19oc59BTXQi1T8AZ1IdAhEo8zw2pKLA7thiyOJV81Mz0VTIzjaQYWIiUshG
Oh2tOCPWt6cLtgldjuKERPHMb15llfVV/W2yoENjycscBaXaCTAshByUA2Hxu3Af
Y0faqUFsm0VQfO2oaHUgW6R8LPBVyFxhoed5Iw9n8V1U6475b75G+Zq51auaYWqK
sd9ttIGieZiP46KmC9EUEc93x1CmKNbPSfiOUrolO4388SmKHvubctcvKvaEoQVa
v4NCpQAKvupAFl86PClMSH1gqR8pLceAvzzlj5ejb8gP0M498NkHQUF3GunCADy1
EwZFnBLq95hy7gUjWMcLk5bwN9l4FzTsQJ6oyUt+FhW5Oh4XVaBXpC8aW2H+Fwv2
ce6omynCcORzk9YUprFquRWRJiZWYff5UjpT1YV42csK+jscfZTB2uAin9CnPzzQ
kTQw297sg11q6lifQoJNSaXR4JlHxyMHVYMP9Xdyu5Axa/AUtvqGVSzoERYpBxn9
1qr8B68XmCkM513kSpDn4XklmHiMbbKe7kGUDKU+qaZMElSaiO38/uxvj39z7Pt5
oFnWJiniP4MmaLztJ74LcTvWfF53NlVO2wvS85wdRRW1GakriAubQiHvhQYHpw4R
xqdq6a0t5qZh/b8TOaPINlDp97ZrWkoptbDnwKeYbeQwicse8xMU6eM+tkClWVtP
rBjtFZr/f2DWsNpfi2mGnwQDw/1+lhTQ0upxLIstv9wLo3Km1uQX/DvKWn+y8hsZ
soaeQ4TA8v/9Ll7v/IFWGvY0zWd3L1oLr1ldmGA/61HwcPP8t5krQWHAU42lSc+7
imZ0bUjK0TWYOYLTOg9A4w+0XjF7XeNA4lGn45ZCzYvOhQ1RATc7pslCuFQZycVs
eo6T3Hbjv+z0E0UDf9nyHakGTEK9dHU3MffdHfKgzBb3YyXMsVFF2lkZgZO14rNk
kN9tpRk5AY1nmUFS/n/xe4A2CYuC8oMFiLqEqk0fGLOU/fl2H4BuGQ4HT95pTgyg
elBM1d+dX6LzHvzuk5atOtFH8v9sWivocRw2Sh1Eb/By47d0et/qll4X8VDeCySL
rECEn1SXw7nlVVk2lI95iAc8H26XAbjb5cHBRv4+1ytgHNV6lxGmroTGMNHT064w
LL1JIiHLRuF/4TVu1ezxXGOhJsngDyFvsbrsF9HcHs1qejb4nkraXIJk9+0UGMdW
pZf00JftvG4n6J8WYYlb2DaPOPcex7QDfk29iRIB5Gz3D6XAuztFSJvboEOut170
pIWVjMHZ3ONZF+BojR5wZe8rkxD4naZZxW51xZQo3c9W7oNClL00IuYtn2i4ZBSP
giOI+V2Fm1HCKp88T8BG3VsDTnw3xT4CHR0X8LPsDC4M9bwd1t5jmNKNVRCeSRJ5
qvHDNlipn32gOl+KuWf56XhS2NmOglKZMkLskhjMTXdCDQj0vpCSQDRnlnmh5QmT
Gqf7EySVSstPo6tUr/zDsQFQHD8y9kdVO7z4GTHn1DN+Qvzuv7RUcphxKlFcbaiQ
14sJtF9kOPxV+/CBuZzmLBoilrNVjKRiZIysRP/PU6kO17RPXnDE05WnublNepSa
8lTL9hqQ2F3pBXby/Lxf65iqQrWafI/jbYCkq5Kg11vujjIXjzy5ZENK7hArsMmp
99EAY9b/X+G26Sb+Og2ERbCx9iu2LgL3iwYHrs+1PBJRaGTqFlaI/p40KmcdRH/f
EHgXiA7HUvyjTtTTKMYKBn//XFb7i1VDnKQTZ/PsFLS8HczNWewpZGPcHDVqo5ix
MA5UWuT+RUctcZmCCUpWkqHUwrU9kn8GIIt8uuB8SoxdofpgQpTlET1l6TR3Ii+i
NP61YMhmVjjC3K/i4w3BBQ090gayUA9wkPVfB+kPnQ1cSpSes/QfFPZfE+7vw8pW
Rt+P4loE6HvcD1wic1qtCZGkuoQbWERzYwBxrr3YnpDtdu7Bln19+cKyg7aotdIO
68cANv5ktSMPi/5K0L7QcxcNRoPwv4O7ROluYHx5r+PXrlGUYNn99wYKUvdMVkYo
0s0PomISilbA+gHAMFLP3ulX34V1whENWL+7ndoWqrFRI2ZRPPISYoLwfGYQIhtb
QHABXeqObqJqsI9xdkdS3bPXzBU+38NZ/+fpNJtsD3gCjO75mFV1iZdj88QV6hRp
PNsKxECt0JOKxCwHRKj2H6hUkv8cPddT+G6mkbHxMTksMyeqOcIiHKGbyNSH+4xS
GnBDNGvBN1DrgqlNfqap3JjMZ6cyjXRIsFnCUALy7oeUpmpheYMsAqcLwH4B98b1
cwHJue4fkEKRnhQ2atEeIpf9wmKgh5SPNSfQynAcbEx7/EwlfgyAhD9uzZpcttmb
e5ut29lCkvrWbuXqWt9sKtzE4TaSbCBvF/y1VsPvSngJP+tkvfoVMf6HfGk1LIge
UjlbVN8kIHQeJYKQdtIC571/B+wX/jBTCGRESK3zXpTOGcMCDN3J7cO0cLCAK3K/
B3PxejcYasqWoz/cnbZr7BJOuUArhZcDdoZb3YYlLoqndYjCExfvYkE7PnSpUBJ1
bopm7m0hr66E45lzm5LsL4eHwdIUE8q983wb1FpFl1wi7JnBaK2uNpyKVIuWIMvP
UgwSsMKC8hxzonxH/AMzJQEXnwtNZkEdHrAIkry4BwR1sNCk0RqJhWoPSSSsilMB
4HCohnIKbOGlKhP6q/ArpSk2Vi7lPFG5h/w3q7YYIOyya73Ha0PDkkvSV/JVB6SJ
Lm31l4xcCocF87jq2/fo0+CBu9z6U/MPQdy4qF4n8pSiEWcBoLD3G3B/oIvI+P1Z
DWoIjc3urXOFZbZijgOSnx19gw/vwPr2lyvNRZSJDMAN7MhBFuYLvaxz8ZNkhU88
WrR4JObco3US1yIPPKTANdbzqSWEXno8jy6Pk3fLt+x4CTPQWVKzoUmUMAihy8KI
IhgJ1d1dlthlcQp69he4EAA3aivMAnpZHMHwNacXQ1gHuMzYEprqrGzgS5dYl+Qt
QxKI5zpjo/Q6qzu1WxNminPcgu32kFNEmgUEW9eIAhPnQVGcTuJYU6FQmuBCQZ87
qjbg2ZokoJWQr4lcCgT86YGdFJBO5vkK65k60QscUZtId3xuvkSS5shjAFXpMvDz
zhCtH9quFGp9yC8aStpsZ9siPTcL9HjxkgQGoCxdv5GsZL4A2oZeSzdyiy42/ujB
xFf3/504g47C4/6VmEmhG/vD6n718U6KnzAvXOANINjJRRo3X6vp0UhhZOVmxCkj
8Yi59PQ9amBi7XRL4CGuYJrbfOcc7Au6AOO8mSdC+OAUU/FztyLHi/hnSA79L2k2
E3cjT5dIP0mTiuaXOQgpvxeufiNM9BZDzXhRBDFjFoWj6zE2MipX8r0JN+O/15vl
jKZzhhgyKQjHYpiJqjXuF5ymzsX+YR/0+ZLqbRfils5XfcY0AJ3eyO9KoMtXjn31
OmDIWY/Nkh5UnlxiSl2vbFiB5ZDtqwp78sV8VX/STy0Jqz82UEeJnfBhotheVaGH
jmxe9QHMX7z+Er5gEkHxK/zkEzKHi2f+OCp5ZBVG5sAM1uQ9AcX9WNOiY+1z0lqn
+tOw2JM15O3x6eJIexn14XsGPLn3TwELC69eCSyy1HVUfFrZ1DYOrjj9ymv6qdVA
54MRJI1RYA2ag/rVFfQFNQC3HgpFcKSYE1nih/au3kfCrhCjrPS/em1w48S3++Cg
gfOZUFe3hvSXjdgEqgJL/NIqs08o69t+PiKD4S420DHDgI3q0UomBR0z1mJbl5tL
i2JkWSyK2Mw+VeWWYzSPOZLGWThB5SlZmBCU73UWrIkCkjo300ke8VXd3acJ+R1M
SjAJ5Dox8euBhd36JXlXY9dHsUW3YtukxWf3cDrZhWGP5olq3+RcP01lVnhMASCx
8l04Um2LO5zHdLFoMpYoyweEZOE6vEypXIK3QMfqbSebO7Fn/d3eiYrp3e41VXnu
LqxxJGapwsmHp27DlGcxNGVAJ1j+grDBIIRgKu7fR0S/etZrtZ0i6ICqe6UzJARW
eL+6F9gyRl/s21NdD7EaREwTLiy2GTzuRavsMOhc7jJCjI0VBqRVR8zL9QgtvgQt
CZyW2ytjtQidFj+NYEBesMQfGN7ij6gNvZu7yJu0PbXZ6EafY2+sY5YdN8gPDgW/
CjUmDMsZlxwMT+xE0QZPRtqukYSYIJY4mrbxJbgK3vUmDFZGf7Kb2CgF8iIGmNI2
VCJrGBgSoUoLBekwqS7mfuA5QvAjK81Q0tFEEyWEaoBFFJYQGpTuv5m3GaIJ6BIk
z5NRq/maF4vnAEJIqaw/dx4X9UeQ8iSqAWGHSnzOC36152BecdFb5fp9hTY1bKMB
hTHlSUk9PdZALp2s4cffxMhQnSL4W66XqfGor9GrLIH8a9ZkH1ov+ox9S4WWz1ix
gKPmX1BMchEDY/nC6gcL2zBFRgo2/JVh3K0PxyFXUrjvuYnZS4fDzrIOsQhvMMoa
zIYK0DutNpkbT+xJ4qV8keemOQt/KQhGEfgMXIG6nTtB6rbd7hgGBAxMUVUzNIxZ
NmPgLrlzNudUtFERQVE5+uLTWf45EPPq2xI4Gaean0nD3rLzOiRI/lh3AFTK4EXk
8C42TdxJE00J9YX6qAw4VR3qYY9emBjyw39vbER9NE7k/XKyiRrp585RFV3Wq4rq
GB1iM2P9KswX5CaGE8wnkkuDjocjPMoy+Z+f6R+TlN0UcR7FZtGZd5B6yLeu7hEP
LMG9GrbUe3WpfEYU8eZpU9oHCNyQqq7ElLTdj0jNJk5DBqWLj+1hewtwVFJDKR3c
h378XJmWSGVXQ5X9IcEHw2oRMxJM1FWpcj+uT+qUfJnq3uVyyBwuNvPc2OlfTtVG
dNr6uYEB8LO5qSbJYryVaCLIEpofGT3yYMdJTS7BlZzMby8HfDYQIFlH8ReGlttc
It24lNgsNCW0D39A1eVINwzWqGsQ5SJzByMDZcs17WIDRtoteKLJRao4D0vmUvsp
yThmE8NOlmeS62J8lqG9otTQWTofSg1q+gmkPH3RarLNZT5MpsWU080wfSiXqz3q
waB6qtXf5ASOpif2G5oKuxaKm2PzcPJUJWlTnsYN9LUd7SRFJXFMlOzmMXYv63Xw
axEkUp8yiEJ37EW9xpAYfhJnuCYW20we1/f6+/YFokG1+D2Cse1jR3fEFRMW8ckb
7uzcJ3x1hlVPsq1ENuKNsJgt9IRGDxCeWAuU/lGi76bc9oQw/5sZbiJDe9g1oeo0
s095Qf23+P3Mrqs9zKhC+dd9B+P9+XRyCovL/n7SvXXjp01ZOb6+UI+XV+IwQjHK
iWRjAgo6WCh6DM+3kNm7Czg37VqB0pGJSTZRLbab/ZNI6KKdDWG3xsXdkwGEpuN8
Sbt2dknLV0vyynxGCThOzL3JT2NAfyc05u+3GDxPkfCce9djcN3AErOXDPwVvxRE
eHXrRQ/1/je14ual78gvXJmaG7fJxnnLZJQpjxogArd1mxzDbM5M2D5R1sfyX/is
jXfZmiT7WJI1IYLOanjfDzjwzuIvkGTmyN4n/zGgyoOPlDexYXTeM7sqzUZjK9Tz
BqVs5Ulav27bQfeMSaYXF2+mqdfbu/iTjW9TR4z/2bJj+yH8WeulNra/KIbHZ4CH
CIruAgWILAb0WrTqBl9ZfD/WTWB2GNGeIiFtHAq90OFOUbnShRpdnROTPYJS8m5T
xDPtLaaWrrd9W8L1gUCtVogvliM+cinKmqueIFcZc2k8n9uX7HoDSAU1DIr2uegL
DJO/qXkbJkWdF32ptEA9gLybOUIo7wo72WGuTpmD8Sxu9AK9dWiuBsz4r+qmk3yN
d2UtE1svMInau7AmXMGV4Yjj1ONRMJ9dF/47wGTJGsdIPUSbSIshpY+hi9QsARgA
Wx9bPc2bKkJCHEcbvUW3MD56HIqT0TEDA5pPn87UQkdMkrBXAbBsbyWUfA5NzaUU
2TCooeGzIAgwoVB8NF3noIjkQjK4+rgQdoAa4CNtODfD+VWKd0rC7PsnGhq1sFK9
8iYy2dtoyNI8X8W5LWNdGdRmz/TCC8cdOsTMT4Y02B69Qm8ah4EuKUkGF34orOy9
LiirVqd3Lz465up+7C59cOs/9SQ/h1JM9OGQLs6SzJb8djlFJ6+flnmIPoIhRx8q
0oaMyoW1euG1pHGKq/0BiD0cG/HCIPb3WlMegYB/u4nRWSaFJtSKwktKuF4Ds6Ns
7d94Hh//HwRnWdpx/o/mKBS6JbobVZ86m9vTtHCGAMywHb///5ZIHufoLr67/cTj
lwVJ1yA8X7sETLcA458OfcHmymVel19oG2cz0H2hMCjkT1yjgcpxJHdz0OEqpLpS
t716f07C3m7OTXoWQNeqMcM7TNvcdzWRbkyiFcJLAl0=
`pragma protect end_protected
