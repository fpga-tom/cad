// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:50 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
B004W5i11Nlwg12pJz6t4IybWzq33fWD3XMFsjnuEC8fOY2AI1Wlu3yHZ0PZBxeD
3i2iLY7ZpdF4LBEESC2sShJsxv49VsDNRk0haC2fm+uIzO0v2Z2dimqgpBhWIGxj
zUGCioA6a/K6RH3y8rQOGSnIiRLNBcARO7NNaecsKD8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3792)
eW0U1D60aZicJPnFd7nuDBkO38Ohxbos54dNSA96yTZW7wxZ9iwBXU1y+wgnxyTK
SXdMLABb9NhMwaMrVH2TOElMvMJDLM4vzD0D3dOHt7gQ5FadBiTm2Rx5Easmth4Y
hJRepWq3Iw5idr2kKEXjm9+8igunMLL62H4rzJcDjoir2i+OHPxtz9dH7VZE6Ad+
doDDRKU6A25iyyuZ4UtbwyRiHRIIT0I9K8YHz41Sv9DPPRizfp6GT5iYXg+Alu/6
VyG2PyyIMkf4fSXt7IG18UKZQDuyGf5kkkJBW0F7ygkXvlEc9iR7ePtQgk6X5lhF
HO/82b+nrsFk7nyLM+1hcOBQifrFLmJIjlDMRvaPen/OopvVSEAwHPfbYe0dwpjX
6KVVGvhG7l9u8J7BWGLAlXHV1PhhAc/fXT3lA0O8bNotasjgFFjNg+lGonM2jl4t
QJ/CL1Ur9CkXMX1CSK/cTJd5Z2+ClbY3zFRwQ4x9QgITZZn/8Cxgo8r2J9TN4VhT
CkNZve3hlEe1fz8wBo3WCOXyT7PmPccM29NFnzgtech9J+CExP+5vY40/HQE+GZl
IygraA7rzzw8NNWFV4bdHsNekEuewTXQgjr5alGnqQBCBWbsONpX+ySgd6aPSduG
+Ffgubj2RugL1ic5zPUe0qrCZI7y01mu3QUO5lpRJTRj2FgQklF/pKUwKYNUa0bn
zovqpvoJyXvCG+U9NsqmWNk02TPxFusPpzKf9DdEbmrluXHfuToSEmyc2QQFSDvZ
nizFZgYofAFaSWl4o7wY8+41qsxFQAb4MiRZRlBmT0tEJREbdOwKLoLsGnzBioM6
zL7scZem9T8QN2JJA7kFrT8OsPA+ME9e3HxQ7deEoP3rBiPFLUy6/2EMuvjCFyn1
+KclVsREca7atdoaTi9bc0rKIbDQylIfa2cJ1daYK1ZIBBXCJ5X07+0Fg1LV4s4u
QDGOxIJBwsh+w88a0qphXLgQAbLXCvI7MGFo4SUgA17q3dOkNUGId5sKcfOSJ1Gd
JvdGpkyo/yR4nyd/3vI7bHDvOPcDjN7RK2qFMb1Z6q349njL1MXRvREJzN2KlYMU
Dd1ZUI5fost5+U8j/mJrQ+MEqKfwJwLUpyOiLKB9t8EGaO5AP0lcWbWpGtVuYhYc
jGZaDgQBum347swKUTe3Dwt9EAn0KFzN7cLOvKZtwbjgwKwekTpxBZeriAOwCr4w
nPl2749WqgJ345WyDznVwivbzGCDS23eLz+xppaxNwE7ytYhtSjPCi9fT1mRBB+t
7x47zgjuWDSJncKgNOc3LirTArLnOIIJie95l1v8A2qC2pLlqJH7xCSCAYBB/zOc
KaBg+bPC/PmnVWxKQLhyjCQbqTvBkW9CPD/FMuCHJ8HYQ2AY/pN/am1Qkw4QdGYu
Dp+Oqs4fk1BBr7QFRYz3gGCt/73UQAWBh+W5YNK/ebXsUH2z2j134L1qhmqNIhW1
HAWfJXORSJfbXLO4dtrVDVCjwRCKd5pETg+uZwIT4a4IRkEtNNXumhdFhpOjPnPL
crUCAqgKwZPNFie4B3UaigOUe33Y3VteDo6OHrldLyRpqWk8sw2V/N2SLu0IFffB
twamZmpXaUW10mXhDkz6UDHjegYAS9Ez2hDlF3tn3kUCIcxuEpY8zfI6rAhE9JbB
mmxXvLbUXAObHmrUa7FdKrZOvxPb56pAn20kpG1LSMnS3E5CIgkIJ+PUz1GoNI9J
z28vFqsKWLqiHFQs1KipzhK2l8ZB/j0Tlyqe4Is7/+4WPmUluB7DwAugzOFr03Qc
okg912a1nIcjyf7f9rg0mzRSpAR0VJkgcSokXTa4A8bJo0IeCm6RImDuOgkCKwr6
ufXCoULIVmLSL4Bv06DR7pmAzT7/K31sth0wzfxPTVUBArLoUAQo5wVQqUeJqmVc
IgpSqELopNGbSbT4sIPZ5amBmmFft+dX/f7oc/7AgKlSnCJIVA/0ev0zglfsWVBO
RGQVNnkn5aPj7CKtKCeqkt3Z5+RRj7NISO5FXFcya5oQTFVks8+WbjxINK975eRT
Qz8DL+8NfjsRGFz1witGVDApv6auULG/4OfNc4W+er3agceP8728U9F/+AwW3qoG
DzKc1uX3qT+4HcQ05hHzRtX/pyKlzWGWNy1porGatQ6xpFmh3Jly7cjPDA6ooLYp
gW/szsZCUuCLb6xepe6boNTXnFg3a7ZhK9UdQa73sFqxABTYL+mloPyXVpxXEmz/
mb7aU64sVXpegFgU1BtQr+z49AmV8RiFlRxGOaFsfiWpTayvUkwWMXd2iG7PrZYE
g7TnvVQRspE3I8QADGxQfmrY0K1fwW0InRSzMI69xns/ipEgn8KjULuXpk0h3Auk
E7ZmnRUuhKYaUxrRoMIbfC90cMqQNjQ8qMecWy26ApDZOHJtsZggxlRLgYRrG34u
fI4lEQjhftXx8A58jG+xQxVwl7gFRvJKtova1RWbJL+Q9tJZZPHNMXvivK3BFRDg
BqHG3DxXHY8JMsaJDmtliD1331RWHE7/Y6f/gRv9tth6cPhmYRXAwCe/QV4FLhMh
pE1USy/xpKLHkErHpY4C4ojLF2IFy8oo8t9ZR6dnj2YnK6Rv2Gg/auVyKU+Ml/IK
+9ZemxtqiDipIKD/ds7Pzgq8s2KG/cm4TwbQJEsi3lcO6xZfDvAwzPVJ3vzuq0kb
IldKLw5cFMcqRFFUbe4XY+pwBKeV4L4Zky1wFEnaKFSIjEEHRUr3uJ9BgNcIaNXo
8W7OA575aoN/u+fneHhiwwzsJTXAIx/1PETcNBEKTywgykZd3bG2qk1oiUMtPP5H
DKeI1vfDYPvky0DSW8BUGW5pVeTZGiYrpwAoSEtaGvLh3QaNOkIiMIkrFR78PJeq
JtpC2EV1tVPkArFuk/0IitQEVwfMWSaJ6am/3N508/IEPuMZQjtk9xUBBCSOy3i+
2xochCMQ6nCiFkUd4BlY5QugcBJwYxKRwHPwgq9RuF7O5QOfCpVP2/mpvJNBRDcA
DsZ93vDxeldYFkPkpkut5Hr7SCTA/uFP5GFdrIPpWLKgNaPaXWc6YF37cWnplK94
tVzVzxBcpIu1FJLTBsVpUtVB0MVt6dPfbs++p8rNflObSyKZBvSYTgSsQg38Vkoi
48FxJMg4qGuql1OVNF02ozyzKcltxsj12F9JZSog+reC5S7lYwBejJMdjUnkZqld
qg+jYRGTystuu9RNWE3xPG+lsJJ/wYOgPfpKQY6mt+w9vBlEd9/nJf9oGwJhJZ26
Z3V4A+7y0EcTOJWwEwr8FgGn6mzQR7nM80HnMxahFVpDmtASJaDdwxX5mHasbW6j
YAJkCrCosXy4/7GvkUDPl3h4ygSkDUhvuQLF25AjozPT0yEFKcir34B3Vy0fFn43
SyGtn4+hLUzMp6Zl4h8i3d/84z7o3XKe4mD1o+QfLM5nfcd2EVWjDCrK337/Hi/S
KpvL38sn4DOa371Y4K8/oPwkLxPuLT+HvNja7YAHjEbVXAv2NJwvoX11d+jqvX5/
628rMQ9AKe9mRaUhy2k9D+x+c0fXg1OuibC79JaV9GMLaUiruoIfPeUlBjeaOVSy
yb/J7KVpGjBcXJGHiqYA+KKE0I5d9S61GttCY6wz8H2stfIhx+rQT2y3t9WjK7uo
pw4XwHaryuWkCnCzqGThMGfoqwxJP0UiBpJhidt813/QS+qN2u8NhfsZ3cktF0eD
KnOrJWPkuhpgSJnfnhva8MViIvdy/V83CnnGC+FfwxKo3qf/Yd6R9neOZiJVqtja
xOoO01MZwwmw3LiOuxwhue5g5I4KBepm5lnqD2mpznQUHv0LPQsEf6niDEhiZTUW
wcsVNl9yKPLoiHjblsjsyqtCNe40RJf63e/eva6RHZqh48vNFVuxYwouuVceN92x
M8G6r3bffLbMJ2z3gYlEe8bivG7ArkIsKyLaSzyUVa7AjgMesOpPBeMEyJV7wLVi
qPmjqNiqbuGRhlBZaxaJG7i0X8ct5Xq6WF1Ta6FBsfxX56oJwtarFeoXngDHfMG9
deJO0AvxUNBq6qN/2igSXGEXMYfaVsTvdfsM4bNEijBfh59l6m/J1201Xi3Yltfo
BLkzlBzpNdPt62vPGryK5UmKWrBhVjVoTR2ypJLN9IwVjM/RJPl1sHIPqvsC9DLY
B4AQtuZ4wvWr0mREMRxa2ypfutrsbel5FQeHczjzyG0Rkbq0b9jOJgjZayqzuQ3i
gk16gIf6uEpSj6YQefHmqKULV5trpIQTZCM4b9zqU4+FyZGE0KLbXXSU6nRRyJfE
AoHuwdkTO9BGSAdohAP8ztbl5XXC3R2JmzmSeDUiLazoO1LPRcX2ldkBxP95QUee
payLxv0SgQfCuM+j/RWt4UTpWT2bT44rwc/K74dsUA0sVmIENaCfnZwBd0UU8RvO
IEfGNvE/gKe5N726P/3iCK5oPy5n/Hy1zCSwwYAJ5Fa+ITcB8hI+gVy4mkcL9Hha
4JErcTXMuAtnCgsTQocOdV2gV7YbJHzRo/0j3btqa4lQp/ik4vsZd5L3OtH2KsmO
i2bJpKrR5FKSU0PfTgOREwGlyyO2MxWSjXR5zw1KhLmWUyZk8KOmGvBL7/ipxZCo
SbXZnfMTrO+tgWLBggMoRXT9z2U9sH6NLHNvN9mNq+Wf5KeHNmEUcZLGZKnyt9ez
Rbynh+44vAzN8MRewGrKLh1xpNSl7r/ByJcMFDLUB2qguSJuAJ8ipimCMk+UdfcP
BeZWzaOw0D9bZX8MfQ7MB3sebaD/LHVpQU8n12C+NDrS2E9aCr+yq65uTWp/3MGr
HpPuOwsLUHlJ7klLPIhmVVRv+ZikuSIOu7BFuB+ONNUEqA4D5H4QZpoH18FoLD7l
Aju6J8MSv8WJIqVP/11RYajkeI2L2Ugjw7ZD4fJHK1OcC3o7tyUCcasXqpOVmkCq
WB4v4V33vVKzsyPSSoTcaT76zMxVJoEgDHmG1XMZE8Dsf6e4+bJQud5Qdmu5AN0J
4FxZrEcOUklZhY89kNrAsLFproi69ox2ecmvwbekU0n0u8svykq71qwkGfCFmO/Q
`pragma protect end_protected
