// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:45 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kLX8XZ6UBAUU5BIs8JqE+1thLKp4e8qG5GmqWnSOd6Iht/biOYURQ2WQKtVHHAa4
lE7cdgJi8yTJWIkw9ml5fofT699wPh8VhaZCGwFmt9CY6uaoX979rwOGNJrAO43d
Bsp2CB1swQaDdtdOLCFvEgzNcbgtl9AtPrd3Pvsmeto=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3520)
4Kq0eoRBjkBD4xagZgyxuT/r8ixn1js178C3M/oQBr23pN2l+DDL+d6SIKWMQiQN
TK2dMYJPthbLLEkNRE3DPGlC4gZSs/FfNm5FPjV6ft2Yx5HG+sWsVG554FZbip6u
193qMdxnNWuTrZqf9yTImL88eXkMmc8hB1LmFZqJnx0Us8x+2Fb9aEqxCCZ5ldDg
+Lc9nK/nrEyZUO8QFtvHarX1iwHwg/YpPGxzzThRrcxw0V4wPehJhcwX+GuFNmPS
DQbIjzklc9bWFCFIcpxU3pj2OUtXqv9korQBpFVMxIzktp3siKXJ2MMK2Wa+GCmy
LBKfYEFaYrFd+Vh0XjZOSpn6TmPrsfJRDDiz5M/v6TlF2wj4CTA4zojrnjdgagEJ
/0UvMmjT+/pPqURfJ5PBa6Owgznd8MmtrvU7kvkXmZdro6mcpBAp4a4XRHabejII
ywiLP3XcCwAbG4Sq7nxnikOOF4nx9ANErZAVQhyw5ylBtm5SwnaPKT44Uefk2Pq/
oBEzf4ZwgYmexK/RgjppKBH/a4pGP/SOrFPiJJY42+0TA6pYouyQ/t8BQmqiECB3
5/ACvyi4yx3oL42e668TKrd8Hp7/TDD2l6gzGeGBofb5gOfRw9XUmKt+kS3Knkgl
Dy+TeFY7b5XIMt3jWtVJe6tixBtYXHklUt1iK7iKFAlJXbml0O4qvZR6BT6PDm64
OpJ3fbv90c1t5XgWwOSuulb41gVrxz2wq5cUGAxwionEcPF0E54qRkAHvNKzCtOF
RL0QKnma38IaOz+n5guPhl5iLsqJdeeg1js2ATWt0HVB9ch0HWq587qWwLNfsSpu
JW38ed27kYihLOtDpMkYogfH3GRhRxe+ENpxvQbljMyVWj/AR6vajgI+h14H4woY
88YKaP/QlYwSNcmT8xsBZQJy8ExiGeutlL18+xn2LX6+Jq+jrrsklz8IQgDDsEdy
d6JK2zYAOELFmrlxYuOcasWyhjmi55NAaMkFHyefSwPooVnPyM7F+IK8BSIJI3+z
Q92hOnrxVt1/K/T3PGwqgkhq+zqycesHuaq+K8anuDdQYXDUnsCuvhdng+JOCyxq
6107YRFpcikcTLT6RRA3izMnq0sPX2T0V77ARTNq7laETp7VK4gQKTtDghZZAV+6
NuVPzJ8YjxNiErV7TLX4m+ELHnxsb6H68DPN8W0RfvoddSunjHUdOfEhbvewq1mZ
bz+VTbjOHQcfk6+APKpvxNg2jh7dEZ1XBL+VX1rbLxoR+CSRyZoQu6qO82wxgd7v
uQ32Xo+OT6A0Xol7Q3omD3yQZz4qmnfWYyenMtj/waztN4nJf/5TbtB/PR8EEosx
3ArrpUaocvhugsxW981KV7aJ1lgmoykzTi+5FhCkWGuwRDXZxnpYANBtgdTiUiPu
rkYAKK9GTWqW/aG9by5lk8fmdRllawSrRHSr9e6U1MvUxRtXdrXDzl/XasUT6hpF
R4BQYTB3wUuHGy0lTYs3HYsgSuDe3TMLy5qSIAIgeAWfVSFniRUANyWSskHpunoY
kIF9QOELgY80XGmB/XsgpvwRCSdBlLXVoFPUqGcWtMXzVLO9NH2vM7eTKBDivoPE
9EtkNDX7s9VYr2lBMrI7sxnHTj2uMJAzbbMZw3dEuNiFPSmQ3H7yuzflszn35Ppz
Ad7+AMtGtZne48FyJINe/AMyjonMxLOAuALGdXFD6A6Jj6BsgX43ooZaGGN9B92h
SxFqisjdH/94JWVqtDuUBoEFUPkeY2enw31P64jXZb8NOydDv5SBY4BD2nlihniP
a4jxOshuvw4OM6KnHbuvfOtJAXWYSaeFr8XAeiFck/gcFhYbMN7LRRfIsfkQlpI6
Qecj0zxLFJ/Q4CWMyKLSgD9EuhEQVFzmhjjqNEA311cTg7ArH7yyEBWqe8g+A9km
909khp9Ltk9tnYAol0oQKTBgXUpsZe0E4WG2FqJqeyl2BiZwUh0ce3+I0ejQ+xX4
hZuQ3dBVnuhEQkbKj98LkTrv7OcCrMU4NU6e4AY/VW6pRo5IWmFpZvC0gc1pqUEp
PmSaViopXl3gWgQvCdoS+3cSq+dV8VMlj0+v1gluiqj6nfMBN/CldhYvmHzACYr/
cIGfKfc1nSPXC65v4jtCfQdwkwRv3KNky9GKqva/o54sIIgJIctk1zQcHRbtOWgN
arwFqIVdclmzeKUKkFllAmydCslAGq7M5UKGdT21Zi8ysm/3vAFhQ26P6dGZUPm2
vExQSe0WhxWgbMoB6yh8lf+v7W9oZjnhIgBdabr0JPbFHNSS2lep1uvLHqPGEyYq
IF6hGpf3R60s+fIxq7BCyyrRg8SeHOlNvVTCbbuQDjFm/M/lVO9cA8y0LGOyrpFs
LSgkHEfyPFL11VOlYKiuzbeH8fk4uti6yFIDwtD7E4EQYTw+fCmUJ3Nb/YhtFNTH
/n5k3o0Y7Z/NmsIDao2KzLcgKgZqiXYO9GADd2yhAGz0zt9J0zPoyOO73Ch26t9M
0UI92HLkE4ZlesxTmQipoW10XrDjVIYtAymX84CL7hOm36insgTypK3B1Ul68JUq
Eo+zarvJmbs+Dq8DMbGEVtY6vLw7vJPQEVLW0kY9OqiYTjRiNHFc5ztgBbNpOeRf
rVLriFZhPHgbRfrbZvBeU2S/0JX8bAWpzBs4zat6pKrXV5D7FDmkapxhDlHtCJ5D
03kl/o9U72/bSFnOs9jps9W93o2g+p/6tn6U9kwH0FCfG3wLrnZea3aAQRUaoXH2
S6mfZ7pGoLVCSoN5w09yEjLUluCRXiUwuIhwPIGkghsuLZxh1LQOjjnLY4PE4Evf
r9hF+hcHKCMNLIZaEFekbun3oGp8iqB0A32CIl5N5nCwuSeBGvzk8p20IyhEjfUM
R3Gv4umecT71cuEPnUB76zWjZqlqzhtcke2mn4C+GyLgi5jmumuTtyuYnXY7LAWr
X04zGRjWhbtB+45Xm/bg6eN4byB8MIPAupdAA43aRfZ/I84fh6vzMZQKIAV3Ovjd
mqN50whK0LpnRzbC1MVQaE4RExxaNg795t4E/tucApqoOhw6wwK5YqIrge1G3vgJ
p25W9k5iLz/z+YAhadkJCpRMJWSHS7F/x484rGUxE4jm7ew8IrGvw/UQ+68f1uIt
hnSZX5vDtpjPJMqBu+NM8wwLUUogPaJNYg/G9jgqaQFd9gj/Jx0sBsyDiCROd4uK
DMAWUSYceOgA18MyxUxoYitSuwuvuF13b6jA6X+wu5uptuoK7ToUPAGAuDbtHbv6
MyKxNGGZX7SUNjvX53fGwpMLhqx9QoORiPYWCdSdtiFmRhHZuexitNT9AMYIUkRd
jBjz3JYNeP1bOLDwqnixZiIiAaHYDlg7n1zGfH4B9WvEZZcNtPJFppsA8Xzn2xXv
NarvB4UXrNu6WyzGSzJpCGBRjyfjWmK0cQaakpbCzn+hzIHPHbBJfin9cgK5eVwZ
Myl5JXfY0SC3OoyO8fxJGlA4PLMXB5DMsLnrl/pcID5NQvK3gYl78Hko5x0PJPZF
f77gAepkdvKuVDNujC5nl1SjFC2c/EdGBiBBxat5mk0YnpTTU0YAttDD4D8x6/Yx
QfD9zMrVRDE3WSussLbSIvwKsUfEgRZ0+UJCTJJ7Bk7eP3yVWyAORANcwfJRl7mH
md8ZcLVZLAooaQsZaZm8ouoXgIRXxGVaKlTEQTPth++lQmJ1rZYSPJ8UaMIxC5RR
WYRnnvsIxgF0uGAG1OSe5GhOiM/M0TfGzBDUi30P3CmwNaYwDtkXmvCFdxO6Ae1E
1W/pbR3t4OibIqPwq/qkGt3qCeTAmAF6+qk1mZKLKGYRJ/BUKBxvARbyQ7uNdG+u
yo09Z8Sctrbf9OrnYy83zfJsyCgm2SjayuUkahxVYE8tN4NsYiAtISklRyzG66/4
/4gZgx+eS2iGdVGGdQlarMXSjNKPNn9b5UzgPWOepWbJ2vXVA8nklmryJX16rvIH
SKqY8nd4pRIe6aLUpfkSRerKmdiQwdGspEPjxQuU14Nnt0RMzvOnSMO5A/fdyoqJ
S4oSeBhpiL2B1CJg4GvYX6hhwKFB3QbLYz2jAnin6xPAoRT+wZCJ1Ks+w/h/SQAu
wQB3ReUbsOnp5dtgiRXpEPdWiYFxoMJxNJ4l/yLUFAnUBYhBkjyE2J+GyCOYjhRy
DSy2uml6e2Qgnd6zTEbPyaG3RDqIcBxPjrFOtWU0YfE1seXRNu7wCpD24c9WrfYP
G4KGOY5YnX9y0BepWCALa1WUsau7n0rCgjyd3MgvluImmPrw2uT+ZAH/hgw3pm5A
an8PDtlateUaDpY+P5Pb5cBIMsYunM/95wziRFs79IhGZ0oAqLYT9SEMBlctbQU0
V5CpjrczYC4QPfb0g6EHOEXD1UVUfc2RKS/ZkIyKhqEqVDGSzOscehkDT9Sw/E5k
M5OPZMm3wcb8HYqC1gLc1ZrmtAfj+H6Pc9dNifzOsGxBwNx8BgEUbcuTvdfkjdPr
PeO+cb/zict9w4SVQK6TEVzpAMRnoMbadAv06k+9IItp8EqP6jsl6zbIn16XIAJG
XPU434nNKvrP9C8rFqJKLIVaBXAtnM+DPW8QhHhsu/5pQuYh85HAeOLAccUg7PAq
ulJ5UTS2UQP0DJUadKcQWeMVwoNXkyPPN7kQ3alYup0m6JUCTOQytjGC5+1Vp8br
C+U8VCpY2m1hf3qXW0tfLw==
`pragma protect end_protected
