// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LfYCjnYapNRNqQj69E+CBcBbqU6dnykYARALu480COubU/HB/wwuBRnOYgqDsgWb
TZPw95TYMFW7oU2qd9IHpJX22CM8c1nR9SBUOmRs41spTumK1T/5ckesW2tQadYb
0P3IyR/Bs8HFHF5EMj2TYaVvrFWOaEy8aOu9CfUjsuM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 174144)
w1bZIeoDV1X24+EuzZQbYx934F5pQDyMIE4y50g8Nz1jzoOYSC0+yzpivnZiYi1X
xYYN9gB9FEj646muLJ5tAwsJHharHdG3bSVk9kS0Uh8FdLbgOOddUjeKIfUO6AIK
ChbX5/wfB0nPjdI+iFBKSXc0a2Z8uoa0cd/qhAnsa4CJSGwIGxn16EAAwogWUclg
OrHoNV+ZM+PQcuwRlSS32O1wN5ttfT/0DKyIts68zIv0MV9gLT9hEojUkbYdqEZs
hKxs2IrewRskTkyy5lNArfS6/Mr+/ARNWtqC6jm4YR8AW7i3YJGUdQSxafkqwGpS
O0zYdkggTFRCkzf8pRvwMpsde7q8joBKeWZG3VW7uBp7RV4NqWiV5bY+r7c8cLBI
Ia1IuyaqYmjhDiNpXH5bMW2u2D25rWs1ZFRPX3U+h1YayMe3cVtdFUldDzaFXHIr
xWNvN/bdNGPipDop9X6bP7YnjQ4u+0UJVoeKCOHvQi0asKwESw21VUSZVrLq+a1b
Kzfn8FU4GtYriQxEg1pAbBf/Kts4LeFlYs8Per6XFXqZPjqPh/zvS/RZKO68ZPiZ
KJ1Vrh0rpi5+8FI1YFLhByTzx0s4lXqTig7UQRAj+GogX9PkKiBpyPRUkPWhAip7
YCXfAhT0kag7hxKZkTrBrZWt2+RBE5zbkanT11YrF+ykjJEouBmenyb0V8rJOfxl
WO9kULEzDZKpEFWuS37577JnJVI4P8hFhyvIAvy/HkwI+LPX08oc+9eupQJcByDH
9I+ULui/KtG1r+OsY9QCvLU2grFoEED4nJ35wiZuclC/BS52yaa3r3DacWoUeWUw
5Gov5dobAAB2YcaeN03gRiqLrLbVX04myJvhSsdjpUUlToNn9jPOx+G/ZXx8pwuV
I3SyMAGy0x97MW9TqObea3APOXTX9reQNpTGc+P1cWPgdpEf11+2cuN/6sc7KsUi
C/A+hlnC8QMYoyVfp9jizFnbLdyO28WvEc6nNkA+1wF83XHi7/582hrImhGniohW
pUf9kRPBIPV9tidaj5W1wKz9nT7mm89jiZsqrrsYXvkmuO1T7DqZLxiD1yWu0Eyh
BCcSLyfnISq7LL94dEI4OFYP4NJ2NcQlCSyMu1WwdSt+tYDzyNba7BC6tktr1TKj
k1GZRmVL6eA27LJWxOI1KlWej2yLJahGrwWo+h1gAp35GkAQrHmCE5IhJhmEZDiT
DaqbvIFDnIxEgGL0rtd0OWwRoX8wwFDyy5CWjsEHPG9WfJzoudFZcElJGBUULk+x
pMI/vwbSyfn7+E0RgteMJZ82R6O3Y886F1MNvjak4L6asdqvS6t4oOfRb8wS3mJ0
suCxeOIvqnu+ZwVog0jyI+7uHcQZJ0EJvo6xoQdAVdq7ALLo8rBkFdRKkwIblIEa
5yR6+h6ckbc7V+ikUwDQnA7tuBwxpMQSbGbAMqyHrhEi8AUM6pxeSleX7d05wH14
432C8We+UL3i1GUgbkNnbJT+bE2IMOkEByLOGMMNDBACrX4eFBSSXPEcJ2NlqW+P
pSDd9Sl/Ua53cVFqJfb7sf3GD2wvlx7pBbGXlq7lczUqpKhjWuYBdZ5WjpNSUggX
CF2p+Ym0/FRATMO6sQ/R4IgoajMBASPowpoWzz3WNi6o4ttdGvTx4II+gg4/DsqZ
l5rxLA8LieikGnwKlWOJNaxS0Jfyd0sIYs9sUVx6wZJFucs+N/QdtIs3XVYjQT9b
FT1Qe/XWIYMuUtGgEt408o2EiLubkWm5648Fun5D6a0oObs+huiiwevIiiiqvtjr
fdySMbeXnzkVBHJWeIbD2Sopx3yfcMSJb/OVxT/M5sJxr4u9SCAUyKf5KxCMFn/r
+MWS87by5gcVlQF0qSngzJs7ISFukVzf293WVHJv+i0PcKKoaQYhzxgOlpAt3i0/
g2KjVUqUFQk9U6EtM6VOQHJK1rRn/5xUOCKx4Qp4Y8Xs4OAbFrIj0m33OH/ckoTs
CUYKJCvrCYFeh+8TPirXYY3lmc9Q273PSkFofRqLVl5O1C/cPCEWkZqXDAHwxKw/
gVugkBZmDvdsLmjE5kMBVgjbRmfuMkL3+RZcla1S0kWj9sgPvOpZj9gw/G2KSwda
gNQA06LtwY5N9eST5LA0i59az5t1TXcs7ANgc1fJvuL/gso5/Z9vNCM1PUXo7nbb
2g59d6XxQZ9xSckRKkzbE6sdj4XmcVXfu9eFAJFDA77j5xxOAUydv/gqpv1Kx+bR
aeiIjV3HDGm1oCYoA5ORipw1Q4fej4XrYBJRV6Q1M6s8VcjNQNXW+R+RS7uFxF+R
P1Se8y2/UUT7RPnTEDGc1eaPS0g/LyrVdJmU9TZPrgAfp+xRsvemqHX0/zyrthv6
Bs3rUs6vnXDOYjRNZ2L9ZrOU+xgqezWvH+Ijngfp2i1R7HgEyj8m6nKXOHaSIArH
so+aTvcY6P4+r9yckmFHMlqmtH/9bQihhVMtgBSRrSKD1rjbyO9WEtrL/YX7BRY8
yFKlxNETCVfNDonMslqOzTkHaN6aOTqX4hjxLEiu4NRiq9Fb3CjtvVs0ZnpUs9Ij
5kfHFK3v1V1aj6b1S3mVGDGOMnGnrdBFx+wtS/iQick4s0u6L9Iz2djW2+DqUr55
AWdTgHzMwKtcTvDXG5DDHb0ftGBEpgcSALUJ/evUGy/h1mjoibWCLAzKcMl7SG+P
q4lOG4wC/gL+hqiFulRYKX2ZpSIQ8y9RpFgv403NSsdv7eh3NE10HhWi+I04JjFz
GHfVqWb/8DkvUOxPuS2w/cRAFGz9k/KcYyWCNeyqD9Z9FIrc2DJPHDWzd+6mMEjN
lxZZEz1mFQqizDQ9eC3kfMB4u8N23kI3tsTH4fDN6STGSC53TTKmvkVsjyHd2gN1
gXIc8PSL2gQR1CCfNxtCHNReBAAzntIDSh8qCSv4qWJpIvbp/dNAEz0Dji3Sl06T
zsz75+GxxTxW5tH0SsYMmB9lZp4gCPV+qRDt015H8r9/s6Qxmf2qxhYn5dwsNJKx
fvoM6lOmBGV5UjkSJigdUS/dSURyylAyL7lOcdats2+CGhZ+rb7YhjNl1nRzmmRV
nznn+MafHdV3SYRulgMLKOFUMjJS1ZrJdOZfNyVW90SJOuxL69hkUjyvLd1Dei/r
VgwQVVEh69ivWgrQiO/QqoL54a80jJQgdFhxnr0+n4CCA4wNrZRa+BBbzIfE9zTj
2WciCVvwcPATZh6vMbvgyz1qF7eX7tOP6zEZ72XsYD5s2rFCLNf1sTTyiXDc1fUw
+o3W+sXm1ku+cLj6fVIx/QI03xaBLAlcJK9Le3PRgI6Durz5+nlFJg3coSY4N57w
x2PP2umW2ZnjxPyixvm11dRj9Sn0JBiuUHYSEPyn77kI9cwBJWR21jsj7pzukgFG
tCRt8cQgFZpS6q0fIeMAwUVUviYVv0y4gy3Ecu5JHyd5kXU6jeST8nKSLm33rTxN
l2qRIPRzjpshCds+34haSIWtNMsPHxc7G/4p9WC5PVc2+Cx3by04y0tvEEOIdK3+
4qaNZhxwurFqdTsfX9a57mlI6NAAZ/SpTaYc1IofUAR94IT9Wpr1aWGerWXgTM7r
E2UXEcrG4Um85uGN5BE19p1kFY2Y83+AB7gJnIMleP5XKfR47x0ABGpHY81ZEV82
YXuds4UXx/EXP+vdJxBkFbLdxMNmxbYa/gjlkU3gfiVwJPTmrwMxl1XgI/INCzKN
U//yWr5dETqS/QVD5eIP8vrRi2GAd0y/pLZSNUSJ+FhgN0kOk+okKyQ2evtYsv53
NC7Esl+17ehfbMUIzgraAV921Q6wKeHL9QCmpnVSlRgRGtYX5irS/+rQHY9B8HoK
mlvPpyKdaNroICsB1XnZwMpXKLkjSPekm1bSpMBqMWoaLrt+K+T2CRUwTcWhlSaj
rDxFvZ1GaBMD2fDnjE/k3cdtyE9oWfN5p8XeO+fgpZmxkQEN7yvIBgwqreegsBIQ
M/gi4H1OS9KfiCKVYHFY+hzJXnDwyZdCdu3L8eIqA6/8GAycxkgFsDbUHZd+ZRYi
y0+BoN2d1bKcm41LaGJ1wpu/LsaSe0nJCBRnhVKBRFeABfvUYY+NN7fdDGvqnWHj
d01YpCGPMi/jfgN5Dmpl/38N/WS+WJ1TffnlQ43UFEn5QztrPPw1Kwg6BSYqUI3W
YSkKWY51+AcjIDkI6v6Cuvy6rwAWOmhSkSEOkkcnQq7S4OM4O7Q1qjGcRBWKUwwB
wiuHb95IhDAA3el7aZRcWw7oRLeIexOAY8v3voFRT9JfTzFtaYVy0fEqhTQaeiix
8BY7apFDqmfNKvT4juEDmYgwo/Y8sPfHvBFxDz7ljx1mnkY1MbrW1yeDARflCnfn
QgMBuEzEUnC2gbieFZRSXQ1/9k2XqB91vxsn0Yx0PVHkBtq/8/C4y1o68ZBBbpjY
kA/T3O0w7u3ndXZKq9KZo2ScR6XO/wFmZI69BD9q1HAobKkv1PQe4vdDX8Gk3KHB
b4aCIMdN5JVIO5JVvjr0/xl4ep2CxbT3ugZEcSyXlyhgKk6dwGlghRrl0cEQGyme
cwdxLGNAE0DDXNqKzwqiqiJOmThscuNe4h8rG8WjAGDGvjuyzx3XQWQyrdxp8zdo
P7M4MivcmKIS20owMZGN56hzyVDKqOfQPCQyGbHb3sirqOSgg34FpVohwFPBftwp
UceLy3XcpmHkBn3JPMEg/npgrbHk0zJGVgQ6j9T7AeY+UYC6MBURa+WWqY+3gHZI
u0b0zIiWaATGcqz56FZp9UdL9noKuiAB6k5gF4fDxG2AGtJ8ENg8w8wJNEa4e5Np
pk0h9P2S16Wliw1L5NUT9fxiq5+vaI5ZaBvQjEBzxy46HRnTFcfdolTfy6Ozjkin
HCtK9/Gc9T5MQLvM/leV0YbqUUO/Jjv3iQoct8AhVlN4PLYhUvKxJreKnQyvEVk/
90TzH3m+rMuS3EnFtG5KYHXjcJB3OjuunPWzwSHifSHPCSi3yYlYu9l1cJllupOi
Q3kH0fN7wLyvhe7q+zFbaiMKonsvTX3J+NcZ6L2fBtUWH8gMLWeW7iBcKAbXXxKn
eMe2u5qmWdcLmKmnfIrpWV0NCeUpnqggmqXYncyT8gs/Vo9/ah2TWF4UfPUsfnIY
YSNKj3LuYNC8Q552EVuqsmunnps6mfhjspS0LZSbcg1ixSmNrkjNb7I6un5tqueN
6Jw1zif9M/YMts/39XFfVd85URgynLq5ERNHCCzH7nSLcVHKzswYiuOSpmE4EFkO
UbdKJcgRPelcPyvT3+2aYE9a/JffgPe6AEGLZjIazyj9ZFAqhD21tn36OYnb0mam
YcfGz5cg7gJCOibo4j2iKEKyLltlrXeYUrhiI4h03nPAwrDrk1l9c3aDzPxpslK3
AtfvTgMC9DiqbRWyj9ury+hB+fId6mN4xByseekF9xLQq+yjIQ8HbfOV7m8PcymC
RWld4PJfsOjfQOjzCBDMoLrSXDS2UL0AmGPKUUxXJra3zKjvjIH+gf/cQrG9BM+5
fYAu/cTzpuoz3ji2X4nY3klkmWrRoJAiH9A02r9y2qvGm/q1MqLkgUxGi0zb2N/V
P9j60FAVYBLe66Wj9I79Hx+GKg2Jfg7x++4rgxhByGLBht41gaJlHEL3F4D6v/Sd
3oDjYu7Ma7k5XlUhKT88gqeAb3zME2xvZvWcvHWlI6ZMJfBeO+FjjhcgveGfEDZi
DNBM2Ahv+MQU4RFf0q00+pxv3FTl+jZuuP3hbK/JYAuw8jqhPRogmGe+Xu78H75+
Ozr41/kwgw6+Sb0Gt/2960YF9ntn2x1T3F4IE4ZMScfVWNORgXvGyWju0whCfapM
zTitIlNLCaWA90fhAwEXzXe0SRr1RH5N4GwWbpMmG+RFZ7Ofd9Sz1OGAoL5D1NPN
qJBO3g2qxYGzLVuiA4kXy0TV+JWqIfbV64qVgYOt4cwonqmLbfgHlPinb+LgKetk
LhNio4RbCb+Y+qTo1Fh+K2R481FnaNAm8m17bWJNcqOUi7+8ur+D9axSsq4g++ir
lKk1XAedkL/BpsbL6ri/RS/qA1BgjFJ8iZ6qYF3NPXObuhpZ8iXIl7g9/fbD4Yro
RTsncbqOB6zCACWOrvSKDn286Wk133pbOKGva/67PxB4VLXJcQdjMMt6kFljbvun
Bk7CcXliOQpeRHMS+ch62HQ7jNpavZix0RY+tQujc/1s7ER/HZmPITKMk1r6qeY8
BAj+Ri7xLX0FpPobBWPsah7eyLq0vXCNIhpev69HobiUbELf2r+VRJV+DaABP4EP
oLb1netGKN9lR38qm/HOEHXGfnYcxVAFlfhwtBsAJvkukbWfRu5Pm/34OuqXaBi2
VZBHVC1ObWNQ2gpvzHFrsZq7AfkLdJDL+wayu6C3iteQr7QW96G5m3+/v04pZeML
whADmX2az3V6bp2v9hzx+ITfIRzv7lkVXIIh2S/3FnAoX+kAO2EDbotNodKwRy5w
XRaO+0BCBwHvKi5OoOJSgJYz9fOc9QQ/UfLscojFopiMBrvNk1WXXhoIquuI3go9
CajRCIz6Pn8S/sqQuCSCqluWKFo2Fb0/sQ/A73O7Mx64u6o+DqorXKBIa8Fgy7Gy
4CdCYqEMTLdC35jfMiKML/lwvO4Qzgm23awQ4FxBO/FE3pkLY95t8xYy3HMQa81h
1m+UliqNqC/Z47MJfMR7R7nuEDATFN8Q+qIpDXyiQianHRECrC3eFV3B5LX+vgMN
FGuw5F1gmRpOZcD+PZlw+MkBiwOjVeL4B1mjKGt4NoH9X1EC/wZUmZF385glvuPO
5PQyUbKJtu9emI54F4YCdNs35ogWieIimXEwcRUz6lUOod5YFqz+f0Kpx5kz2GOG
dYeVLTFT8skM8Vls0goFCG3HO2K0fb+nuqNm3vUT/Tpc4HGiyzS9bq0sISVWSLD9
vu7hEpFeI6nhkF6zbMfrxVMIoFlIG9KNporDbzL68IRVVNMgg4rhTrtq49XLsniB
a1msqPFf+G4YujjG+JADvdKwyM1NxSr5vmdG8ScQ22/yD5BQ7s9xOAwEa7SsqW4S
WLuvEeZXGvzG3feRc+QWgFqu+UrMV0FDGVB4dn2F2q8Ab9kkNJMli/enf86LGE4D
T4ph6BnaGR5tGc42wrN3FfCQdBVhUte/i9j/Dezbqic9u/opYwR3V80LZPbg2s2D
87ChXAghyFaFppZurJPLDxQUPD/AbkVLEQJDnqjij46MO9DqrU16dXY+YO8DKjvV
eOnurTYbP1KFHF/9o/f8ms2fKCBs8XYjwn7SinrQDvi6nRTPQIIf9ww0L5mQmx3j
6qBFH0ZP5wUFNTfGmk+zToa0GPs8xRMFMaNmc6+FLlENo3Kl6vteYmWjMgxMc0xo
O7LiKHKQCshzyGsnubdf3WwXG63PkV/OkRJnVXfREnk+GLBn7mHrd56qRyxgC4lK
M8mZyaijxjmQgjN965NQivoow7LmgPQW+r66TK8a1Dtb/jhzHFLpyWSie4DsBQWa
wc7CBmluEEa/Q6mtEvhi6PXbxfs5B3tae8Osnx5odA9ykLhxD7srQ8HBozCgBN5z
z9E8+qKK/Whx5ErBtADIkUhEsF7/i7KjBdCPysN4dfIgioh+Any7etfOKLS0Nulc
q+a0dGcJ7bdANT5XiVm3Xjh2VdRqizUZQtLnAIDOHrJ9JSGtFfTmUTbsbYQSFmlW
Syty1PjF5g7R0bScdD1/NI7BrPsmLl4O6vcYU1jBfAkp4Bajld5omZyjUwftJ2s9
4CIspHP7wgV61wEqf+gWs19tvc8ze5ZYaauaPWAtonlF3jjEm2dVcf4EmMXgXXEi
/7ZtpL9I5GxOFNxuHDFvLvKiJb7V43Gsy75aXasOa17wwb1HuCEpZFTdJN/Enu8o
SgWGtsE1BqYBYh7Nn8qRLvFKMG7kA5siW72NxqnW2Q6pL2QhzT991cJ22cSZ9QTv
118HXzxK3+013h/UjUYcSzsr+oN8+nasrYn7y45yVbLSgJLTzDAr3yaefiG80sqS
L5kd2igNGSL3G5BILvgXCErxowEK1cUv0CIqm8FX0kOxolKFWDLPJVeRue1Z/5L3
hHk8pKgTJyPwlBogBuHjr5exC8LMmgimmEnQqlSHGE6MKcc7nEAJOfLRmSbkRPTJ
tJiFwwF/rlNlUtGD5wfVkqA1sJkldzzAtZCdi0cnFSuxxuiKYKBENYTkw0XCfU40
8vQrxEdU4lKxhUAWft32zrWO1uVTTTNaAdgoGtlMMX9jQgTRrLKpsjsFYKpyMz4Q
utf4J2HhQmWlB3sOYWwLn9FvxUzs0Tnvetluk+SPxl94osHy7pHGBwBpuyEq7lM2
Jp02zEdMU7IPY8rOO6+9p8UK+4WDBATVPYMTkzWWK6NBWrv4LKdsrl5RL3l8aIlD
c2t6f9FRjFDD3vlj9A9ZoZZr3xet29r//t7Zp0hHSoFAsDK7LLvJMx5SABdl7WJJ
2NN3TDhSZGQzCcbz3IetIidaF3mYbtrAt8DsbRR/v6WQxwtPECGUedpzCQv0UXbP
rKHb1lSFBIBbU/uPUKe1g/0sd7vvWlDy21M6+jBNaLeHnqLOGQd03YhrpqWhuL/I
Vue6k0IKZwznEqNMJMg3/WzNlXw2bQAA0WXWymyrdAALs1AH/oNsaEmbamUtFzS9
CfjD3optwOzV8i6jtkN1+rpIHiL5Jgh+HtDwIreB/6cTQ9zkzgScFC3sEQR7N38a
FPWeKV8Zf3LT40zD3G90jpBAylP6Az1zk6ZZCYF6lHHp42PEpilkRyK3B+NzAgRU
bc0ycnzy55rG6CooJ1E3fo1p/R49HtW8lre06aRQOTGDPFGNctrLpgLIKGhpy5Vb
8zhlsgZ1exKtbQrbt45s7xclasDF3UjdsA/AeILojpkKgb3F3dorae4dk3GLwtEV
UzZDOFh8lusiNDgKExZO+QyfaRVKiCBbJc9fGLD7GQvHBv8SXmquo/c+R4cbkr4h
ttm0dnH060psh1pHvdt6BqC/rI6gNq+iRdkTyAyZI77M3WxHHraa73ipKEgcX6O6
q9OP34foR5HNk1E0qmaAns8zjzAaTe1mdMstTpBczj42qvtmrh/ruSeU4H7QBRBp
ypsHumA6VOFcV1JUPEXky4CajEGFu+nJDNw+dDnBY/8lbDLLColhhz8cFEqeObul
27ao5ibTnQ1RXS97SvWwcbi+7TQp+bs4Mg0yaYRuxEugPWIJbyLBj07PAuuPxDtS
SPHJuy2R+1n0jEoRSxv+Gin+kPzkeJS7H6EOZ9VSoB6Y2tqjapwvhU511uolK6B9
qgfGDre7eiU+bN2YRGICNmLzhd33/dXBshWYcmM5Y7N5Xvl5yAM/bgzGYOztBtfJ
uHTSkfhXmvwXmD2qBoFLEUoiF5zjwLDIGqUV3pdUxhycAz1ANXilGsg2oUHf0ncF
cj1frB6HMZ7Kxesqdpice4C+v2pvgr7w3RHCUpedd/qZkdZCuWkq98HWLv90OBId
lXYtf37ZsGqlIuEsDWsBdW3mKdKvPS3Foc9tdp/7c46zgxvVIpH1JtwimQ4wwKsN
iE+Q+3pfTWD/EmXaIDcX2OiHD39x3wU1PUmAs/YyZUZk6K0KIlD7qk7iE2Q72ymB
FSpJqMVuvAvuKobToG1BnH7FpHglHAzLgyWPJHnhIvy46SjwP+oTe+IZNo1+kwMb
vDTZqsUM65bvyh144/GhAv2iBfHJ1KWVtEpEejzTyPAH+KWOdOrZ8rl/LFXAmt8s
uO1YZsuvTKRbywPxO1nbG+S2ZbIHseCpIbU1t3ZMyoDc43mYWYJvbrvlu6GZ2Ueu
rppBt9knfLXcjYdRk/GelAyjK29kHHZiKmWRlCVa5dpYPLqcbXhYNGij1uVswayf
o+loxYFfquIw7pPREHfN7iasTUh7bddQB4dwxX1asOad2uJBsAwl8PNHPloqu5Wz
AGmaHwUC3NoZpOylQatjxJ5OkDSwohVoQ85kauKwzBQMzpzoCxch/o+r+nTTgPTK
VlAnTsWUd9q3MwA5VDJOyKHynA9CzYi18tYLLvzgw9n9y/6+BTogphbwRCriYeMi
d2J/3uOVa7pob6FL5nBPdYL4LCN3EXVjNM7TEHlubOmGNjxKcIMmoDudRqNGbwWx
NDLRY7CxvLa5RSrJBHB/UWzdTX9V/LMHzua8yb1zRb3DKSxkLhfjMRYP5Ykn9n2f
Jf2TJh2cxa24RQVT8iO0dVR1UUKccMiN7PTM0SV1BVIjKXggzyTiigV/zoEbVBsF
h2l44lJWYer3X4FNKAXI/GZ6JkVQzTzSwetUPXKJ6yLzCI2DvTucea1rG8LJ/9d+
b4KZCUVrUYayTtpoxYZ1z0qH/+bshSNKYQZNz4T7NuFmYw41m/jUMzql0/y4LN+q
WPcsIWW5gxz3J/S2mt7BziiWVyh+Gjk/6nGSogfPF06KQN2gxGnc/9JC1WC7zqdo
paKaD+UB25TrNYtdNnw8Hk5vOIxDJzTrjq2r4Pdf8lxBeDXHAhZfo6kXfcJos83b
Qussto1Gb3c3TLVm7t7Ol8t8BoQNZSByZnixpwmRESdfoV5UdV3pGUrXx27uZrZ5
CrHgOafM7PrHdwkbpSVRPSRMi6ylRgU2GESpv72sr8oUW1dSIGtIavACMoqlQXa/
Mzijyl+XdJnHCsMz0RYc/uM6vEs2dHevF5u99dglJiDcf3yZylaQO2CnPijLNqoi
yDahY307ZFlyTzsT1kZ9lhQ8/StTPOP5uL7jxFz4V0jDNIL5gDwlBVOVgjDiHnYp
UKJ7tZaCyO4w59q1IYAlpJtNvmAUIlbtVVlEjZH8G1GLoO5y2r6nAuYhozb4HQSz
ocFAxV9qKoc0tccIsOzDcwehTsYlHcb/2PQsxdVThVVJ+PpkoJg9fsfi4g7RuZAH
zdgzt4VAc8QBqlm4scmLRhl4Q2IDYACy4pyjKJSLSu0Ta/dAsclH1/28JB4WteDn
BvATEl1P755/wv6wnsCekfIn1GJ3qkShKBjCW9D7L8hscXbcr08EMnpKKBtXBh2G
bEnXc8S5Da2+s+4iZC1nDdxbxKg9XBweSkME9C1f/AGGeCO1fD7TDXPfxtxzp7Su
Y0nTrCdvnlVf2ixkAIavcs8ZlZtXP6282s5AT7CTKDe3eIw5Cify70cUZsHGt1Is
sLVdikHNfSE+ggkDEa6Ucvg262Bkh2gXJppWSZsLoeWrKNfHZiuF2E0nJHJr+tDV
xe5bXnljFbwWmBGs4R5za/tECeyP1IeepF3JTOAXbOq0MeWbyS4xGqqnQ+ScNqFZ
52f+J4WnAuUDdjmsInU3CiqQttrLd8H7ni2qYtGylmtX6rDTlZbi+zIfeKzg9qPB
9saZz1krsdvDF2RD2oulkAMtj82DeaKq4akjZPOB4Id8G2kGeYb950BSejrqi2vQ
6JCoLmDllIjyXfAq8OlpOnbrJmVbVt6YIXgkkm3tdxsDd3bB/EG00ThSWZ/7e5Gy
3Sj2HQ4pSyZkYdDfdDPPVb2+lCngo0i9HQRrHSF58CVJhztcumQYh7vvGbRXQU3S
qJnkIC+Ad80rl87ts6f0TfrgUz9fvzeN2bfHGJl9ouoZM43cmCmBdGSUaiVoj9ji
iXaNFTPp+bN1vHVJIQ+UvwNE7ljPvNr6AO3sEcIv5jPVX57xTrJXkPFDYmvY225n
RdLsPZt42m61rE887HPfEyMGRlpFOq5upCyO2XfAHSaxxgnJX69jsEw5bxFJAsVi
bAxGlsBhT/DFTi6NxYCVFwgbs4ZKfQGlgiqxfPyAIJC0RYUb59F31jUCwHYEEL0o
uMZnRU5pzc/RO3ZAIn4y7OrwZHZ2MKtlrED9ENF35iNl/6fF7kFXe4kHHR3OqsBu
l7fVnyToc5bO3KMzJoSNHGtraCJQRivL8TnxYQyt97/ZC38z59z0sy1v/hG9ddOA
EGHd/gaXbyPqEjEQlIoOUkij3+vahedPLV6HXgZeVA6xmOI77IeSdPIEi/tUuLVQ
j/LQc8NdP54hsG57NYn3+DdQZXF23LD1hlS8LF4LvvX5lMLu7yj9yXywA40v73Ib
KjhlYD6hDcW1rVKgAm9LL7nBbw9nAN4a6117dtIYkVV8EBha4PWdlFRZbCteybBI
w1Sqb5EZurF4xeMFgSccpO3SmxL8AiRFFdIsmndc2vOpQu6+VEZDLQO2TMkjpFZH
pzmFQQ8YV3j8oFiI6Zuylb00hGH0BF/wgnZENRI3L/AFPVgJMv7Tlb6p9lLD3ANB
eydOa7T5SDrCSA4irB2RnK8oT4sCp0Av4TXZS2qBFPllVPx/gzmXrXlDyTdVQum/
b5YxoKCLMOCML0ut5DaWdkvVx2XY+O28FyFYd8kFrin2zDlu9ayOOXFAzlvVpEQJ
5ETP1nG4lo1+BXa0nx/QOaN9yVuMqGDPpvIrXkeq2sR6b2uRgdvzpR0bW+/Ev/vu
eLXD9YnyvK4ZS702tqaCR8sCXZ4FSqftD5KJP84pm3nnZ0GlpirlCbSti+EgUzJL
RcUb7xHQIdBmVwvWHDSALk4HFwgew+lPFYdK8L6BzllixBYh/jTDK6pO8dSlYttd
3rcr/oozmT1onZGuUnNLcNoSmL8ECdpdv2dc+YyH1Kvb4PHwkoAfPox+ftvo2QQp
X8O4jkFQmg2ZiNmLVrAO0ni5ci1k2LdYF/YCN3d+rsh0/nMEOymbwv3IyMFD7Mzr
a7tREZYUxd5MyTBKydTsV22d4Jpt0vcG3GLiS26015bK5j+g5fZEIfRtvPed51Zd
M2ehstx1M7vyY79ke84umdP2Da2Ae8OcDnIsfCD35815NiE0IG/jYOUwpU6E5KFb
T4s4+MmAfXt891XDPdtW/M/T0AHGPmR5Yewpz3eOcnjrA5vf/CDn2jRJw3ylN6BX
U3hreAiFZk6cidknz5EgBofjuvb2rDuu/7xWhfq/l0jSKaown8Dtb4wQ4iWtdoYy
v5FnPR4NxYWOHyBF5Z3SS4NR7dK6IpF1eSYb/AR6Aw9GZXZS+/7Cped5/15Q73mm
j2MFi932B9vpw5WpLM86ws6UmqO6lb4eFMGhC6GP71i3kTSbXZmW3m7oE75WqhgQ
CJZDoV/6PWTgD9aThmBhWY64a14ZXUcJosyTry+tyW1GjnYymBWn3obd1U0g9xCW
xxlDfn3M+rt4EIUdvSnXWgsHsKHaJGMzSItZCMdCJ2pULkccjqGsu8vsDXR8J+Hm
kCDGvxOnyDBKHP6wJgwYhM5jmWWnjuRRr0Jo4WknosMZuFP1bRN6IEvYTx3SIFLz
ZDsLxpJPR5adiygxtoLThvppnQ0AyXUD9a2cDuM1zUGpUCWNCc3LTaoo5oAS0iVm
/1wZFPDDTRSX0ACIBAAei8/hCLz/WCRvh3WJ1Stk3sUFRXrHCfD78S6hhxF0kAa5
UuhhTqmJdd+7z3HzdMjlaegzZCmyDIoi/6GqqPI6WBC+Jmu0EavtNLPtmvwA1ogs
LrZp9lD5kK81fPh+7ryeEaiulSE/5g8/64WitflADdLVpq3y5FEP4TVG2ybKu7fw
1eGmv6FmtMVpqrhPnG9mpRt06RTSzzh9TFIBquuW4jUQTrs3dKFvGXUdmDGBMIyv
L7Z0YAdOOkIcF3Vhzvm36ubCp8+MgAG++7l+/I8O9TdGDOOogbECsMMHiv6do7l4
A+BtRK3gtJ8Ogh+UmhL77cVfTGz6xOrheJEYMwlZiCGZOLhuuAy3vBIU6ODkiGjt
2KacC/sMqqhCVCPNGIHnCQgQLl0iYNzzSXj4Gng5ucPyOaS9lVD9FtdmvnFGNCJH
EprfjfAKMBvlBwpnA0MFNpCtLAw6o4CdMtlvZ/GbNEEIthqJHZX99SgDNjmwhQ+u
ehC+yTj85GQ0uDqiiUUN1MSBW8x0gZ9Fm2RS7QqzTMvPG4udJL9B1SlDr8jBCebD
0waf7hUclz7phfM1TP7T6HIxguJ1wSooLPhoPNnU0wiKVwkglxGyWbCl6BvbFYm1
gSJsW8oYUSowd3YbEpjY3R/MMua0Nv0ROrxNPMozhpKUQKZZ3QvpQwFIb2t9JcgM
bDz0p/b2CAvDUptkC4R2tLfrKnUBSPBfsIoIbadOCmuA9vdaEFcbxr5pb9+ZCUeZ
LVoiwFYDKqLiSQ/r21Ea8Pe8QK/GynULXTkSoJZiMIHjfTc6eXDmdBe2M2hJbJ/7
Hpqt3yXI+6fAYCeJbQVHinFaZ0C8E/xfugqW/eLUZA8H8LdFODvr8AJWdkY/HQ43
ZtEp7UJH+u7Y3a/kg8WNF3pPK3GbBjWTJ+0Fu/iH9812rKbxWwC/yG6fzlgleASj
hZC4WV7za1X4Yr2TZqNchPwsClfAKcXZyLMdS0oEP2oP3HJv+0bpjD8ONdTewypp
KhEOkvfPDyZJteHw9WYXrFgJH6Qke2PEsryi9LvIo/E9Hn62smMmDqNA9o3LRg17
qQI+yeLLlbG7x9qhNNR/UxBl2VJGBQ6UvCl2lAwHkMJW714TwYQHW0KKQCR9gJAy
93+aYcgVvlTKjR7gjOKP754yRodpyDi1hK9UI4xgT7lASIyrhhc5yhDaebAsxtpW
/CaewVL3Wstc6a6ot+wYyE7isF56KTXr0FuqZ+hGExNnOAEEz7dtLfbTil+r6vtY
m2aSt/xtKLcUDhUGUI51Aw2lCaN3bhpG/XnGsU+s/5skljrJo3DLlrq1EEiFruTK
l5xMpr2jeGApveX8shl2BRtaPdjvno6MrBgsaLpzv6pAHAQI68CFLLcErzzslrvV
L0idIbjrMQCAg8xsobEcNrgoo+inbPiMYAYBBBlAH80vZcY5RFPYAxzC/M/MUfZa
QxLrvZQq/dT0VjFyGdD8m8Ygw17p7MljwwMhd2fnbn/RLB/SeFrcRj8yZmW65B+D
paoOFmdzybHv3hfoclzvBT/AM99z3h3sKNZHkuU3yR22NrXIYqlIzVmrkGDboZ4z
snPLyDhVtGJ2asYRZyIA4LGHbAO2NQA5nBE4iVqCTW7inpfb8bzWxWTSlbkLHXX0
n8OpZ+MCJW6IgklHdcWxV4evJ8Hww32vUqPgpWp4rMk9JBJoz0t2foHHEwBmtSG1
fsAZy4U3XXISgLcMPyImsi8Lj/PEN6hhoONUq0nb32P7fjggrh8NqEf+2+p6W9lF
aTn8Xb+9KLmP9hfmKvOCJ5WGEokBCiez9HIEigta8XJl6drBKH0c+cKSkuKJ5SyK
cifwPgzJSRy2612q8furo7EbOk6QBiuBo3z3I8ab/vhjth9yKbBZ4FmJy5+3Brd2
gIbJ6rQPYdTlaiGVOGje3fKdxty+VkTsTTSZHhVHIBDv4MU1kya27/WuB/0S0QsQ
xHTT/ApATBf34NjXnrkylZIlyZ1JO8fGaYUqFEvcbbzXu1zD04toRlMpticU5n3w
dy8U5ns5H3UfBq595vh843fQ9SvcUzOKVp8EkK//E8brnYBMGpXolfvcXhuYUkhI
o6j8fotzG3KmBqSnHKZEzxkunXF4ERR5mkKyx4YIVf7nttGFSu7WulQ1k9K0dFtt
FZoA8Lnw4VdBg1XGzxklcFYCEPKy6t0Uaq2hecllb1ftJUW6OhVDUJIU/16B/b7S
4T5oesi6JAj2ZULhRr7am3a5j65c8ygf+yjtHOjS8ElTBVBU03HAcSqTxqQmYEFB
rV6q/IMsTppyEYfmgXPU6xKFj4DdIIw/Q+htKDPPDNt+EGnuVIDdIjTQa5Aho4Jt
zv+2/P6YCJoSlIZqOECnWP8UGtAm/Chxg49H2sp3uVbNo9MuvT4eTGWrANpBhK0U
2BGRCs2l6FmBMoeW9TVhZlUaSpQOlJvIdj+MQW7pCPWhy7m7YPSpwZxq73OMr3TE
3louwds942e9X4QhuhTmNV7F2agubD0t2APteKfIhznWoebA6iH5o5IJiALigCG9
HFJ9qPgo7FAqcAHu2uec2Ct652yidNi3A8DXUV+1U2rQ2WJKWkNudQeY040k5/Ez
Nf7MxXCFv8q3dEktV9dwbr7j5u+nZxcr9s4k1seFEDQGOdLumCPTOPZT5MLgsRQN
fhaSi9DklRvjFJ1nNAEPL2qfYb9LYLtcU20q8m/PPSTI1yxTTflq7NoMAnttKhd7
v8MZXmGuxcoEHNRkY4x9UuotDYjcvSkaCv0P/9QkV0hF02FDcW4uvYTkzm/9WaxH
gieqy2nedRWBmFk737BZFzvluaJsl8qKOOcJU6XTP0wGrPs57susVRRsPVj9PxHu
eYSzN4NQzI2JzoGUTPsEo7PlMO9uSFwWNjIY4jHly92ucYNAvZfbUxstLe/LgjCv
1/7GvcAWpIkfSJvebqMrWdQaw5/qxbJSJQzUpCBpakazlFYNfv6VKL3QFiRwxzQu
mM9MeWVUTc4vubTSHYMyzDikXf+B1G+ohohtIUo1n/mx3vgrJlfO0hQszg1rCFGF
AMLq07L11PeiSNl05/Gq2RUjxSMzzZtWC3uP/z5zeKV3pam578DBKXezWXgAwlwk
16ErNPE2U33N29b74LAHPWKtIKXvOeaQuViRDy+5TIMo/mTMTb/moKJo5knlECCN
taN23NmDKdTX+X6kdggXeOzvUeICb4BV1aqeMsknJ5XgY1px/dSrrCSLKeXZTmvI
5Ypx/1cD8REjM/VB3hNS1OjPr6Gr8GiTvtIJLbB1i0QwYlIX/e0yh9YCb2VDMdcJ
QE6fHTae+w8xqUZqSjL92aNtO2R1o+TiScwjkSVtr7pnikoJobZyAwbsCEhKrQ8r
O8TEOrhnK2vmeOAl69WLX5WDBstMSY7AjnKsroiB/LRF3DBhOMZxrZZ6Hh1thKce
ig8PaFD/Xx34r5hedRBy8rN08HaHaKV06ihyK/eo0vSbm+hS9XZ6uH3buWzw2lbO
VBfp4o/g5+gFBxt17q/0wL5SlGWFGwV5EZd58A0uB6PSnSM+TOLx+tF96HQ20sXB
6JjOtiDHb0Ah6SJXgLEPgiY+Hr65cNYjDt3H7J7dWTU7q8dUgFgAHeZlLxXijA4I
xOkL5fKuVDXg6CD+saBfOBDWUIIONFjm2w4zmfZEzDoSEKBwWaKwaenvRaVwepjt
Xe1nvCo8JxVKlaZDa5Gs2X/Q1E+AGSjM8wf3sQM/NU8X4Q/1/mcQwdoBDwIUqdKj
cqWg531Ch+16eCnsrs7j6GlSWaM7fDdMPYbqNZKvV1BcXQQWhjrZXTgBSNIn1Cnj
Xh0YMx60rKNAMs7ngjmqDY67ZRUsIRzu9cncLN7LcfUgyJQwz9l0WMXbtOKulGkV
y60BKmCIrNBBi2Pn4Rme2Oeu73hNxfckl45wuf6aSgTK7AN42eyuZDIQHGukZen9
/sGEvONU5Y6qRHseTtvd0iQmSj2jzhFDJOxABvm80kN4kXatrrzKYsWSO9MYyj8+
ai3Ysl86BA2GTAZPJpfwud1nOfsGO5w3DtqND+3WTaJBji/Azdga6a9jPKI0Ifu6
O33i6+LLQ8N26rcuQAJpkBJ/8N5ERkhRP8j41+4I59T0czdR6kOWomjAMmWom3FV
HXC2osaAI0cZ1Za5V0aplCBltUrs9DnGD16zAsTHMXPNjYQwEMNxtBeebNAsmnEd
g8Zf8hw78uxLsXLUQc/z36lb6ts9zf2R5mVNpBDRxAnTXTkVGN092GWA3yU12bJN
Azm4nupwioO2eiGrk3Xg2yIwIb9KC2LNsViNcEIjHz0itJJylsJYa27FkofycI9m
8YywDupB0DudwbsjCBpREo0rSENgpvKPFWAclSKQzoSFI4rBvJtnERhOQzN+kd+c
8dnYJwwHq2pEQ3iY1xU1ao9NRZpK/vxU01na2eXJ92MMeET1IUwQiKz6jGFpVuHY
PzGhXKuzcZqQ0ef8L9Io4g5m9sgl4XuWPUBUa2df5inRhI51K7k3ZpOnb6pe2bIz
A5wiNFp3suslFy7D3qAB8Q2C7gfIZMJEXbdMXm8GSTUyhrvvo/ZWTaQMnOSI39dk
f1ZVEigFEqekpZw++GtISsO5/1wkPSItMMKN2qAh50OzAFPagtbcBqbhu5bz9C21
RhWhfHUkO3s/wp1gEfI5pps38D4xFCsdE04mpC3b6rZU9XhesTS1mw5w71wH7VEI
SPm4kuyi9+XCoJjRBxkg0VSByQIPXtejdXmrJq8QfpEBaVtvjmWwt7birH0wH9S7
08Q/kFWmkLW/ehNrJwxRvQM5fTxx/rdVqtO0AS1DLm+/oELgBgRZTfkO+fUj0Pn3
E7BFhc/3L5GmCqyYtJNRViPi7KX+Oip3QlLqvsXDpgqH/Mn7EeosF0MKDXiPC0g9
zefitUJ1f9AR2yg+dRjJSIy9JfyVCeIUGfhwQd5MOA1HieOsRB+cqTW11Ztjtse/
48paY3YkhXlrA6D4wvNwRbVCb6p/yzeRf6A1wdDEwejpIs+AxF+1EZqZyFhSu+/j
6FpXQamJOPGQ5ZFUtCI9N2BT3RP3WgSGSb6W9sCTGGc87rDnfH90kBUdTG5H6IP0
HCS1lfgkcSideqiITD1xmm0J5vAmDXvpqTZjhPTPpAialZRj1FPi8NphgPhuzWMi
BRyJc1xd6Beo2sEc13v5Sa2nnudvNMOXnhT26mgnATAN619NztWU1/AZx8WObjEz
PaB47qoFTcB+gvNYX33oqasWv/kwm8MlQ2FQK1PeKnciChZTDjf1s0SBGp4XijNV
CTgAeLVUCAg8g50KWnzXiBncSqlR6zCqqY0sjV+Z5bjVh9x1nxyVO88D39ftFS5o
68GXvMrEd/XcsRVN/QDgP1El0Bd6AC70I4PWUE6jWao3wjo3mIEkCqb51E1NYgml
xMdCa23RV3YiTQsdp4pT1zbhWPZ639KyaWS+AntO9PDm9NjNOchdPfeRrJRM6QMo
jkFZAmD6AkUDxym5xvIFkZ4D2RC3mCEIiPsuV5zjFCNq1N17tRY942W4RJfRp+8i
ciT9RI37ld1RJbsY0z+JZTfnx72K8HSpGA0PoszBP65YPPP1U9abHEalT/BSlekj
Nn/YEcyKQmyJA1XMq3scZ7iTmdV7AM1FlHJzfw6slUNmjy5D3DyfCUYlDSl8e63k
jfa4r1ALPSw2wx99n1PPteryo/vuNOt1FlHa9Swebbt/WYsj+zDX2oCQ08Zshwxh
acnteWBUKgaJAkDXFMbPDILqu+hy7ukJs1HBLz5fwDFjWpVPbm6eqT6Aqf23qzZN
DMyTr8VQHjmHVW2rjdELn1gzmTHVlgDvDn9WB+GZKwaPRWy5JZ89CwWEUlLiilDA
6GFCbU0M+4pCJdW55aXRHfmy7M26bA375jMsNiOUlBRzdFuTvmHsPASZkjQfCIpF
rJGTDoc85Stk0ScUIZtCToyS28GZ1OrQf4wVSM4kGX+bRWM8qKuoEi8Gl41V+1Gf
ho57poSAVJsmZ6RfP1YuroO+mH9DQ7JhjCJOFS/D/7Q7nwMmDLKVwrbuGgKByyU5
cW4m2pL28spIFJehUJMmgGMx1F5snEujxxrW0f7ClTp7Uom/JS3h8hnK2FMyI/SP
L3TTkEFj4lrhgL07eeJS+UviK/VSQay/i62nYpQfnyjzWUjO0SQ/vEfphKWr/bw+
CmIDrGNt7p4teAvylS/s0GumgDf7OlsaswZT8/BAk7mghmi2jkHDc7Fm5knCw3bC
qupr/cC6fR0ltoD96mdY5N++A4DaxlA45XlXUsuaA9UQwlmlb2I1swNOWvJZaBYr
EnqIzWALD2TaigZQ19RiFBWjTdZGLeAceHcWUrtjifmXOGTJjcVmBLcmMMqxH9Qs
8zyJBEimeBs/yQX7fhcXrHZx52B0Ljo9vPAvdBunLTkEOST00Xq16VZNhqDIfThF
265k6TlObrjxaVr6FzOWXrXNjXAXUJQyRyq74j1YQKrzdf/Yh04mO+ndozOSUM9l
2qED1lUAkgusFSPrIOVcUsJK0ix82VCMh6odiKL5m5FhttzI3bC43p+R1wUGhAbJ
Rjwegu98MbXss+UFdZpgRqhq2iRNlDhAYgXIBA9O11Uxxn63zx+OYxKEizdFwOkP
OHugtiURyZwp5VqDKYH1Iwc+rCQc1m3BK99+l7lGbgQ2mhIEVJNI3oyeYIwdP/P5
FpVjDjEC19jQQt3ct2dXt+WX3wQj/4XHZZAPDssp02Zq9H95dxys7wc/3UxHb4Dn
FMlTOScyt6HNLAKi0NCpdE/ZkhO1AtuUsHcbEjXm2NB0SxHzVHPhJUyOmRCTF97J
8lCBSFT8jcqvEHKGHpJT9IrJTOdO1G9ADiULbTwkqs26mKKznyKMEQvGQhVl8wIv
MJd9eBJKmK7qHjcH9EHDcAUjG8PB7X4nVOo/d6TYUTC/STx/6SnUPogOLZlrMU8G
CsKXpVeLjidGwAJ3/Nlk68sXEqy2y6R5QAiniPQLs4BPdDx2WgPqbsDMkImVCOsD
x3DfmFpvhw01rY5QQ4/j1ZhpRzaZvRdCvUX4aVXf5+PpTJXJsIM1ahA1hE2ktBuv
1JTR8bg9rwS5Gd7UAyMdVT8U2cLo7ggcd+avktQjeNU7BPynkeqwFBMqL0IPxD83
yGlUXaMWrCWiTYYQeariq1Pg1jdjBWDwm3slF6IzypAippWl/MYgn04BF2IsVHUb
RzvjtvxFi/qrSexIKAzMoPBwGUtfoLWXMo11WVXTW+e+EkHLLfJjR5Gks7MXnF+j
eNWV2y+zlRsNapr24A4R/lYrCiWrD9T4l7e0QQEoywpWjBiKCt7A3WYAbeUBFe1B
4TzqqtrZeU63sjYe5mPhMV8yRk4QOiDU2Np9NBsrcgo9fUwway2AV/o4jiY8kChL
+yiCIB/OF2zXZpXhdCWZNp51Rr1WOqRn2sRjxXXjkgAzRiBBD2BpvgejmYRJHwPz
l/jC7zA8rUvCQJ3d9G3TKJOiTe2vmBN6NbQ2fbO1dJEmCBimgmWC9IintodPp5iu
7L6h/CMqVl95hwSoebd4q0AG3NZtN9M97fVHk1K5lAb7+3lv9Gc3A3HIUMgLvS/y
oKVNtyX+SQC1PrDFMIK8AAA9655ppG6bmqZXedxZOfj/YuxvCzGbI+pyClHNGwqd
3bO2uJKrQ/2zHOA1AwUz8eimrnUGzRadCHpYZobRpisAI6oCzXt0uPsUBdWNVu3F
T6f1qn6R86v3SZNdi02jOFiViikpHLwBKtIyZjTN2RZ87KUVjXwmIRP/Uyavweof
bxVpcVx4p1KEHbfYZA8TPU1X0vhn3ecBotFtnSUkyLCvfSbjtNZF1zn/3WSv6+oz
t3GFQ4Q28VaSf3B8sWdNFLIFvMky/7/9sk1vedOzGqJesXqDs9Xy2juFOPyR09oM
jNzM2ZhagKdTaCRwLFKAumnm6iezYgpRaB0kxVaW4pEBuG6WYwIEIQkuEWcZv5aw
CTrGYEvhYP0ZAFO4czLkoPIWkgGi7vB+SJ7nBbfIwivf7F0kMisfprinD9bM0t++
YN3sqGcOdgVQ4XlCBaugZVxtMVvPU2BBlUiGFULza61GY/DleNOtXuPo4762NCqU
DT9r1EoJz3+1C7As9wn/VirDEDmaCNaA9s9FrhTQVwKzMbnjueq5evX3pJ2Vi/S+
1fYqteDZpcyOYS8Q6YwKhaZtwsoWCPPfO0F2wzZk9zQAbsQ3plcrie3cZrsuUoL9
xsrx393TDApHXLjLWDiDJCOb0XIk/fs6+AdVL6W1w/Jt7Q/Zx9UMHn67xvZkWgPG
uiK6MQ1AvLs0TtbJzl53o6Y1d7K1Zudv+EpCYKpWsVvNQPN/6GVafnrDErBCxLDA
34FPXYJqFvwXbr97tnfSKbEkwoXrJBX9+VX7kacf60dMSpJJ1lLzrgnDjcLerhMy
Nb0aCx77vhmiFW47LmYFq9Q+56Q/b6MfP9RcqA2toSsgzxEmGcEmxLjruo8YW0o1
Lk+bN3RVEZHl5MNFkivLok4Z59cNa5KRvQg2cXGGvZyhVDKzW7mW400uHvf+lqUh
1MpIxKo5kKlAWrPLYpvU5iAnRuY+FYGgr5Ym6UQWVZcGQm/WXDXcB2u4UrZw+y4o
hjTDrwLowSwOkKo8SAevJaWZLxqlNMqgB5IPZhZmd1ZqVWPsvOqV+YmnX4ac3p2t
2UsvD/yX06JHWd+pZxNgViqHUfEa5Xuk/AFAjm5ePReaRT1DhBgWPPEpdr7CAPsJ
fH/nN4dreFgDHtl4V0boMoUaxIIStpV2CbuSaRWje6fWAvWw7mN8w35w5/LnOITU
30u9oN70h7/OSNio8c3ZOiDCKTzfoYLKl5+uZpSN9jvbzI+PLFWRcU9hrJoePU9o
GUIRfSq8rJlmTv28ySghGrd2d1iGFz+8C8cTVDkKKz6h6/qMkX/sUc0r25X3fAtA
bztADnA2/SdXKjEPOj12Ey1n3r4mX8w3PzOfjIV0cX5qxx4ZLjkJvMq8wvtk1L0i
182qQk7zRkNDgyjDfUNK9IVhXumbV1rK6yvyT7a+F06FU9nRgQJCTtMA8n9CliH3
AVUSZ0hRdjc2xBRiP/LP/dnHHLqfNM/dfO58Gep4DcXyvpkt/2saxtFgWpNYKgrA
LCx758gzRjc3VtHXZLwDJREJlfV3n3gZiHWq83u7gIbeDfQPBrovh6EasUv7nXPG
LRNLHtbFmMxwu17KuvF0DlzTquth4VDRM6bzierDty3Eml+1X4Ebd/YS7/vmIjHh
H6Sk2G5MTmOXw99d91Oiy/bT2cc+5JOE9GfqOsNBpFHWY5pgnAUvt8u4jXBftE9+
gBQZkGlo99ahkJq6c0Dk5de/AeMqR/0iNJkhnGvruNDLLmpBdziJ/wA2cTs/e4vC
tY3EUGU/LVJJjohlfTfdJa6EbNv1P7ZJBYpnuD9BVju30hGSV3wwLiAC9YZiiEp7
WVGATtMm3WvqsQKPSpazfnccw2RBzteBXOjlfiBxwIdc8h+JNvUnUy//hPK4aVcY
g5BLqPlLvJ7ZoVKbdLJfQWLRyaZ6tJp1vhP2HG9oD0LA8IXtU7TnRakvDFTDgUD2
3kpieqvPIrZAcGXpVSCBRXOgik/XKlc/Q3epoH8FiFoIYQPChF9AOvBwYCDcfOkE
Fy8gnepRn3VoTZCDLOIV+C7k3HaAWxxrzY7ElZaTykhYaAiyZOtmoMyS0aWGru1J
SRLGEitsWq91yRMZacHncl6a3OSoFl4yk7Qk9ckE3yV8rJBpPE/6uJnN+qyrHEIW
DaNxVRrSu178ACsPHyqhJrPjk4tpNTcuaCBMxbqxgD9ESpQFw2PigA/BcSNZt9QM
0V96HaSJwjknmoqJLZXsK07OrCZ5g7AGjARcIirtEY/FJNcWN+klRXAxg7f984It
r87o7TWfCyhn92yOZeYoYhoc0LkuKKeXLD3nGvEgp1fEKul1bGps5MNbDlO7Upl6
0pum9d49s8nEOTyS/dG7AM3knL/ZpyNuS30FH9BcoUl3/lvz2ywX74VduH5Lzq/J
a56P/CZiFrIEgUSXJzh3kUjtSDnzzyPCeWIzOYfpl81QqO0X1JAqP5H2kXLY9SQi
7emNafCyKcRVlNYflZGNQaPdxYmbeAJ+rT8uEWiIz4eVQdEC3sPC+vQ9D+c14BD5
oL1FwbVbwFvcU0X+HzH5HmYP/5xYZ5KnQjGruS8MMT+ME8EYLYtThGYlNJtVpl07
1l1Q2fmSghOUqQZ/LzXvUeBnCGMFFB9/Zi2n/xY0pvQHD/dhXBKrmcItEI+jwtDy
rUEFrrCvjkWJIc9UeiUVoXAfAmvxf8lobzI1DzITvRavHSMTVgljvf9camve0L4v
mzTGMeK9rwUOYIBsf+BMwuxO8TvOKVSmMfNYpErazjVX06T7nBmhsmu9n5s0SAOh
uCJMvdaj9GoQfMCBY9tk5T0PW5QkDlyfOEvH2qUHFiFVR8LE3aohxIa3wtJIYtga
ACMGEPp/EQbIdP9gzvYDFhiuoHVwzn2BD6ztDZrm81zF9AKZRDcSpMk7Ep9vQZI7
E9eOznaN0rquKF6lklrWOjCxO52J2AxPkw2bILvws0Tm7NVml/sdvNG7WnI0XI8A
ayd7vfIbbnG7czUaj+dqEI7geBLxR9vmGSBnL5zjVN1eWOntU0umb6aM4aq8qi7k
9D+eFjQS+qUZ/aA+UTo03OuPpahPO5MfLo7Qkb8P1+vaIjCDPzu2PK1I4YiCxVPz
VYa+bpi8NRRZH+YrNAAxKeATG59W75+LeCYlkyyWBeFYiYtNMjyLjadhCGYBbrM/
JyM7OpxOwIPW/PLdLZ4gGvrTwaCd0fBJp83it3+Wmv5LKUNJU+6EmzwK7ct2uhxR
dXJMTQogje7F9kIiDyu76f2P4N0pOevLwPAx3yUQl2QdDnD7KtLdvsUEEnhMp24y
HiCPnBC12wI1gMLH8VdsYYjuAQM9gXnam+sgv+d4Q7VoIRcjb2A0joHemNF43uc4
VfgJ4fbxrZP05xW7sS5+tAhmb9dUAn6r7wnMMEMnM+ScIK8wDdkUTkodFdDSNDdC
c1hOKDSpc5sT3AjiY5Qe1b83vmKo6zR8DwiZHL0WR6Yh8q7k7ccr7hcL8c5+/1vC
tAt2oo2kOBSGT3grEsw9eGfzO/32Mdkm0huJLmWfhxeP0pgbD9YABFtIhhmm4T9k
ZQjZd4WBftglrpW9Sf/xWUXUYW7fzOcFIYTaAA6kt0rPKi1KtnTRPuMzY4CAR4Ka
Ge/tLPS0Kv5W+Rajfvld8rqVw91Rgnf/hKXsZbbNRFcCkhvRxSwbDBLMFq3LSE7g
3RDbG8/F5p0Svj94nPa+xisUoADsTxR6wig5ZJ3G6zs376qF9LlRdYzK5mcp1xFY
QWLjFjrMHiEvyoUJ18kRzzpg2Yqs6GSHVmpI7UO6W+nl3VyBSO2T6fU1ycBcVYnW
rg5CYAgirp/7p0x0DbvXI8rrGz3nlOWfCcUBUce9UQCWpJCmBow1IQxU6DDm5U4i
vAL7nNzlASWkziWP//JuqE8G8hBm3fX/lo7zdnfEnUNrbhDW88Q7MpFpGEUep7PN
UGvyMXhk1ff5ZA4uAJu+2J8fhnFN5oPcYT0CJ7BwqAKoCk5nEPIezbTXzA0HWNmE
Afce7oYt8xMxsJkpQrAp3YOtmHzf1IM972ayFRw6bBUFYrfpOS9sqLzRO1jBg91y
8aro1dE2Da+39VbgrA6wRCAe4XdStmHOrrDa0qEa6WIdXDhNaUTkqollMX2KFkwv
Vwh8OFGzyNl09xHx3lr8icL16xmYDrcX4ggaOwI2N4kHBP1Dq6EVMyxdJkY06KPB
UWRolLNXfdnmjyBLWMWJPj78G77Icmx90v0Owr5J59OQKPe3Qj2wM6LJv0Nq/GoZ
05Y/e4aO5QVEz6sKrC+MG0XcCVigspLf69eOlQtdkkVvoEdObjJvil4zLKFVtKPJ
+8t6RQx+Er1rpOK4ssfjhCSCuPijci1LPUEj3VCN56Fs/MP13LjVC4Loo5sAMgbq
H2QTBGi52nQ7a7+64yuwrxmeX8R4lI+yN1jXdJ4Tu5j9FZKVw3ql44o8dgTuVqbv
NGpHcE69v8omCCPaSnY4C1O0bGZwZhsoetxacV9n/TS8uuiiRzTuJ280v+xWdrQu
G/mT9zlg2QbnGJRDrq5RAQ1iOVwY4i6qamXwZ8g6P0HKjfiCB9z/3Yiu2ntKtOG0
DYHCyq7ErKGX9As7n8rwgI0uLRlidOxvGI6qRTbHkm4Hs1EyVB6QSnzVWxQCV7Fv
P/wJsTF/Ex2BRaGPpxBCOmVdLfCgH2fCaal17zcWCC/ymdigtoBrp2Uq/mXTWzLQ
Tby/bmoXwaOCOxqiiWgvEU3xSZg7b1Nd1ipipsBMQYh3AwIBVGwGnNgHvWDqvLjj
Ja4MtfEpKdCM7QkCoZiiIPnrL7wvO0SJeV2kqxxRm/uuk9GDqrX/0rnbJ+Xnq0EJ
J4UJ+ZA+pyZNnxUkJxkevSbGc+CIyZMoxnq/bIsSBC+it2CtwIRccVRWvugjSwcf
DyLX8v8/LlAYp+GYbgorSzRYa8UenemjdqVzHeUqCSYEWbPV4Rme+R1eUAFQTHoL
mCwonjAd8cJkFaZ7mvblmmJf08aDsITdbHMWP8Eg70rKIGWicAVRNCBNcPbM9uEV
5dtOxXR1+bAPraXdE78fptGpTzWBtvnNWIhyPPlOTf4VkUAkJaZ/N8gtM8i2sTFK
hJq5+01Sk7Phbhn6lwJgUHe3jkhhUduvV4hldAe4NX0g5uaDygIcwiQwk6U8A1ZO
n7YfmxewEv1dgkuXUZ1UuFhoBZ5GMucf6TUrZSqEfM4Jv0y6jxo7rQvuYlY8n8my
80GWlQBPcfcFlPD8ETQf9KY6baM/bpUwF0w+1N9q2fNd+pTg8ojMu4Hs16VsT771
esSSwkA4LaG94XNtZu1+5EB/3zx7pWCW3PMXGYv7zaGc69ZriDLbIiU1Z/GfU56n
lOzaUKnAqdkMp/c9SOoRzYBDKtcIaipTgqYqOyU1Ze4RuCdyoMxZ+qKNL3IlDJf6
KhCIP0lpnpDIwktEOPrvfxfz37Ho0W2S6Nwfw8fJVDr/OQ10hqkDs9edg9UZPxu/
DxaSN5Kqd9yKEnM8uangiIQ2MxVHxVvT2CTwh/jYCF+idcwvfs3cij4cMWNC91qJ
Kwu151gx43nxJdkOyK+2wsG2FZFnOJtCAyrvyj5wR61r/suwGebqsEOtN7m6vG5Q
btx23dzPK49CvILIn9p5JwK27AnPsNIMYoYtkzGGeAvhfvHMWt09c6rKC8RttjXO
XozKDfj5pqdghOfhKkFKTKKisjJ+qRWwYpbqtWUAFKrly3VhBNw0SXCONkUDYc71
aB4i7wyL2CbwSbOk9bKaBjAt5wZHB0I656B7C2KUFNVgoR5XWEQzHNBQmZfXSAG6
XYokda4rY31tAd5TfK/y5u+OD5HvLlJdUSyg/dDIOlw+/mdifkBzXqPz6vVLDCch
V3VdpXJ3t4KseiAOSx3lKLW4k8nlzlLsJE0Hz9JhDlUzJ6FF8k1Vzlpty3hvmrm8
+qGPFGFWu5I6gtkjHYdbVQLpllfDuCsaiiGkwFHzmvf3cAllTkugJFCJwLF9xfQl
acA84UZmQWPVgjkTOIMzBMS/UFJnJVrmT1Q9bxBeuk1FcymIYg65By9TVaVKgCPv
cpriCgxpiDieFjoFAEssI+owmBkOxdte7hdwov6I4mJ3NZqHIJXEs2F88AfnQitE
IXwyu0Bsmi/QRwx95Y6x7IQ3gONNQO7P+1alKtnFTJgWhklSbbyZkos3eSKVUbs8
nxJgxBde2qdq8MKzkN7JVX/PHat/nUySsI3yT8CSUlPubtZfNuI8PJY5AejwQzrt
7AuEbKh3H1Oow9JumG7F8ZYMf+ZC7Zd8ZFBtjovUcU83x3Bnv6m2Qiy2A9s2EOTg
+zOVvE2nZBWXQBrhYNFI+9IK4dKYXRdtAQ0ukGEDfjNODVFCkPx0xpyCLnQ7bpU1
BWehwz41cYAVIKB9dI+Xv6lmqgq16AzkCULdyjwOckv2x6X41t7LWNpuKVqP1u1k
qIaPIfbPm00835CBvG3GZzLEcI2fukacIb64AYZyX4+joYYzXjutVoEgsBs9IHIu
9U91dr6mjCp9DADCCEHpZW7iiIQkZQn2HIDe5wgwh8OnXF7ZdrLxI4+BRHX9uLix
5Z5Aqf8tXaLv2IgUOPPcgYbZ5ZnrzkAfNMwTx/3uPO8ojzch/YMWp/O/Pm3jOE67
rd1bHsCR2i728PK4oXASdBNp0o1An9MoASETLh7cxs/R0pnjXzHN2qytK0y0oXpq
uGgd+Vdd04ZGeCuRYvtdVWgq/9tPzN0FdevVgSFAp+ViqwFLuMXQn/Edl1Uz9Sfn
c4ZbIgZ/hVBE6YDUtZtdS7+3S7K5KGtuJT5/DMYOTtLiHoMSa0zdV1HwwVSVPTEn
VVWzopIXv6toT1ZKLhpJgeRpNU3Naaht4pVEq8XC7a+9bvWx5N8iOQstrvgTnHSJ
G/gfPMQUFOOZX+vMAf4G64W6EiXyD150hmMXNX788Zi6RQHsw6ejWd/rf/JHISmA
NbQ7IQna2SPZQgq0/w3/fFipz8fcEPdz7+ofa0sl6POTeRkX+woix9x/Su3GZ6dx
fQNFX4eW/2r7Nx7ohazjACiIfph0vrpBPenYjQwFXbORll/Kq9SQfpz1D6XaUdkr
nquAsxYwbk1DN+zUS0UxQJvN96LYzNW/VBgdncuxeZ2dWyiEEK+/PRwtIuxbxeKa
Q50HFzXDnRwV1knys4X6vb8t2YVrDOaCQMeHNFN8+LZSQZVlAWpCZYPSro2lSW16
NPI+Ge4xtVEWiuY/dGVAjFZWLAIdRmxLquUZeB4wVvdsSCJkg2aLcHgrOwXhlVzM
qBS359yJL8A1L7UUmOgcYhuIG/4+M0Fbl+56J351uYxC/Jk8v0zRT0CS6f0EbPGJ
QVF4Fye4vTFL3PClHiGB4dEELZtl1fT0MVZU3e4IU8K+hilwnOEIqcp1+8DqN6bX
uEjkvWNFdu3dWvkjVeekaF3To9l13Y4BvyT0WlWYWWr45v7cSUVNVFBhX1ZUw2XE
lUDSIbtMkVQNO6b+YSdXfMGDVYu2PCF8/9Tl24sWmZyyfR8UEJhRAjhxYVEthZIB
dSxoUzn5nxGfVF6Z3k3XOF4hf2gEKQkR/ziJhyo2Gb3iraP5dR9I2Y1IgNAVBtD9
h0vc7Fl9QA0dHWaVcDl2Qgtz5Va916V1bIajZNbaBnm9E0P7DANczXzV9kGD6sRo
joIiqtsvrlZYomtp2sf/J/tpqkYJE7hLFtm3EnL2lQQxTgIAhk8dIzo05AoMb/E3
Gp6/gwJxvo+M7YBiIOHqOqAf3L8Z+t7VU+mqH8GEDo9GXFzRQdYTDRusFmR32VyT
xrSh7Fzawsge+himS9YfEBOq3Q5xCu9bqU5OB296Geoc3hjfuCkjdX8hLzl/m7DL
MD10luYXTUdMmPGhsEO0Dm7P4q30zZQSfFx/WqomVyYI8OUXR3NDzmXQeUa/kl4t
oV4lMYWhgPGy81uauYiNQj7qRoxc8tCsQ3zw6MuWquKZlTavqWSNb/2TdfbVB8c8
IR31+/lHHScv41COm6CiZ59K0kmw6e2GdBmEkVGB3VUrPrT5qlGDOSUrScJ4YwHc
eovVBNCsfrBJ+Iqv6w0e07hM/uhEt/jRpYeV5T5DP2P5bYIPkcm8TEBAiLGLdFnr
2C8YV9Jpn9ZBIzP7/zjmhxhwXmbsyUp2TBrNt5AN84KUFgWdx8TcKBLdXkMYXF5i
VUfaVcgAnhBBFSksuPkHCGMjiN3uxqhLZNKl6f4ZZaHcNcqVzDdYf2pPbD840U4a
8LYbG2m+y2cjIYL9eoLhiciKxBjavVU3F5zzc1KkBNpG9LdLUeoHJp7Y+hh35RMH
Sy4N8QCBLBO4u+ThuUPXuv6SJhpiZz7I1eGK0KkNugm6PjuM8FhOdoYaQ5jBA7u2
LwAOLrpq59W3HCfXSPwcUlx9UJxoTuuP4yLqdF+BOtHXUU85hnlEcLnjuoV3u/dv
vfGtG2ioiIXaGAeQE7cyh/307avDEcbkZl9E8pdO37Qr6Bp4gl0VUN65/ZVY+nhe
jley17pMB40bcs9gdW3n+pYb6M3/666im6gjFQbeyPOEhW2Zf++45BUVHsGb2BDj
QApIb/WLl95b1IqsEdKREB82E79TymyH4RT8xu2ggGQxW3yefgtVZKyGelftOoJn
oppr/1Lvb5iIZT2tCD2YNuyMcGvcrkydVeuImVxt1GrcX07uKNx2RhQEcz4LDyYd
x6WtyiuDQ6MX/ZkWEHoExkZCwZREm8CPg/hk4g9fpjHgDfSyU1Ybrpr7jqLrCl7J
uko4rEAO4+DWC/Pjoek7AdEunr7a5Zyqdv+B4bVvpDoz9+PucWxe2lIE85b+UBm+
vpciXXzzStHY7vFhp71Py/s4EZwynud7UtTIxo85rvAK45M0A2v6GEDiMMj5bZSn
9EE3x6HySme3uBLy9+aErps/5u+vf9fXgUbdXbRuGkqDElpD8jIedn711Yr79XFU
prE0yJQJehcGxaprLUed7qhjWJJ0SL3Rwsy5w/tLvaw5cjA8H72xWHj1Gmq6iViQ
CwSJZdkK6b+ePl92PHc8kHiJDL7vGXbzOs/bSUBoE760CazFfXUNE8mSfmDqy3t6
Cgm33fqkXI7Cnj1fdTXpjX7XkeoeTC4ORguLkn8aNu/WNDMxn0Jj+FXThY6Rrytt
giE2k166QsIWNCucWCS6tWWJrT7ZScEDBA4Oixvy5oQIb3iLhgs7SthqdvmHmZyd
g2/8C7u819ZLok58jK5JLWjPfoO9P/dnSwOPcwb8A2qa07DYb9Ua6KoVUOko0BuT
g+2dCHkXocDUjeKG9O5xbwZfbF0tuJo8SYAXEoBdNpXK1R3j2OvAoOQTO3R8BlNs
mkl8gZMkuigmG5ukTgH63VaJANAW/CA9+Aw+ibUWYTCQAFhgfFToKvXMn8L5/Mlu
CSTGuvXP3+49z6+wxu7Wbx1+zkoOYKI3RVYFEOu5AeTiJp9nmvb30qAnuDyu2Xm7
acShAGAVeX5mddeQfAcvDeFPBhGCINXDetW4K76qsQVBOLTTFwgSfEkhedBWh9ny
FkoKQCPfR0rNcoaJQy37ZikWDIW4Oec+cXBH5z+6yBKRIm1XIs4BZN6htJrLjz5R
y0oEw4iezar2dVcSe9bRoxq+FO043Q9oR6CDHxyWdHp4OQJNtgvocToIsKNKqqiT
j8+s/jzxiEYQdI7O+DbRRw2XdhPKmVojTu82dS8e9Lb5YbphmO4YOPpmSmYTtpK2
j/iX8S/2zuUhV8KCZ2tzK0ofuw6curAcXXio/bWn8dHk/QeodR9s8dYuKS0o6qFU
pAuQq1o6v4bovmWFI3Tw+hs2J46u11RWw4znUPya8Ej1LVgW3gN9xCK2fW4TQGXj
GY7IyXc/737VFfc9PIlUmutzjl0yq1vyZJQq+ytOXWkazQuzt68zX3hr8C9n7p+k
rSrJgczve3cohS+qHhdXlwWO4l/+RVaHOhqwFXMKX9hRGWfG5YrWoBu0+LKkOty2
omwLD/7+wW1vDxyfx9t4x+PIqx1XfSUzxQHCFIJr/gXMaCNrGKifWWq5qGpSFo8t
p/tNMcqXp63p9L+kiRpi1iYXdDd8kQnMr98unQRkDlaMe9n/78GEH7wxqhNuX5en
Ke7aVqiQg/mQ3MNsJNq/q6Iz01jxE6a9rjlePzPRUJ7kaN4jZUHbLC+sl7hTHleZ
0x2SqQlLbejHxhEGOvZTnXg2jJzX31xQZl6h+zMUKA+ZF/GiZAzpWw30qcl8m/Us
RM+2COulCvlh8NrejHBxwit2IuQtpLG3ItEbggKDRhIJ59d94f8AaQ8rjRJsKUcf
hRrXajBDEh/xjEONLpyqnF3QuOCcwWJLdpmF87r8j19Vo3FGTryDH9Nib0Wa1zh1
A7DdFVpgDh38VLEERlR/esRnKgHOQ09uFG+6C+Zo2QCO740trqoj6oAH2IbOkN9q
IjZA2rYw7/12T557OxIcmk+J/mYJaMyltvNZc304nE9wVd/GMm1lOvPambXurAjX
9kijGKtvhh6btKDH5I6NZi+JL5HlByKqqmN8lXhU1daprf7+cOgya8yDErrs3U51
6UNhoXTpBTIkIT3ePcQ0mkix1ULVxRWQIujyfVpergY8bLQx4+TOBIv33f5uOSC9
+Rls47m9f11wFMiGdv/i0GRkMQ3mAKnNuH2Sn6LV0AS8j5ieUqgWBqeOjhnGVIdG
EIpghi7YYmm10xGJ3rXxFpPbPGHX5K56m47kRKihmXkSwM4Q8utbAOOYrai2B3yZ
8UOcgiOP+PhH/8tcIXeR9eR0Y4BwZHAodXfWxtDSd97yZ3NJRmQtgxv/C+Fy2dZb
51ESalbS9klG7ec6cNxwML84hq84/rsX3d3JB2UNVfifrOqIOhMm3VaP2YqVLREb
lYs+oDBOlXglzHgMYEWTG/psFt1iPjHjMa7NZtHORdMY5kuuUFLycT+XrkcXlmSj
2pVt539Pz0041fZ6Z4AGOyBPjoWikzxf3C6bWfMFw89A4BmP8EF98BMTkbr+fo8W
VXUGrGSONsebKfGLgRFDaJWNVMHZKkfpBe9qOW6Im1oJZL/O5nEl+9PNcog3l7T1
ZnTJQ5W2hwPqZJ2z6HOzV1kvIsu1mPo/AxKDoXYy6bdJVxKtsC6aDpWBxeCj9FaH
lkwl3rKh3lNOcvLlwaXaTEOyyv6ov+PYNyQW1b0VVYlpciG8HdnROhlYOB73a62V
JsOGrbhEpHJo9fleFYm8TT1C0ukzImdgXgbAntf+a0dR348fiIkZ/5s5iGjORQgK
JSFC+P3nRdehaW8oo0cupjam/BiGlSCskluekGRD4NLxmLxStWzkW4uhyHlb5TkH
M+TXdiNDQ3boeH0rVFLkziJIPynPvBwm9NmYj53KwXqSh+Bsfkd67ZL2e85DFbq0
1s3xKrsWgIRVgGmHsLDOZF7r1lnqXpMOXNSunFwz9+4Mpa+AIN0Wp8Ps1RqYmMHf
lxFyxWQ+RduJtsokYKxc1i8TCFtFz8++cmgsDLCXGVueaufZ2r73+Xstq1sew0Dd
D+ms7SR3blK8s37jCBgx+XtYg3bCajmUEUHTBJoC9PP6zxXGgfvhPaIbZAuU4YMg
Kwvx2d6J9hSsyKg76qeNc95JD3ylAdBKfKHpc18ccp3yxatQ1iHr2fRzmyy7T9wp
agtpvOmJq+gI2d96mbF8JMtdZ2DN0HeXiioti2yy2ePm8STt+GQW8umYBx4CTOVf
lJYaDZqbbmgvgyQPO9C6/jXWFAN7Vl+rUMRKcS4FOTYnl/AGpPZ411hTAVXqQ8kt
9TiZynHmhFtwhpIQX4kNZjVe4KkxajBBk8U1gW39QpuKWB/Tk+ZDElZGA65S/SSf
/ZII83IexDDUsuP73QMVqU/OyVoiyMVB8B9A9brRdvEpkJGw3Ysu7q3uU30SZTtA
W+cQXWoYrMGAsKV0eUfN9KTZCHFMWLrq8U3n4cG6wg6/HxOzdpCc8abmk1bTjvT5
rnmmDVM4iJVOTX4MYebb0trfLGIoTJ51XyLOTNBloUlrzDReltd5sER9OWehrqgh
t+RQlAE1lBwdAjlCEWJ9JdBU4T6ApgIvZAJ8lok2LWqnWOhDuhjONIYfZpJEA5iF
5yLCYafuUzVJGZEJDJRa5aaA3ienwI7WX40qtnyRthQgXnDQTPPid4BY8B0oKFcF
jmA6Gfodua+LKug9yriP+DviHB/PWCEwGUdlkeKEfQI4Qh48T4mtiIJRWg590KYo
dgyHAn0X6xdLBk3UIpb9rI63AaH94eO3U+eNhxh3do60DTQST9tu1vHQQw0L5Wpt
lUD4bUes+9ZSbsyLJaYemaCC9heeV0x8vCtDhts05i+Lx8Dzjmrl4V8pQ1Kmha1s
HAUfXl2BOcKnoyJKFKT6JHAns8G95CkYB0otvxEZenmadUYSMdRjj4jb1DGSs2LJ
qWKdIlHAgxVOek6bUV6rcGCrKFZAeWeWr4qT3Xxdb9eODX/dwhmQe6OXG6b3Cyr8
jjtPb3XMGk202dpS7Ia5Inp5Mn4f1HFzz4c2iJ4h6Kml5YXzUxuxzD4pMiyJLo5h
+bZXzkqf51s6uw1vRZAtJefabiUlK18tRzk+DqJIlAt/NBM1eWFl9XvFzGKcTCWY
yVNd2/umaHpXcG7fsEmy3kBxoICjkjp2XRuido7wxT7AH1Qyg72to8KqQ/zXhx3f
PNtBtPtYi0ZcsNJQ/DEh6YwQcBfKa1qjhEgp9tW7GvpCoWxpKChMwJHec0I+wKIy
ZOIrtvmziRj2ftjAusBZ8x6XsT1DpPNCvY66O7ZUuOAcOuE1j5WmDNTPwMHYzrO9
v5jAedHPrp/Es6VH6peTbeZMkXVlaNPN1s5qsaJ5D1MBpfXRlrTvbU0rXgrjtkB1
5DTs5pag7KwwBoCnrFb8jK4uKOqMyBYkGOLx/Gnck1EmnoqVLBXaefOl0LePnoRd
9FYNjBUT7qQJHPX4amZ+Io9N7f7B0i6bP+FsANdgIbelDc32fVmM8wZrioMkioJL
Le3Zxp18aiBv+vwLk+yTG1i63yjMswqCXpNX+Vsovd82CQvMCVD6nDxr6b/G5CzN
FhnduNS7NnfV+yTde1oAMK8sWv81HFm88PcMViq0FpW15XNOdQ4HkO1auK/NR/AQ
w1GhiFfFeVPJsuHUVLaRxJ2GaHBp6NQ7O6P6hA+Yg68Sysm3nmf3kTLIe9qKqZGG
ar68cGxf8eeYBKjbwH/Jx8pAicnm69PUrvZDzgrXOPAwiKwpw9fyTHMtZtQa1Be/
oKnrLJZYkblpEQ/jpLJbaCGB5xzdPJXqxT1EYpK647qfP7viP28EDZz30PrO2s+j
BQ/kBYBwbHgaS6TPZNgFJaHj6nhw6laq3xLC614LhVh6q8XdqMO7attF+HYtyC2p
6LDkwxCQoOnw+4ubvCKgwNtn7lk1fyzT0b/aXzqPJHFaQ6u5asvjbddNgqk8giIo
Cujxchyjx5QU8HRyUNX8B15UwOi4juwMpc3jggXboIxphHIL671q8f5gX43TNqjU
kgr4Ff8Z5V2jwIuAkvyUkCOQZ8DhcmRPhk50JtkljcnZQ977GbBG+BlKGl01HH2J
2O+IRTgdukBp+iE4/LRm1LFyuYYZFDHn4FovtjCFfR1WqNEOCe8FnaeG1r226S/L
/onVFBBoZ5+zUFd4hoQNsidKf6p6sRyeUZfFnksp7OmOpp6HPvFdG/3bML/l98zT
MtBgQHbgfqi1leQds/ZL6qqCjgDg3WnwzYG9Ok319LiuxV65WQKEoNstzGobUYpq
FwXd0xQXqaFt0F6s8oKvlz8Y+q+1EGk7h74Cx3k0bZWaPS8n0ErgoeY7xgohe4EJ
L6cGKW6v9zNfvWDzmyLNArkunhOOYw7a2+/WLnQT08Aw0iCxL9qqpPeyUrydx/qV
0RGL8KwrE1mkGTAcfIzHoXCcdj28uboCDx86STa9ugutjtXuTIvEvqQTOdH1xHC3
eFjI1S7SN9qz7Cck4ZyybuctwjabfOceF092twJaR5/nzHquz/OC8m/3fTvG0RVj
beOn36r/6Wsf9xhStuIvezuyfxIL0d9A0MfaBPqLl8ywJknIL66OEj/wIM4ficxR
sUmeZqhWmmNh2zkppQCIQlL9sguF0e+4K+cZxEAhyXY3WItyfdcjdbEZ9DgqvN8z
AE4Q85S1kyCOEKR2W763ph508S3XnZSlfpE4rn+qlYnUNdVY4CoERcDNZDec8UbA
oreEoTXen92oz9ieHwQsY5ftqPykkCXuigJHuQps5TRs7VjhOWtT7L4UiqAD9FCF
7sWN+S1mMMMSQvBk5CLTxYpVRazBinQGsicr0m9d9zul3c9Kg1RF9pte2GxOO2RS
YU9qMnqN1U5ty6LFczrTDI8SFRV6u9D8znu2yBt8B4kp3r/92ZaazAsvY/FTK48e
pwJpL+piVhDz4GE2+CL09Z+eUurh7NE1oWJbMDvcMWcUaIDCc9qW38/bjfY8/nPf
3uwXgBm2TwD+9vvxsLd4IEK6GdZF6zIsn5Cpd3OJ3dssv8x2vK3+CjS+/U/6WONA
CdWb8uLlJm22EQk/ENArKBbb+sUP8s4m1qiXkzWZqYmLV6Z4x3LYhCJez7H3NtyR
RpPE/5VVk3CPyiD+nFlf0GD3mL9D9tNUt6uDvfdCHqunV4cBZ0igTktAeK8LIT1v
k3/v768lmPO3zWhYjCbmJmZC+DFY+ar6Vj/w6PcqkVRtHgTY4LDptJLJ5Xhtrkbq
e/MnIEVXs8j3rm0jUhmj/DoaBNz3HC5Nj98OjwccBuVQhXazullAtk6S3Bk7IzYa
Ujb+nj0YR60PdHwcYd+ABUyT6e+JppQgPypsSdvS5/zOhVYTMhqpBC3wlRYEufnc
4ol7ymMvDF/fn7wqIA0cc4cjr1LNNXVXb6AMcGry7lBXrJ3k1TLnblOtRQtFpDFv
uHfqWR+RfG7Vt1JPsbafnziPGf2fjeWQNRbop13JqC8DeDoBuGVe5oaAe6Gg3kr/
wd0mnPMaU86f7gTNyU9TI5Ol/sJ10o2/O+jF9Lnc2YC876EbEyNGNnWYMCprwK2+
WIEz2zgLsbDw5RmBj4oDmp0u3v9NB97/iPRxf8wM80TuQFhKnJfFfzJa6ajY/iRD
ZuAMqfdaP6bwhmsKIIRSwppvOv0HEitqw6+++PlFq5hD8OAq2Yw3WPHXin8ct9Hk
+s9J9Ho6uySD5L3yidoFtVhz4oG54PWuFH7KgOdlNXt4J+8EX1GM/RRrcUvsY0dV
rawLISJkVZ/Z2SgMJsAikO6/nPA3wgMcg5jS/EW4VEOESrmbb3RQ75AUZ9b902/y
T5MjvRRUgchiAiXwoMsj26h+lcDblQFUAg9G0W2f2LurpfniXMB+XT8um/t/l8P0
laMGRsf/L/mfVuv1iFRY19adC2cxbkhIgFzx+r1T9t375xLFQUPFmTL4yozZ3hhe
7xG6ZoREze8JP1jpuuM7+Kg4Q6YNasZz5wBlLpVJ6EGIxivCT34SE8zk12fjZOlp
yyj8LaTm6R6QRVSR5mUGsDThTVt4NzIwEk+f+HjlxOBEKWD6haO2KClwefKi6NN9
/5RPKuXFAjty3qMSinafmvl1t4Uw10eKfcaqDIzjuLbLOIat7R3WwTIhY3+PkaKf
VQySrF6MDfYLhFDBlhFctXCdsvz1UPe6cn6I92ObARAHMe6pKxrpJvQS8whxtCxR
sj6Xh0Rg8czViGxiCLcJ4BPiWn+DHp8hHid7fxR0ya+AMhb+KVgHIjenSCTt4+6P
BqL+DmWEGgqtuc31tHjkZMUXumfXBACvupXXBubGmc4oCo8lL9WSB04jB8HN6wSZ
rrgtss48X6jwkkulkeB5Hl5RMjLRlnwvvadUAm2A4zcYH0QRggErTE5JHnz5N60R
XZV4quXprbs/w2zsCgLsqoENvo0Z8wWv2OKpCeOEZd+9KwOVVbFb9aneDMBbQ0kF
3htrT66Y4V9W/uy1AuLlWGRZ5CCFtKTyMrBjuY5ANKO8gz5GqMt4aFcLyCd3zMkH
diG3ii1X2vbZKgMmA5MLlupR0RwTJmqYfA4+0z++RxTFxB7INHgi8RpWo2nH1JVR
+57UuQHBYf5efsbvzqeCDOsNcY12a1p3RiYRv0yg8OTGSEMxOevqAn1wBl4WGM8H
5BLlXK1teqsf51GSfONkHfz5Y/L568K6y/rsnYHrrgXCfkYU8KYbRTN6iGoOx2XA
39jKQ2gFnlEUQ7nB9Z46SmOi49/+5Vgydi/JFqf4mejSpnaSTS0PTilnhKwcTSl/
mUdV6jWv5MGERgMyvYMGZ2uDbZ8vjQ3rOL3xe3PSUDty5RLIRQamoMVLH1E8SzWl
r4bIK34Uk+nt2u6AhngWw2FSwAdWIlX0C43+nPR6sToOLMtnbn4B1RH4ywppJCLA
cSEPkoqcWhlWkDqsUos12KJ40K/Ymvt8TMCFJyBqEtfetu+pzmo75fwYItmXWt6A
7W6EBGf1hlX4e+z6JuI7bYbeaHNM7IqfBTa2UkhuI0zpj/xuc/LDM+osQbp4wlg+
xRZG/h6n3AXKqvVlhYWWOb4t0Sd39JENX3ng6dd30VBPXgZlLXBI6KYW0Y/2w8mf
J8SbPVJRh5u3DeqxS5WXcYKZEtc2L+0WM3HAno02JMyI3gpgEKad8cS8qoZBgxgV
i4tR5NSGEK/S4D57eTq72xJ44+xr2cad9FEfvWdLh8/ec/moHsZMH5uGgqgxFpbV
99QLAhwC9HsRwLGqltTrU6KdtK8yDs9ShRh7JVQfn7xY13M4rOSEGKJANcKJr8rA
eGHM6Fa1GL0yeqFF9kLHrZ40uwUa5o/Xr7nSsi8mhkX7csNXVVmLwTpj/Ep06nQ2
OKCgWl+piVQfQYaVL17nCgsOsBJ8btbxWSYpFBubfY9d0OGvh1t9r28UF+5kFoNa
mvPZVE5SQxpkUw1bflu+MAMfJ4OVGzEupPrXsixqfy2rPouBNSs7YaLuQXnPqbz2
mROeM9qAgtgQyLQXC+kb75K7JeaFBhGA5dG1W6UIL6YzcEmdjJC6RX+eUkhZvYRS
BQWUhdWjoWAPfl5/azskIhsX5GvjzI3oRfPntYrsj5anHFhF8C70cA7Hy8eRoqxV
/VxQf52S/32jTmPNsrd6UAXObxZOgitcAIbZKeSWaKlPnoqlZR57tm3bEjFjCtUM
XIQi7XKnuCw1edu1VYLkHjZViJQac4PRmxVthue0eF6yhZIshhsf1xW4SBT5YNAU
M5xg+aJeiknRyMELg1tVUoozaZ8hkG3qLARsUsGpRdwggC4gNitoeeUasB31p5/D
BnAzNXbOEWoa/ViinQv7OEsBI2KDC6ZJU8BcyPdEe30w6I/mBFNaXhTZRjEEscde
xexC7ofdV21wrXy2lU/lXVvkSj+NNLLc/4hip68vBBGmh47KSkeTQvF4BNVhCFSB
/shXaGHyFoP6sWS612UGT2uFBzEc/PMUnS69wbxpZfKrfALqUf+S8noGnMewaXvx
jntKQOZQR8IAOUsG2r8SVwPsywUu7O08TkOSejDPQ/PknARuIXusXfoBMkcILVP7
T0Frdp7FLk4kQJqckVOXPTgg2sRktJ5fdCjuYxJg31It7RN4ToML+ILBRy8ISaHw
KJn/rxHo2sGkPSk/6ziPvW4b1fSyK7khMSK1th+ZkLGZrXnGrW6YyZcNmoi1tuL1
uYkogpUKS1MTAVLHRsR5HigGYEbXNWd/UVbdeQF6f3hECbU+hawN21nRnlkiwcJD
Cgmrq51kP+6qIzM2PUXGWpGEG4o5lhZqhMfNUbcb1chnkG4SGNoYPDXPhC5203Ov
BoBxEhVwNqTkZZXARUMHZ00MMbt8iNA9Pz+pBAfQ8spIve8vRpqWuXySPzU/Yu2f
X2GkrJC4Lw1bOWbZkt6lrOTk82y7g8wR9+EFbQ8WvQk4E091X3PsaLkLa/nbkAzQ
I/9ix4KIw+aSjbQQstiMxLyoJkZAm+f93ZjyX/srIkEB1SRG106rub/IgRBViZwe
IPzcX8FD4WZcGm7U6jvhyQXq4Z421EoP+FYggPADDEZtdqA+wrkPGFzuZOmno7+g
fOuFNATM3iIn4aZ75F85OWtWzCPxZMCYzUyLWn3hzdgfPQboRx+LXPpXMn+7ByCV
yX6cehmdp58RAk1kLYlxWb+zpdORz0NXc+MIdKLlCnzVNVvPHpDO9IFQIBd39Gy3
3fmtWP4XhmljXhzndjBNAmi+4UlppKB5Ir0Lb+fprCmfO+nd4SdDQYijx9VsnGUb
x1PNxLre3030kLHTBkLZzPEAM2p0j/uRGzZcUmMlljX3R9pSYSNRTvUj10j5/O54
PfCszxfQ9oMFfng++sehLVQGk5wgM7D0CwbBuneW1SdiEyJ86kTs/NmcztwGhh3B
b4QFb4C6fapn+aro+kwVAZrwg4DPjvubnyThXsduxoGwrKLKAvmYZWsJ7WtCXUmC
pm7PxwEE0qOOGdgQnMMSgARIxAP9DVQrnpn7X2sxMz40U8OLAbKNtgHgEDkeNqK5
Uc7kV0MZN0x4Nn2HQaNqow0KDVBr+W3BzBI7TyeV2sFwy2GRxSDzLdTPFG0lhfNn
0tdencv5fBbasIhKwsqo6cFxjzxKYRAATcG3PxHCjDL5Vjz2Pv4I0pkB1wsk87fd
99vxDQRbwusbMWJ9sNASnpaN0vvBn7F8oidv8BvWMZMMTfrag9yGJKyD2Ga+amPY
h5qGwGfx8V5C4RO1mZcX+q4VdfbznvT4O8i70tG2XZT7l5oUvz3i8w5p/x4Fbqqt
TpB9w9hdw/W2SgD00cVsQaR4tf79MwqgIs5VYdqndZRcXcVBeRPLXGqwrBFI4Ib/
2uU66Zxa0e/nulYRGGu5nc+qAQMmPyzWI/iiY5giAAeT72GxnQcOTzfKOUtIkitj
QZoQk+AbbL+uZ5E2Tc/fdiv2AMOU0gWkXgaHNSxMixmY3/SuySTPS+54awjk6fej
8IGeMe7qrYqJSAF1ex98LISNkn9laKbRU4+6S2bPfgirKhImmzc8QFjiSSatZMfC
0TM5gR5uLU2EPgtukKFeT8pz6mcr9tTihT7uR/Ls1JDKHmSoZ4skWcC9GrodnsSx
N+6rULkRM7SnLNaGDs3pjKHBpcMlcfCWU6JTPB9FL8GBNnhM2Q9X/NCkV9NCvN+C
w8Ujx4gtJ1xna1GGmGccxgXu9jAtDWYVKur11LempC+4LObaqVGtn8qYVJkcWsap
Ub0hOeT7s9yPBMVNOFWvub7ZvnflPATwucMcerujYkx8a1V2Lb2WKGYt2KfDcjlp
FpfM7eWHPZX/4sCNTUV1Y/zp6IVru9GPdHu0M5CLXFbDcJnNIUy0q5aKxZ4zgK/p
twK6LWC1Z8sMo1V4ektZ7g5GvMXTZ0b8JSNQF019NJ9taNvAvpyKchMPcq86CPOj
rImJIlpt+1xTpqm/urVOLHzqeiGzZPzYZY8MvA7QqKpNUU9J55DZ69sGo1EIY9ik
hQuwdv/wCqTKYJ6qGb+HgWhMu2Bhgw2a2JUV6atdj2r4JV06k0xcugk0LVnO+kch
3l8QofuGHuBx81JT/qG3i0ybR7NpEo445suVKlNDwjghWMreG24Bgee7nbehdtpu
FvqnM3ihcF8K/nhRXgJ3lcp7chfqsTndWHSCRpTCr/wjIsLqNRBI5neqHUHdJPZh
EB/dByp5M8tFEZojDsE7volejC7GkDWnSB8dEaxNEa9QtxBV+xiWAz0jP7An2XaR
4TDk3gJEVWPd0n7k3iAIGT39sFbfUi+9NMw6ZfMSwsg/AUs6j6qytD7lO0eN0eqW
Guxy3qMzOo1Op/MykjX7iW8NYH9xDylnNrhdOTrObCcZ4rgycNPJHinx6M1s5rlE
LjeGA4QEtpnYL6yQlXqDHtUPeZURudq4i4+6Ky9nDx843yCTUONbTZecICZXj5X3
TZz2R2xPSH1qcRaVr2Oupb+P0AFeq0vfLodKGQ5pcb7OTpn5g1woEetkf1KW3yka
FXKDqdgbLe9+5vRBFF3/GYy6hxKkFOowADOVK+2NFdTUCBXBh4HdFDSZeamIKU8x
9v/onmvQxRPGektpclvF+Wr5cpCLvsciwVnqp4V0TGqFFO9bIkQJVm4RxOBhNHC4
j3jpEKbdrLV2Urb95+GFWtfRIZ0OW4yz48kss5JOm5weVImUXWTVO68db/kLSOKP
26diXVwtvI4WOD/GAS6IsOuBS5WH6LLwM0HNfZltLWnUwLUCO75zf1HXg7MqHshx
j4FkgicHYpJ6ohx2LbAzUOWEBc4oiDUrle1sUY9QP9G170YCzV8Abj5o4Y+fvP/l
ex3ds8KuNDruBkOpIWAzHMt13pIJ6+fKGKEaGwkCF4T+YRKr96JQRsqSYwyhANbG
KP/Jkkeme9g7BiWSjDnLOWWNFVLZYrx6kTBGULHA9DLnJFw73eHuWZEbUIzr/TXP
UqcxnXbp8nDDR8JaC9Q/zWS9OeLzYSuYFHuR+z92J/v3Zd1Wpnx3m9JSd3n0xR0d
eSiO7TrXsl8f2rBQbuE/w6bDY441j9jEGYlPsd7eVLM9O6yWZA+S2Pu/1tWKWCuW
gucrbh5/PIGkSG+lHMXHR/RmbMQCugzogcOMFor73zOM2q/653RkTKDVO1Si1E2+
7OaaO5XTaICOwBAU/n1hlR9wathYVT3SRUqMB2gY5yLUwvNoAwWKIN3jAiHAc8yw
fh3h+eQwWDeNs4HOX5EPo+lyvFhiroKvCzxesTupFEpN9Uxd4d2xSjRY7QhoW98E
ZQxxVMI9T/HUv6TjiBIebQhJXy4hOgmqgroPU1hF+9sK2Kiz+ehAerd2m1CN+RPt
HU5nqclQOaY5r/uK/Sw23X2Zm7P05zDT1QjAV3W6e9vqyfMdi/R9nKpkIu0WEShE
GVCVF9ONI4kkVloPqSRWWuglD2rEA0hNBR0q+I+LdE7hLH020PlESKyzU6fbqTxo
oqYYDUnuFlDfmyKEac0x7RgFjIp7Y/czPgHc3OdPmzGWc3WfMoO8kJi77kW+YFnK
WEJslTmFTBWsWHljsWSBEJoNhKX7lJj8E9O9u8GJ0HFvkPXwptRbhR1EIAul+M4z
OJkj3VPdOB8QWg7iG8T6+mKiXmypA5o0osRxEkboZlil7cpsliyRwR9JTkUIQMEk
pKi93OS25z0zBHQGvW+VSc/PZtvVt7gUty3ZbAch80DSj0aqO6Tzdti3qHRidMcb
PchcwqoYfablfDeWMW09e/bSs5k3aEUkS75h6Pbp4ixPC5L8oR52AMTEU95BrvWC
KWOaSBq7uk+tLdBooetCvQu78mmBw7kmXv88io49HpOAVgavT7w0ayXCJBuUS+rO
SJf2gbQK2WvP3A1iMZ0z1WNtZYItnxpNJBJVRSELWvSgn3XRBBmXjJpmWEW4Grvo
+enT+Mm2Z5JtflXsDxZSP1u8F9XWRC6SL1EejiSaDfQfGocJKcIqg0xfVL+dK76u
ylGtlNLM45Ywl49ZgYt2J6+0Tzd/Ctj7mIOEb5Q1EkGYaZQfdOj0CsviI4G2JCtq
+K7e9/MRCwm95xekFsCl506NkRLZEC/ph6IQMLWw7e7lOKgwKhCsTAmGdX0ozUhL
SR0QCYmp1t4A+oMXLKUc63Ttu2J81sJrWO5aYvh0GbN5gNHcVW23S71q6a4WXTLN
10+JeR8VIsibk3oGUbVHJH9KfKIuiPb4Fja+wGjNV4ffLbcgTn3Vdkzhg9vT1Mj9
wXWUPkBiFlJDenfDsO7Y4F18hME/04WNIU9znvaoFqwkF4Nf/ndcm6N4mDrUJ3hu
z3fTQquS5lYvpwejYH5mLTBA107EiaBaFxZl+mzjee+hkYaAhqE/ccAQf7kBQrRj
XqEfiXyynQn2Z5K7I3oB0OFYIhsFO6nvXTZQInPBTTXRffBaLPaIProw4wKFKqr5
o0TDqjXjuZXgWfq8U035P5i1l1PLGkMqlwMMGs8eO23yVqOFe+S9nkfkt9Vl9/qL
/hxvtMmSx8i/P04U4CAJfTPsGODmmt7R7shIuiOLxDReVpOIYc/7QunUA1pFB7zd
upAI080qIYqv5OmRlprl6G2IbkrwBECHNjCrrJU3+1bx1GpO2iTpU8iENEmxrYRF
Z88YlcKUgk1pMhbM2W7jfjJFuEcSZK3H08Of3WjZM1vcSeoV3EpUZ+Et1obQsq9r
/8Y3rz1L3SCLi+vtC/a7OFDm0/29+tj1v7ta1w97OGzKYTc8V0aiEf9Rx2egzelI
iQTy/sosSmgtqtxVtr+vznHu4UK2boTj4IY4TzJmWVVNGZHRVy38oIGl8pcNXrBd
dDs0lzjIwpTDfJfS+T/DvJTlVtgosO+uOzjf/vvKf6i9qXeHjHopaLFyGwzs89JW
MV7+3ANP2saZB55I5Kwaq9IoiXb+TO1UtBS1rb3PeYiyAKQos8RV+8SzFzNkZ64V
ud2RC3+gkjKfbkTADqe34suB3JLtdzRigrWIdecTPLZt62g8ou9Xxq+lYpsDoq20
dWKYgC2JlPPtQpS0W6ovP/ipQ524fRJ9Fq5YOkdV7k6cbDcjW9Paz2MH6bw7mFyw
Y/gLDJGHb7xeEV1amQ2X7i6eJ5F1YsJxrGJVTWHLY1KK+6l7SIRFZCR55NdnYwrj
e2N8bhAHuq1bzN9q689IV0acLUZ4tF+s9ObL+emt1cuUpTU65IQ/coDDsahizYFM
48986cAYL5IF97TyyqWC/LN2Ddczhr6s2AZvg2Ez+ggGpctwpuv4x0cN3NP476Ct
NAnOZDAXH7Zw0xxv8Iexy1pkGOdxY6UOF91pi3MgmcwatP+x+g3XwZsUgJRxOIAj
pULr4r3O9+P2yRq9ZdG0p1TU7uJM7jn6WlW3h210AsEjBO2kj0lNfQR4NBaqQjJd
xIq/HAztTwAMZh568ICZhFbI0Wt+m0EaHM+BvvPUh7FERJFPoFDEiRUGw+AM6Lcp
cXD10LzYmMIxs8gDEvNS+7EknfzeYd7FEaMFw29YO2pMprjNC0PsgLmJH0RXE2R2
Gj9IC55GiBDEnOurbr8eajfWqwDVxqvBS34VEOSIDOZNzg3CRdsOWW4kYSI9KbYJ
uz0jMFiX75OVDNfNHSRAXrqJRqe3tHIWzXxBm4pmeMloVXxyc/Rtlv1SfgfHi2Q8
ad1DPtkQCxdh97/t77sD9zSogoi7vQfFnVk7ACuTkIUW9+lUbGYTmz82gBIpAlUJ
pfuXJ9OeDlVCzZF8oUikeuSJxzfxGom22mw/YYsSKcY1EMqz75sabSjC1V5NiIYN
rZ96S7zt0VenDlCA5g+JS/2AqKFbfLmrAXMiB7l0V6TDjuBVxH2LO+n/rg61FtYP
ShmoyfmvyfeWogfFvkbukNcwBAuFcEL9HA3Vo3QkIj9U+pL146qvZm+AO4ySc7Kn
KmbEvaWogOz4U6UY+9asF9RSlJytI6wqWr0pvpV1DIac2lcNMQhOubazDQ6mGgJf
2eFD+GRt/9Y+Q39xlIysopgHxVqC6G+G/rBKGdsUQ4wXhyb81Z9MFx0jFh2uxdzc
H6wJqt66uvDtf5qL+cJe7CXTD4XOoxLKaiQ1KoJX5NLWXkVVvrU+R9CA+bH8FPCP
DBaSrGJuLlcmfhzWqBYNHIDm4kyg9pXVbVJv9opSup2fRDlw5tj4opyBdhgOfSl6
G1W//B0IVG/7rYzuaOeQHa9IfxWWCDYMR/0sgoxl67tbwcuHlscmZzKtlkbGb9UV
eUdPE4mZh85dY1esLfi1qfuei9sCprR/71BePjMx/7ziQHKCaVaYPldY5eSLrrM6
SNpngKNKqRMi82a6g7oPeMJYO9MrvgSS6d5Z+4nUIAZhDgY5+w5E17uWNLhuUTOe
e5/6xv5O8rlDa1nLLN7VggVznaFQCa7WbOEA8cQUJC/PmQOmuDyTAMpepnqNoES+
TG6U8QMh8U6ypojhqyACcU6yUWIlCZae7CVexX24gUSjuKVWcsl+XqK08GZgtyHx
BGxU0LTP8AUrjX/Vgtja+e5X7qovo9fKvkkBUVV0LZk+4/SQkTHNKqXFtFHZJIDV
zgvbITmSgYfFDMVzhvNFhURn5QkOQO2ADK0iU1xlbToMJmEJtqKLbaZWGXjxZ4xJ
p8FEg9rHo57jIsCmz+5vyxmTiYuqSmkt8TWOusLW06w3qRDmpfqIzBMMxJ3vhh+8
EHpsP5fbzq2aX1Gz1ym+nPz+NxIP7+klRYKyt5wCuurjY3FnSzJwXjkr0+V7kA/I
4w2KK72lyECI+NOpQkQZNVfMr1tG026p+eU85MCF9QUCW58CALy9bM2LDRmPQK3N
wH3mjvRcV5O++nGlC/jDuAaZFGfcegZsv5x3QZO6k9tCqPvnEvBJ3CcjMQOGYU3T
xfIOAfV5Q0npiKixlAfiThuaZ2RnyIYTBVKBNLBcIS0EamyfUQMvXne7zQu3LjAY
v3rmDoNHxI0wT7Qut6zMxHhfoiaOUPQ2UvOjK1Fj5SItLQpJHF7gqs4l2FcV0JYk
9ripDKli+dYCpwXAIfHcJWRgczpUJTjSPNZdySDk34BF5kYdC8ZnL3ltOt6gPBWz
KtcHy1wj12Qv0lTIO9PYtwIcYGBW4eFrTpQzpofgeMe+3BSbgXJ6JQTCboXLreOy
D9duKsupZ/AepcKsp1j9gIabfUbChkWc7WsqtUvmFVCp9PV1txl43IroJJ9IGJep
Ww8llB83nipTGwlvhIjyuhNcQNsXbCvxAwv1m2AbsIkIXGpyXpLnkaIAdqf/1oxb
yxgrwyx5fs0PRadfLKxkO+cdYACWCW0j4vdH/BE9JTM0aXkL5ZCTWWBKnlXEZRHy
KB6X/WbIWaT6TO4M1oulm/5agvsG9814ZPjj68rkUTvWdC9KhzfC38o6g7CT/iGc
o2YtVtPshQ9J1phT01TYhMuLgCLgL86pq8M4NhBuen6N9sIWQeO1rSDytoF+lPEN
3mEwfxZ0HBAxEUC76nbTw/eBQIv84jlKkIv3VwAlOtbpuj8s5GIF+ExdTm/HOsTl
Gk4O4SAthWGCkui4h5JbAp8pkRThLyfhTDsGsRjTGzlK5FTjWiD+XOiLd9IXQdum
KY6iS+zNz9AxSC5Nwo91reZEKR+uG8qsunf9kXbrVp1wASOTZaVWIn1nUODfeZfl
Nnvj3EwGxyJQgR7qYw2qG+i1G8anZerRJqC+qhCYc25NaTDiEQ1EAhey3GajaO+v
6ZliVXspLm7XgBHwspnMmgxUOGOgc04OeH4QlislvwODzc2OVPHaZeQ8aX0bKBfh
RnDying0jI1ma+zc03R0mKS41cETFruHSsDS38Ib7xpa/eaj7zF88Eb8eQ9ya2rj
br1T8+DTkn+jPv3TxVl0pUE4NK8tUI3LV0F2gGTL0QqoFQpfICc1KyxzM0O6QLGD
S/EEvpFl9CKgs6iPgFQz7C/GMQMto1pf0kJEv8ioMSOlAqtMk/0W4qY+5QzmQrms
5ZdE9nbGVf87KLyZ56hysddedS+z2Qvi9vPay7MOotbz+Q+TangpXYuCToLeRscf
VOicJXTHBXxxwszHvShTDWRW8jUeCvpkgtyBW7FKKhuSdozuLL5zAD0dnWlVeVB5
HAxosD9/RN4XDBpIFDzsH92c1nIKXwSDLnTMVGU2kdIuuoWpDVucTmMmpqm+OoYI
1b4YrKcnjl3NH7j1SGX0dC0Lb7kNHKKIDaCFNOxgjBP+Iri+Nl4E3hIkEr+PKDYb
diZjr830SOowecOa+zeT9i84M6syqVqDBn1XQhOmA/rYOk6Si7+pqIFuExSz1ypl
GJ4eT3mAiEWCzzv5213bXZmloNJ1Z8MIzS5ov44kxN85YGFBiEmAGpVMf2rMjmWs
KgS6yn2lGKaQ5TYEzrMwlGed2FSW9sQaPjcAwqo4tdhrL/64HmRlsdcsoF/rgyBS
LVblPBCkoQaEMcYwz36OQFUUZmoTjUIP00pSihu2t1dE3AVesKaQtFwXDmor+KJd
En4w8bTKfBKkkkj20AqkA8bEcwHdwUlGDnoe9CMGOEkyQBpj987+rzD+ZBmEP548
IHzt7BKYH14hP3rSr8TkyRZGifko7yfWPA304aMK+bFM69XHDswovK75EyUa3u7s
zWCXprngzPeKQKUMsBTesRRtVyc2zeXTwhQT09fVOfh2C7HcwdpDxF8Iwnvl2Sgq
hjp06nt9rB1DvXFxf1LKBS6lEXEuC2W0DIgnUD+AIIamY22xoK/NlYBvdehuy7Hx
+5XU/l+AfZKCV/lP6CHv8M8jRj6UPjEH94Rl8DHyj3ZUD73ZyX0Opx88Z2FXR5m8
wHfqUdlWRuvHWupJmrNi17j4Edi3Ex5chbGwfPUd1J3yAzxCW8IkrChe4WIp6piR
6LS14jlBXWE9E/GGwLgWBvpwxzuFFMd3QcSsKCjmBzq/le36Mv/WaNDv5vOCvxYC
q5sqXe5QS/B91nFNw5iWCBj1eIOQemSuOF+RbyrqctXige5m/KQQQ8FBnEq/6VYM
C6d9Wj3OYnZKLtl4f5tQt6fXKErGfC2cWtG6iWwnLFjY30gYY3IejWpbQoSkamr0
Zv+KpUE25EB6C4SNN/1aJFTFllqgGQXrnR2Hwgb58lEXQrjiNyUwpbICmEw+UYHR
yWXs/xzHCMTugt8gUJtm1y/T8MHqfn2D5FiwvoyfzpWiTFGPca4J84ejcdYZ6HTn
VvZXyGA6AoNWo7VauvlyfVWNMiulysX2zm/dg5Qh71d5ENAQKlSS+1JTWjsbnoe6
9Uw0yzrynYRcspFjC0da3lx8g9R06Z7zSXMiPPc5nZQcLJgCleT1usmtyevH+tyq
dRjKTBCchrxgVWCIElFCbnDx4uSsVzYkJEYC0xdkmeK4QaCyoRP1uJ7jxGL0kPwn
3UcZQZzgxnuD0YRgeM1MV0k5ucB23YhHbH5kS/Gi4oEXefizwNO5nHFG/qiaIN4Q
hNB5x7R4c24LwRYS4/Rh1JQQ/LjEHWnMeVZFK+BseY5nt6fuVQFwBMbDF4zPRld8
Uox50LC29UASMbZhODQHuoRuH64jb2LUtBTGQkX8/qVKhF33iSVHchoM+dnnsJJK
IXBRUEw2JsQA34kv4buaiHdGftFWHNssAxVSAOpcTnik+Jv/FG1UGngD0F6BRUjf
t3ymxNjlerSpjWWHHaeS0NS9os+EYxz7ACOCgkpqebsZxsKikn4fdzBbdBLn2nPy
ydhf+5TqqVKRaZpnXTCtmLZWkvCdP7Lsx08RzdQC5TdH7DqYQE5LvW+asbIhAQls
Z54cakQJTsmj+k+Ti4+PYYowL0b70GAPf0KE6xkJ7zJ5ardmd/GNIMvkAhZX/Mk/
uitAA6MgYgXpoXWv+sblplOfF0HzMLLg/VTqB1fanIWCC3AhcCM256QNOyy8wRz8
i7+wZusJufAhPs533AGqFfg3rEOR3dHUoNxwROf5sq/MtZiLdsu6yw3DD9hehwCg
Vvq6p/e1zDp4WPRK84Riq0ItZudp8AnVRSC/gWdNLBphGKvifKtwjcbjmNr40skn
d3OOCcE8EfUfRPHjg+PQlRMQuNqSvQHGUWXJJCJzJa50l9Yu3i3P0P7+LyhAc36I
u47AgT8g9ewEbdBenJXj4cdg5zmQnieMBFpdM3kJtoyleE1ALGkGGpOsXud/UBvb
gzX0Rs8zzNTGuU4iP4uPqGYJgO8Vu1FVJ7500Zyo825BYXHmQDo3pdiD1qpq6DuG
Lf6vm3BOpD4UdhK7iM/cOeWokqq+c1kM5YXkdZyCnOBD5ISkicu0BXIc7kx7V9fx
eU9lQHcPSvy21B5O+UfcFQkqk38i0+6m4eBPLlldvj7tWmfzkFYukFbB58ErgugF
t8aSIq2xM7S/OnAPflPpt/f4YAQgEvjKjJOv+oPKEvbzn0/393osRKZ9LpbooWOv
ZYPf05lz0Fh3C7WtlKqeoMUmzT4rxY/LEo/lFeuZdqm8WmJf080U7F4iNF24tZO5
gpKzssF9Tew5H/r3XZVxh9VYdMUL7SqJn6Ybp+9x5q7lHbz4WEHP5YCNAn7GW90B
zg/Vrzg8sM/k3fMpWKHoGz8UmdI2neOCcGxqG7KOw7ol4I4cJ2T0ADTbHvO4+wU0
BL8jW0RE38XW3Y+2NNlI/B9wzR91eJvryWhfjqLGz7HxSum1SRmJupTn4iV6aZ0B
5r/u/CKRvXQuTkYZzh32in5wb/eYCR3jSFYaYGaQUJyWqi1coaxNuDRZkj8N4Q7+
Fk6j/cQK34Y9jvEAWmy+4J8ViSrFOCmLU7n/BApOUTUAvXVoUYPJtkYLCZjCp1oA
rv1oVU9aL7xgTE7d6cMBSdfuko0u9LeTFfZfB2ZpE/4cicNI7gI1Q9Xmn2jJcS8t
vz3RJvqmhaC1gm8EXN+Yk4VRad5Q/rbm5RNcz3dfIu35Ina8qISAJb8E1Hyd5OKf
zJIeLEQ25bZfcdNJBfkr1Nc2OKRBGEqX+6U/9VTG94ZbQOtBzSUNTF50f7AUm98b
Nr2Hyr3N+I04bD3hHvaPaW/7OwR6O6zb4FuhxsGtIB5brYRLMCR9jKTxm3J4AIc5
m6PrutMlSucAJvE0gO6VQ4TP969JC9/fzTaRw2Z6t1BRTvnFTA9bkHzejspxhuge
GU8POm0wlP6RdyT5kVdqL2IE43PtnSMrrB1hgrtZReBc0ruqvILG2SOwKgLggstp
3Dl63RRrpFqB0/HtoOuUXRH+ci1pPKP+eCxSzkEg2Ti0s8rKFuBBQR/pCxrHBHmK
5ce90BQYqsLcy5m9zkKKp2bX6Kbt+JecJQIr0cDoAHQFJaizn/j0kC/tj1zPZQHj
XlFZJA5kvEcX88dP6cQWKqmZsCzpC+rPwbGt3aEJYtpq//8UrTTdGcHmQ1g+eDVE
j+MfEgkQPbXhUhwM9IhmBOCVhtNI5QMWbJvDWJBAAEP8Eq1UT+p92vxjXNpKHWH2
IxnnyuyMQIMgvWKbUQPfXVfAxNCjCHvAxbRoRFxPyC3FnazOkzsizyWcT0FBnrmb
WnHkteNLtuYDtLhaWGVEk1JaVxYf3osO9zU7pnDMSfJQX93Z6E3qLIVR164V56Xe
7CKBBxapiinNDdbVQVpG9dkmbjK2wwhlMT7qbKNGip1SN/1rb7znMkX7kFh90VaI
PDtXlMuvx7qXRXgbouffyJEdlhpOpO3ojFX33yozWgmNyaM+BffAFt6m6YU8KHwg
jbg4jFaZOYS6oP/lnDEpCbsJyYMlRUtdksn3/IASHm20yAXqJpLGLPRZ2XDe2bDv
n8i6zZQSMcO5WWxlA3zeFiH58EYs3a8SuYaki5WpS05zKPwUYYU5YocAi13pPPSX
fMk5D8SJBcDH+OnPaAoYsWnh+Ojgwa48n1p9XnJkNfmY20iFejOAmZzIAQ6eRxTQ
6m40/zwVvvBgV4xMxYfxZmqwTK1ZvoUCXjrz1veWGJ2JzzKo73hipj+nL7n+hNaa
8Rf5ult7/ksz+5IRu98T5UL2Ma888b1NH052U4WBjgiPeROHqgsbXAn/S+PBuO6a
Lz8GdIQ2tU/YXEXENUUOxWkeRyWLr4+IMUS+0ekrhq8bno3yPzRYo0UPieLkVB4Y
KFjaNzsqe8YoewNJEbwMnSh/4F8ay4z/7bN7nh3bg06pTNRRULsO4Jgc/XP937Ga
ynaNSTC2wD/BSFnV8CjAga8XXKgvX8rykLlaecQ/BMKoEtmla2sImtG72sq2VpoJ
1CfYf0XmXWFbGGr5udHV1O83do9pDRe9UWBqdtqy3nwD00v/8TdHoyy33eGpfvGT
ZsG3qfqkmbFL5qiVgAYRl/vXKsTDiCMg6m7iZ9jK4yXkSitP5X2mAPd9QPPrQ4pQ
q8ODsvGI9xS4bzVVp5Dc2fsemQSh32/gsi+BYsvK3N5HFIHKixqmPMHtGmuIcV0z
LNxSYJztvauIPJybW5JF10W1ersE+DvBiSKfUZhHssjQxu0y+zp7H9KOsoUlVksd
FHNbWuAP3goFJqRNdL+7hbFB6TKFlKGH39sKX2LPlB6rWnh0iHkkN0ucojs/MxT3
euE7xqAFgnZPDsu+vPuauIiexFrbreL/pSyP+oB7Dd/JRR7VHWX6d3JoI5Rifstc
f8+S/ZWq2mxUJErasP5C6WAxW+XvvnR4a94GNceZQjotFdBUoRk7aFU7MzNECSWz
NGkHRjRRt7/t5JJ27DdCi8tF1xF/YNRUhWyyBAxjUSOzRItyr904oi13M3zOAPHd
pfROW1H42RaAtQ+uwycOVq85iRIXO/PKhmuSSChtpsBsIi/pra/Smv4zCQtgBYGh
y76TXI6MCQbjjUpauU/qLOzvlsWzK8Xx8AKx94hs5vh5hq1UHZQthdFIV+gPM0qe
y8Kj2s6xXrAOfO6JhrcCbV24EsUBUi8FtiogmZ0RzYWuMYuiXohOs/SdzkzQf6/T
7KzQGRiXP2sSUikWJru6MLTYHK9yToTxtNpHEofmLBNVhzCuh8PFHNS8xgOp0JPu
XcisXFXK6l6HDmEgoi2T/Gh4zHDtZ/Wh1yWJVefTRrPFVbWRhL3AbsHU8LqWkgFs
u1da9byNvC0PRrMFrmzlqYw+WRBmiroaBgMu+iFneb0bjWFHyMvttuEMwm32UNhs
VFtukU6UXx0L1gsrvgo7THFM6SWrubv4NQnsz++/SLB8S1LW1aTscE03rVS1VzuT
C/glUFdvhOXS60Va7KkRSCohZpZvTSp6o084xu4C+F7VqBmM2y7+nDsXr0WuH8ni
A+4EMbpRW0xh4aN29wGarn5fa5TqxX2zAf+jFp55tiJLSIr+jtf2atPWwQ2WAT4v
km/rppXb2cR7hfm/Aj2Q2tlrwYxs0c8PRoSGEFkZdT8K49vskn9SYD5n4aosGaEV
wlmyPt9w6R4jjPPA5dp2hiLlMDA+/btXUlECF5sfXygKcyjN+UxAxWk1ziFgtql9
bjzmsz9aC3iB+s/RJikHygvvujZq6rQoU5ACbOgwvuCOG4RS6tclSGqwIJZ2Y8tb
PTHbiTGnNUHHRguBJJgp99CriAXAYtKnaBMC2aFAz8zHndswW4FFWfhl1FM5jT26
1e+oNTWB/XNV5u+ABMxNBsMbwIHe0HBy+IgpnqofL8vyQU8keVPBoOOqsCg+Xo5B
ekNe/GY+TZ+00JumrEYT9U7SQenj9tSbk36bLXD7jEVuU8QuVgiUBUdSWHAO90Et
EUxU8IL/7+wHJP27BN2S8GY1YWRWiljrwY9u5CEslQDhcAqzy3fvJEVcgwwg64MH
p5fIZ7lAwF8seC8uAa9DRCuAKFpa8TEOJNACjp7PrxVAR3vNe1Qpj0OWFi64LxU9
hbSuXJ2PLo2TCqPaTGAXDzXPr8swJB1/NwE1o2gZlgKLAICU+f1WveBVTiNJu8yd
O4ys9q56QnzbeHHTgEoFCigIrHKdqVB6DXsh/4W1vLTvReVEGOc48hYKySE4/ptC
a8qL8grUwNCLUDBFw7tv35z37qgS3ilImUt8IHyo5ngqOa3MI2jCKYgWBa2rWeRO
VKHhTXrXleieKcUl4PxZIu0pjSmcS2kqbpj6GElB68DasoiRCeLWlFZOSJpIfGHl
pQRU1PuIW2QW57zFyIqIg/0NuhsisvYViM5qH3SJMNB4OuydjPbYg7KjJQ1NS97e
StKlS5xHh36uXnCKGrOniS8/Ziqis52BM/OV1hM7UDfODq1txnwrm3sP9kgqZnKV
39w+R2lN9JDLTlVwCGY2ZDpF+ybgPh4YwaVKMHh5IUiAKo+MRVQzTM2Xqkc9HA81
3yT0xLgA5sTGAtujpwOIB3gIdWcVG+00QElXRupD0m/3tjYoyozQvuBeQ69d928o
+sL9hXSXh75o+MVki2nKaVqVkdpUgCn8Sr6nK9njeMWQhYXiHFRFC/Bmo4d19xbm
yjpMM0z1sfREQTBHIZDKHCcsC4W7u2qRehaRS2ahgpGBa7LQ2Lq2dP2I63/rmp60
EjSDebGY1ub6pn46lghhnEfATmSJ6B8YZsumk7DCHLSQLMIxLPqCdgrqNw2YTNjL
284Bo1MRtCZR68XodQ5yRoPtkgS8/O7lZRqqz+xyV9a77iGIrmwCJmuiyb/hPJU5
x8abwQ9T/OyEMUvCRAFDBCI5nt82QF/He/P3XY+wjDVB1/mqIglcUm3kx5MdPrjS
VaZRt3A+7pkzrMAoS/8FA2mCTPjNyeurupAM4KWgPy9fTqzshsI/Ulh/BE8XbKpj
kcUWbWW66gSlf+K0boKG7wKo0ErZbR4Tp20mFFzGJgLeFkMwaaSOA8ThJw0Q7aqa
Lw4G6VUVZMBpXjvTltfQMmjIeP2prbSUxfq4oEWX7jrb/0S6ofqwv+WhXKzK4kep
e0D6zMPQZOaJPK0H7sQtZppI4VmCHnPwneeQitr0/MItHeuV6nHO6ezQIGY2+UoE
IJwK6h3EV6Ttx7H0+Jx/RKv3nWXeYHsrxi01RkDED+X+8XE1Ivsv9p00fDCQnOS8
Vvhuo/7IrRdhQK1/xlMk9vOKuFyUPuPL09pO/SHhmxMztIdOP3RsE+5CaH+BzS1s
fj5VoD0h8qNylmP7fqYOzzyr5xtEUePOiYY2ie5hB2dgas8GwOyMoIXZzD9hxX9m
OGxQLTPy1vSXrBG03AwD0XkkRjvzDnwXUp4Fnb9cGfsFC3WtFNtX14LaGEnsX86m
inCBaELUWgNkJaF/wQa7D9wQ4LXnVReZb/QUvRoZzaDgcpePvFkzXtnPGpitXPo7
LwVj7FJaPQn6MOBtMkJjSj8rRmZdVHOnS3ZX+tVN7hk8zCdr3sarGKWIGrcD0GSq
Y/eO5I8QXKpIsxWBhHqCRuXTWH7x7jj8kxjDrQn/qfsyYoxs4BolQQL/PaR7dvfo
XwVGP0cElyGna2phRtYnHQ30iKeWUI45ynvuvZKHE2lpJjDV7zVr0siRYY3ewWBf
8gnRz5cmEPiRrBliRky6uj70dXuGS+ibDYDJmS7dEvKpY0eD4vufg6pOq7xcXtSw
U7arVSZ5MzAsrg38xcZAI9Yzd4bfQw1rVxpc+xAEPiY/RFTUjR4yCYMs/o/Szyi2
Jshwbyob+02UHL+4BHr38pu44FqpJOO/V4IItYN/JGuMbsO1TxkEa7OjnLySSIpq
2QQD9RWs/4tsY4HnLAk+flEwzif6Hd/sqRbdLWrC//55coQz8XN9VCOwB2vvzHeA
l+ysb9pFBtyLG+747B32DMK7j2R8zLg2tUezrHalzYwUnAvxeI1O+quWxxtR2s1C
QYwbHwyU1H4KF8EnMHlBdb6pw9NU/wF/VIDIcsxBONzHPDxjelVCtWpy7XyoNMbw
XkiHLfcuHiwMgW07rDVS1yeNmHJL3UgE7bO97UheUhjQqvGW9r9UX2SRbhxDkTba
ZOZOB1+AdiphnPH4Cxtv/8XCNxpvNSOUEOr24daHFEZf4ynno1PlXnizgKPbB4eW
GpaVao5j6AWMfVcL9rnE635XrONSxp7PZJYTKh+iJd74oX5F2mZR+1z8SoioaXHK
5rghNJg9yR5IvUTdwMOS3rj8HnFhDyE0f9+xgk33aqE5uBronXboiZt7LCkqTqzx
fYrszQAIeQYgPA1D7u+2/eNQXKUdjf7Ifv6DMw51tsnzJutRHSB+3l7u1G++nIgq
40JmYpdp18iaWUDm6ZeBO+nz6xc6t4OfH7Ma6L/tZW5pqXuXEtDbdi58jBnF+Twy
7yVW8XUQTxyVHEgXEd9m+MoV3gABLLODC+l6aida+ejqkMluZE8pa5bBev6Wpwy8
vcPGX3Ix+7+i4IRK/qlaa1J+pMb0r+nWskkkGTMqJX7jGlny/Z2uB9LBHbpUqZV0
KWvN961bRUl5xhhqabEaWb6ShdqHnUV2RyBeAEKzVe0STkUAFKT4RDWjeDF63iuI
10pQhk+t3pz/tQ4DFO2kzmg/WurXNsnSP+d2eo2OpgKKvF9MYZpBgI8X2uo9P2B4
xo1vnY5t4zfZh5yAX/33UbPLlbR2DStlOnhGJN/1OrRdqW9ytld9AIYYXm/32tGH
vKWwlE9AC7xQz+MDHcRHZZojQJYGhsDQy4otKGyrWMV4txRkxT0uPkV3fnR4vZO/
g3ux1UTXOFC05UXpR1CpMh7qWHgHgn6PbHCL9AEQC+Xs0KCL/p4dbaA9U/xm+9+x
xLBBL+YNg3OoaO4kLuTebuAmShaMhDo4nDiOQpR/Rj3U0WAmtKzSQWpY9sUz4u6o
+hMdCnqDBOR1IlznuPPaa4xp18WvY6FkDHWX9NlN1JAiUxEg6dIbI95C7MOV0Mm5
S7zskY+/dW9aGmGXQLkSFDAxbARWW8rCJmbsaAlRwUJeaAMdQGpp6qV7Z2+19OQI
DAZ6e1OU5tF8UjvKzzXvy0Rg3EzxLe8tpR1W+ddZ0G7Fw/nuvWFqwWSho4d4ZFoC
0caHyMAonyBicd8OuyT3NDarc7M1OAQP6a+DEGZjY87MwPK5RjyhwbgLDX+I5pEy
1FJg0Z+Bdrvr/xDiq4OXIPS9rmyfluV6IAkCGt+TWOKHjvI6Tw/l83jfwlzV8xjR
KTKjRRAPY5uD5DJXIcKrfkRLP+EMt0obLNHaocdKoNZch0rCSN5y7kcKmwJDFyvr
EmcJMWXQW/5dUOhpLE51pwkPFNLEhDXA9cOLbxXgB4abTnCE4iSUzgSwgjv5LyGT
IndTu6KyNSVC8lN67KtdrK2MS13vzBpbwEVqQtYYknKi1prEwUMVm7qh6EijQvNv
j4xDFGKu0LgotARnAptOJ5f9H76zAwqC3vMjdosL8DYsInfOjCZ08pvlGgDLM+KV
hj+5l4i6FimQC3Oa0Mt7v5He8vNmZsF5+EwLBdk6L7x/845xheE/uqLwzfsUEU5v
uvXx5wz/ZiGfJzpJSIlZtZxQrVV4C8ow3uUBlz+y5q47JjDtYISiTz82VwoFk/SF
B1tCmmu6+2UWFgXjp1JFsk74nJTOFvWNDov/LfpF1bmOaUItCF89toWm5TDRaJ5i
X70U8eKBcSd2n7yps4N9eZN5S+wpIJDeVEIkeqS1nSTq277e2EFicPMmiF0cF4+u
UqvsDwHTdpT/EauLqhSBeqPRSzX8OeXrdrgkTgjOdM5ak/c6u02yAFt/8p0tnmcS
VdjVAjZX9zxqbjnCt8TCzKWs15+6Zj/thBz4Oohxw5I/jcNGcdbcTABHYBI18Am7
8gDe1MfOezstuqd+PZyvYSQRu9pzKcYQ3icmt2GoK4Q2S5d9kKIsYR0/mN7z6aIE
4rX3+sS+3c98v/Dxb8LqT6eXh61PNpBRayBO0Gg9I/K+6LVZPrDgi73m6ev9VZVg
UX26ll1d6BNReMngWVTidPUhh12Apr0GU/7GoJY4V3KGDv04d/xLghsXcXkPPGCt
o0g+qiX7OaQE0QoyEzvxY/ONJw57gQWvOS5RF1gQLpwUqDkB0R/5XNfGrT9zpSeE
Fft5gbDss07r+22S3CA260xnncmYM0aEct8nSSW16LxsMHrykiHn+kMP+gifWgPY
v/ZphpL8sFSnbglONLreavbeEp0koohgnjIm527IJx7qgMdL8tFFzUfH7JUlLI5C
Pcrjz8NkjLmbbyeWCTIlzIU4pcy2Sd7nQcCdw1h9l5h3aS+29DbD762CItbmaoRm
9lJxbvD/4OKHWCr+PosxsJ24F4vEkKO1giG1Rd+F52WE6j/s3riLrjPv3jUK1leG
K+A8kV5xEH8i2WdCpmK2Biisdownmi1mvlLz3+66PLMGieBSQgw0Dwg3fs5iWQSX
qT6TALhtPO8s8+hBDCFKKngV84T1mpQQoUtbI7dyeocu3L7lpkUGa3N3lrEg+xPH
KEKDNKuaOFy89C7yjnaf82j15cenUn9Yy0s0jQttm1olQBWvOiIvqUYYz/qBRWfJ
T3ztCXLd92xecI2+nz1BMZJP2/kSG5f03aCeNIIJLyosruRZHJLsD3ZLRswxfUhJ
fmKz9lEfjE9HHXtNcNmh6dJx43/D+xOMnqtc/xW+7+gABu9wjvJrk8ZPDH3qvjBJ
3mi29j/zw+oGzF3trxAU2tzcVrg6kC81bt/WLgpoT/9CP2zmD1WAjZx3nMGE2tQj
GchqcwenC1wriSHe2zNPb6ZkpI9kWGa3i3CHcyzVrRicwSGmL0pyTyVdbegMXjvG
5Dx/Jtp7u4sGL46+mTPofTjq/MzA0t/M4Y3btJOjhutZ4ICVFKDQ3lTJ50RgnlSe
sLjVtwSlc93IRuDjjfGph9eh7JwJEcT5RWOxO9c6i6rIvbzi34RV9o7jvUQbe9zn
M94oVaarof2lheNGWCh9Oh1bKGB+E9Ab48OmRuEh/0N7O3zrHFly0PPvW/QaeHhN
QHKAYKCUoW9ppbRDdOq2V0KtPYnlFC+Lrxjr+H0ro/3AXKc9U96wa6wGsJwTwreQ
jA8p6iBG9WZBerpX1h+hROATDlsM9KAS8DZsZCfCaptQd7qF6sIFTdHbWLDZ75fw
2mc4hIMKy+rZMUSf4VVH+JhyMwQuafr4UgGmsNJ50rU1VnIlOr0+ZocT5CwR8+vW
FwYRyugmJTjdN2K30fCuVC+mwODIFRztZSHhv0drMbfRF6BjhIMXtmgeIiJ8scI9
jOkkA2HApSWOdv+m97AnCKlTg3sYVmX14UUiQKhYIZRpwondhx0p6Q2bncADF9W9
1eprxEp6bb+GUZM087KAxUSckqTSnfovUGvBMPLVvgkT8FTtKOJ392KvaaaicPfs
fZcDurvX0GVMSDVR3LCZ5ellNv9ZaHHPQD4q55PZNb5N5DEzlxqO/lBR2zqCvItC
KTub9mVHnwtp5x+Xh1ofiABoyH30QPhwV4uOPbuMVofCxVL/QJqmStLZeDcX052V
4Q8cDgtfrn+KX8XXzzBHH4//fiQ4c+JbBUO+Hf6WE7exeuIFcaCUgoGjqCItQBLb
N0zQJwiaz8QNKujyiKPVNekP7kZ1n4Yv5jmUL9OBl2QrBOGJHfZ2EJG4JZvkNMBU
4UtzEtBzfT01yldBKBHBctvezRbt94GHolojJW37gC5ILZclubDFJVbKZUbn9vd3
nE1p4IDZ2dAakC8niLa4dQJExz7GuSs2c0TrS5oQ9RFCLTqUzpvKI2vbfnopdAJQ
pSaVh6SJSrllY47FUAWGzGLpZ0qDcAYKJ+0cgeIRP71923Km2Ny67u44aENAKj9D
yG27oUgD9SXfnSwVpVp45n1+5d4wxZX8f5b/KBMdYJA6BdTZ4KvE0upv2WWW3XFx
nklzeFw7qzuUmmkqmS8JakUI4P9qjpsJTLRrsiPOOpd90h4Xz+VAMZBWXGqWML1U
YN5A0+ZExc0wBIjEbVTFOmgaAt533ttnraJoALant1RePjiPzDl4OIiV8y1fZe1G
ZKOgm/m9AkHdYEi5wGRLdrqK7hUHcK2a6KcMtpzKxI/IJ4smXs3Vxd7rfTq0Famb
HZ8UhaItNA32UI9bnKMQvDc4T5oqryi8tC6Q14nwdFR5VA223y9bFXk23NQrqxJr
vLgwpnj1M80L4ioIs1cNvfdM8OdWL7PJaLibfAlMofSQndUi2mg7A33itWDDLM9R
4pBffzrRtUsXa1M1DGcIrRaCl1uBt8H1rFbplrbczsMb/CIjrclAlrHUCc93pc9q
00QTJ/2Mi3biIUbIuWq4RIcwTbH45Tw9Inpxy9w8JT3o114+DPkZigIGmp9H9Iv7
ZneZLhsNTKNplTqfcg1/eUUBq/ZBLOauDLcxWG34k+XsRl/GFq2zxf1XC367ytRK
IWdkCYSxOrDzik9sKQx3EfKYNmwK0lo1YRlJBcntKH9NAtVjSUkP1Qg0DebBtdbr
3675Wf/s4/0Mz4Y1JUrkMYaPTvUHuhIgmle5oV8/I1kUw3fAUFmFGIdSIFz2FZAk
J8v64CG/P0h9ALGG+k8p241GU2cRPq4h9avGscHHcyv9SLCW3eGePDZm+/6MQ92H
Aes7SdB7aQVw4pnviNl5PtA1/nM8+HBodXNjOw7/lZJjqOyn4JrBBhL7sNkUIe4j
ZaEBSd6gv+elczBcKZRte3CNXfxE860Y8fjM6hIaywd3BdkdtfkTLZ+Di2zrEfIr
oqBxi7q41YFwbE/6/hCi/vD8hUhzx4DDyXTLng1Pgygp4yHtHUZrLzbQP4lhR/BX
uBCLcNY01FcxBTacoRIylVA0INxaSVP4CHpJebVJhH+dTmFoSPQyryPMJ+acJPP4
Fq12CDmAf91oGwrIAYIdZAipS2g9Vq4B3/qvIPDKw4g/dTSxJpchCZQn4KU+TbKj
oW9B2sEwxrD4RrC9lrlzTmXa1wk3fPDGl4Y1pLywpZQKxm1CpC3OXfvjQ+VMDqaY
bvTKyFTezOR/L+ycIYyeXguAVAQftK6oE8SWE9KnTWpXOmQTEjukTruQ2M/QL6mO
YYtHlInceApT8H7V3iecSJEP0RKSBSi/QpZ11JPq0oFWOk4AIARbVYdMUM1r5CQj
7pLPsGrpHfJEnWVG9U5nAOAcGWet6FsvjcfPoqqW19aSYZLknKhdi8RG7LIop6ww
HOKPODVmZqbPQE4VuzNYtbU/DUYfngmi1FKRE4o7CGieQWiGWb0XZs2xNu37H89E
KeQrYccyiOp1+7um803mjOYV7Nckz9ZUwhGTO0RFS8ZX3BPYfh5EaQsGvUOMLoJg
iiJPJ+x0yMAI1n0moMvJAW6bFsywfH/szOADHY7ES4MPVUF7nZSvW5k1zbWoaaif
nVAvtx9Aam7Cy6piCs0wsH67vLOC7sZDcHbYdIx27PINswCJHbTU3eU4FzzX3Mdr
9hxwoUu7gfngVqfrw4Efuifh1JDr7r9c+j+hFVwoaRV6oz8AX/MRmPkjG+U4VEWe
Vk5GiGpEpDz8SRJ8Dal9lKmEqnHICZDUXMnDUO7FwopQijj7I4utsc7fB6N8ofzO
JsCw13ovIE7d+IqV9CjesXEE4vV3+SlfGDAWT4wRYUumYer8mcIclNmlgnAKKNvA
elWm3UXLfda+639IgWwNu9hIrqPXuqZVi4uERRh62cgvRF81pHPp0wSL/CkEGj/o
MXONWNcFqjAHpYfF1CwOO2f0CmGFHsW/+yHuwzIluXI2d3EJk+sfpHVb5o3MOMvr
Amd1s21awf+f6sNAWNuli6U9hwOaQGl66s2GVDTWSnJfNmYAlF0+7FrnII426qCc
MeHwssRBYEBZwiUzxJKdJDBdiQj5A8UfsUaaFV0jDTJYyfgIQ+SugRY3/NSLe6jm
IEjQBKH8KMiZjOB3I8rW7NJ8MdPDsrt6sKruicpv850GSJcOrwfliUoHVwtnvfGf
yQSfrs+Vkoy3tvfEeErGk8QSnH2Bp4YHo69S3mWOSgK9r/ylXxLwoLQOESCrg/RG
pfC08Amux6GD121PkW5PCwWTqhAuqEvEkauCLXjg+2o23pbV2kIDy7lBuRVijD7s
1WgvNowHD2wxYpQyXvW1uOgeRqSow+lhKuXpEI/JAXsuoPMwQmB1pfNL6vHRWjD0
IwU7gWngKKBKOfHweEiNDJhfhHgnIYa5HrCgvKs8FLo3lvQ8sZupRNW1z+NRbYBH
/3aCDSrZfPYPjOJg2b1+BLOve6XgJBjMATluqWMAYOyuXTbqXQvSrCT4HmTUgBHR
80ofs+97Fl4F1xWZDP6vaj3X92CxDqf28/dFkKXodZ7kd4Z4UudvUZDJ4fsUmieK
g1gGl82riihRWNdIp9dMJThy9RhABtHJPi8QfuxvGUXK3A3DyPzQCvIOwRLmN6/Q
u6fHiHWcGs3UGZsFNdd+x0cdeggeDSY4SKhBsqVXhMWOC1njbmDimM+tPfZhAxnU
471FwfTXZ0D6MbDUtqlC9fLBiVpk4PMQTob8RFRL2pgMJuqAv2WXfkUX4Gfx23Ao
v/4UXf/ok71ObkEqwlBX8R6oS9p/H5N+fK67ekC4Ns28gNTAI75nB2y8gaYuo0L0
+qCUw/DuE11COFIuI11rY/wDLjS1GEWjn4fgvCqarGqQGb1WK+PWrZHvgPudTrV4
/dZPRQ2hZ0VfIoOK/uf2SvD0fME7idCaD/AsYqAqGHjOrbBzxrTccjG7OQ+e1LEV
g+xbC+EsJUA8AG3bE62jDDpB8D+wreSg1HaP1b8nuWlNfE/ZugGYoNOj9/Dn+hwo
jxZTOd992U13jfFTbSCuDt5F3V6i9H3CSnE34b59A1Ymkw9Gjm76HCN7Ch+AMnJe
y9oFFCbHvtgd6aAL+imqih7Ki4KvHaTB9+SVQPF3o7Jkz3CMnavKgwn6wR93BC3V
jPVQrz4aVQKkqtkyl9e+Zcc4u6gklhgqH7ItR6e32tANVLr2xxhd1OksGVmoZsR/
RGJKCcXr/HJ4mpVALX4phrho24XGY+zTHelTthawhJFcPyC5/+39OEeEjoK7uu+R
mxYMGZrbsiY28Y240u30ZsX18f0FwcMyX8NC/gmd45dYpvg846Vj68OMJf4ryacK
StDhGn4oBL2Koc7w+Kw+QoGG3ZJw6lQj5OjNx2gaLyxMs5UCbGUpnFM+OphKBOr5
V5Unb34QZRTGhSXrIg85Gh8S+WHFxDmUcV5bXHri8QFAil8pODqT3WopNqAm9CRK
iqBM9pyQk7GwszPwGkEEEPGwScFEicEn/vzDoRd4GRKUgSJxgS023u1mV6WVpNfV
3dFfPaPDMqLxj2Vht6qM6R2VyjhOhKgrFhr/VR3T3X1FYo4w/XQjxqtgntvWzCpl
jjUY7Fn+3EzBcN/Eez1StIczu6lcY5wXv20OZFGETmtFWszD8CTVshvtcbVQZGC8
qOOX32aSFfDVCaDM9wq4RqSE0qlYEwRK/8wo9BiHLN+7YhGHaQ/h14HdRey9C9WO
pZ5x4pKuH7nfV1gSghn6E756u0V6yVpK7fj4aMdrkV8IVxJnMAK8Ff/WYWGi7Pb/
ekA9KN9/yYAsqfWXT0pGl5WtRYV7Omkc5MrfE8U3HsfJli9Wdz6px4Sd2ZhPS1J0
IwhLasbPqtvLjWHrntXb03FVePk8cuHLISkv44CySQKDHxbkKEpnLK7Ik9ERAMNf
PgDBWW/UFy4vvn/czFaa6Tf7IO4SXb4n5qJhQ2MJOCE1t/8T3v55S6ALnEWgP/q4
JtlS5ZYSnLhMvBmf3vbJlqtdFt+VRKQRwOOFdfuj9xm3p9ASQAun/xAgLi1/8/g1
FI/NbUo1iCQhMlFI+TfRxTpDsCvX0nP1ZdlonH2ESV+JHbVnG2OpzDQWEQxmM8mh
0Co7Cfbhd6vj8jeDg/OsuaDWh+2/MXhu/3MwBw+mUDy4twoHesx3biIsjJZB51c6
yzME4eUr5ubDRwUrEN1I5vA4jOllYlSRIfmD7U9DV2D8jwZajDMtI928w3jENTnC
usg4Rhc/Gx7JnX2BcLoiGVsJ11Zxv9ACHtJXm6/HWeYtDlUngZh8iVgoDlX0yNUR
QKDmQKGhkROfTtfJJ4e/kpP62orlcRLOsdZb6L830VWvcRBjXzAG48eYdnXuv50f
YWKAHTM+wm47cz1Kl8KNmxVDd7P1OXoixDOxk90R0CY3USNjZU4JXoGPZmy9OvV2
ZWtB1P7PuZI+W9X+Z+VY5+bz9XlMiI1Qnb6f/hFu28Oc8QOAiagLuJCzpnvv1JZB
V0SG1Q1gRtoa7UfZQNqjk5xfEgTLxzerD2lBOCaRmrpzjNIVoxFzXIITPz5pEGkr
KlT0X4MlTejm4Byft4fzj9JfXmD7WUjBhSuIkFRPHjlnIR7Hidy+C5kivOkVn1TV
07XowR9cupA5RdMn8D/Uow/v7/OyAZHHSZSJkSOeS1D97n+7362MN5sofhD1Xn4o
BSz/j3SGyqV1gz3QxIgGyBi+sREwBgw6wailCVL/7UJTBU/mH8aCOxHOpcBgaLsx
GUDoad6HLHejAL61m0/Nx1CcZ7xN8S6hTLEmHt8mO4gPYDDZUXmwzXHSsSLQPhrM
gz2XC04KsQljj7MwYotx3xh7gXqSSS8/C2xkht/zShN4x9SYX0mOCYB4KR68n+Hq
naeUP1+SorIGKxrYKXdzH5oNMV9cZ8v63goLTew9nJT17JqX9h6RLnm9pOuOPxy7
XOzd2/lg/UQYWNT/zDlsNXodTa3HYvroMfJdFhFvrVJH/dG0kMNxEzBa1OycdnOp
JdskigS7Ht3+q6VHzMTkUQV65fbhKP4BnrUg3DJgKsbotyZqSjiPKchSQW2gmI6U
s3Rd2stL3XzdTmfNTH+Dc+T9hlxIbt7EMkdXSo6T6QwO6B22iwMetKQGbacO9xa1
Cl37fQm1Uf0t4vqkwce1eHjnCDFm6Zkb/JrKcqXHkGGeqvj+/jHEoVzUyoYnvVBM
qTe7Zl2RKyhdZhfhluvsusxw+xp2sMdmBHrkaTaMzvGXsryaYdjoeFT9zZTYaOWK
x07V9oYMeLi1P9A/yviQ5JZNr8aNw6C6VTlCXt3OEMAGFiAq0omUCtL4RPaJQsSL
sF4JUJ45MZ8lo7KK3/1SCFqAK1D2tELw3aqKZkl7Ukk3o9bFRGByLltJ9R07Jf1Y
SyoJBkxrIKUvNgkfMHQhayxh720I3LdJsJbki9qzYf+q7rGbVI1Qa5NM9+pUXDmf
NP7Jzp1uWKcur0oWqCuB3dpIYZ3dJBzMfR48RBRa+udLYUGvOrQH8onaUv6DLryv
SOZRLFvWpiJi/LL9ZJXy9GNNn6myb8smowJkTCq4mkTs+CO6SiYAh742TEYQTuiD
EdUdNLlesEGNBUnih+xb9EdLZIpit1ugQlLKixcNg8rTqg47SFrdHG958sR3tWNm
eH+gEOarmuvNT+ZrfvBFabKyKznUvfbWU4LMLEzIU6JCWukFoTalBlncjmlsHdcX
G/Lc3dCHGuPXYgp3z2pd4MWu+I9KQ1vXK76ssicbX4yvMDem2Gser9FfDXeaeMAg
D3yIpzNYsWHZPqUQro7Es7e2IXwX+cQxP10RkzILedYyRky8DuxNOZaw1alugrlj
wsgpdAm+gQRlPHMggMh0RDR9NiI7GwO0lQ4JsTzurIqfO94UqkrpgpxE5HadmYZY
ccp0XBRQgpEWVSX1mZpkbpGZwuKcLX+u2fi56OVtyPBb9McAJ3Th/wPQ/kPwIJPY
dlliehhVYpjk6wVYvmMbE08fiuYI0/u5uhpCuCO0dw1w38QBI5yPmIWnt44LfwsI
wQ9TxMGESGtuIMtXPuyGWM0r3TdSLFhfDnV7DJIVF5/TGmORgxRJRYaySnZ1bgCy
nNMQuxVnAvHA5QCumEzELxq0tcVwPVY5NHntffZG+6wQhECFOPQQ2syiPFnMB06A
nBLWU5dmXxdADLIuRlESVEAcvHsCjDbFY5+vZl0RlOyXtmcKnR6KDYZqZSWbaUO9
2NVtuJM6XNgO5vQ0VxLDfSYNbMxuRbo1guE27aAcG5QggECJ19iTxSd0yOqK7x4l
pcfe7N7nFzicvEv/QIsMwnApf0A0nsYfrI5Ll0NBVjBjQ/9e5fBeQXPJbMzTeMfy
EsdZ8lxsomL5ZMy4OOo+Udq75OdGkSNEhQW5m63AipX0JwA7888vIHjpFhp4QhMf
53Y66eV98kkbyc0P1mtH8tjVe9XhtS4F5I8C5WTqKXWKXEUQFp8+0Td0BKhpoI+O
iUQ9Y+iGe0w9nBKcp0HI9BDyh8hqme6IXalIoTOBLtPsk2FrARh30TKycTLdBJSS
AsPQwLCt7jdpD6BNk0RoIUEJ8PcpT9P1dKYZMDleCuywkJI7OZg/xCNEZTc/a4vB
9rdOJIJta8fzZVTwwvefdTsBW1S1Wv3qnAJMYCsvW7DgY/VsVEhMvfvAqsx7Fyu8
F0YG5mUuRSVpP0e5oaEmF0libSOYiswgQu+GCll4mwWuWq7JXDiaksPs4I+clAwh
ZDdnjnZPIvvbepRsOL1O+1hc9UQKTkEJhwYHl/s495lh/EJvFnNsZncywXyXMN5Z
ZKOhdE4wDQbiPbMu3vGtwBicWdmbU5ML5om8KOxbO0TK4QkOmwvc/7YM6GwvKMjJ
R/cXHi/04mmuzhtHAtoIAIZv9Q2bWlxHDDS6nTo+WQ9fx77FMRQCzXgnXw2smxuw
PWJBMnuk9mJx0GmBWvs9J6X05jjK1uIO4AnDkiif08Po3p5cyZY3WHv98QlCDHza
bhImkW46LSx9OZKcq4FFPVIHwZkgF0a7Xq2+9jitEtebLKncOq5PEQqATTu8yQK0
YoTbS6BppdPav3a6SkASPajqjqNlX2Ge9Za7zZnrg3CVRxZiUkBNfcFx9zWgcFUW
8I5mrPj+t2eCJk8CQIvJPRhHuQ4VnmNEiv/R0+BRF5wQmG6JiPSWcAUvYRywgq9i
JaKz7pcGquWmZYetTr04xAQtXu5k9+huIxHmHFC9UgYf7tQ6QtrkFwIKSSWzEyPV
xGHh0bdcvK6p2SeF8g8Onp7z3roP3attQ7A5PQ/gkYXFYbTl7iZk8zBKCBgRXqZ9
eaSzn+OBILl3ZRjZyGshun5eKllOecvfTNEeq+b/R+QRmt38LTbiDLC1NOpQuwQQ
TnnVJR5kJW/ybwf9/2vYYF+LYd3z1b8TVbd+kVi5o9U/vr/ZJZiTIykl9kS0qmL+
OSDL2t1uszysUE21kp+V7+Pdx21l/Azr/TyG26nSxYhOTm9buAErmrwOJVu3XWqZ
BGrI7Fcfro6dZegAfVE3wg5ZOb9BXvatEkbz1Y5LNDsMlWm9l6Tvpr2kVmmeBXaG
Go+Dj82ZE87NSCuFpsOHbE0uJSmpIRgO/A1pey0MuWIH29NaxVuXWS46FjAlhIrQ
6+0fonqpxGVF4yN+Qt3O+z5t/XT3eW2kWyD/0WrnD8Cw4EpdgnGWl62ebaKNwWy6
/E2tEnm6pRb2SiKoNWvSjABWgGBN2gxzAA2zGQpjhuz74Gj9BrVg2e6hiAOnbWvn
0N+A6iOAm2W1JJBjRJuTzTIewdz5Q0LX5RpMS/bHsrGqW3JB1xwHA1oEGguJL/7t
LmFt678Ljz+TiNXdXzhXY0gVTMkkrn4j0cFguMvdrj06pEZ5ch/8vnHdVWo26IjW
uGBESTSzEPAfrkHiQ8hKrFu78rOlW/lm6jHrldqNMzx7SQPlS/DbH6ZQQNcoCT+t
OQmd3XcdIJA3WSeSOyhLlEdhaM4AXc9vAYyl6GIn1B4pZnaRcduKOWE+4wmlFiBw
Rc5TSSA408JwmxQ/L4a+7sKOrjyNvfbEXXHVFWtKS8dDerh4xBo+mDTJ49rQ23Uk
6WM3wgVwURLDsThrn88arA5MomVEwIvAutN97egIgoD95kOQpaWHEglJmA/TV/ud
/tCk+jiz6YVwkser+1T2yfusbkYvozPtjp64h9KD2mBY19xysnVqDPzvQE1skx5h
9+64x1xsOzqfac/i0GN+k7UCL1p9tgNAeFEHnlA/ZvNNF07eB5804s2rgAz0PKld
P2pelLUBZHtUP2+4dilzcmn1gS9N7etpHSxgJ1lhDclI0mZ9Z7i3AQRqXsJLemxv
39pbuPzGQY2r+DFUQoYeWUaPbCXOf8pKioVKpMps2/mQ9FqF2z8dwMP7YMx3tlod
H4JA5QVtMH5OylvT6UmehTulyTnnAo1lD91aGN/LwXhvw/KTf5gyJBbRdxziefx8
XvQZdGj/uLUoU7RhiCxg2AX5894SHH9z2t2JTvvCL31YGZaDXiet5Kirb1fMWmj3
J7WzDzf+bUPJctAl8KkULw7Lpy3hkwx3B+H3LQw3gWbqs1gTuVvl/f5jit7NrcIY
8MT1f6EYOPHct1njTiCn8NEOeO3Ql4silwz+pwfw47Ik5sc7Me7VGvvWMeGJqbId
9rySK7jSoMZCI7Alp/TCbtRI0j0d9XOYOoxcLGKWfEcDfrSI4lSvrf2O21t6ahzO
aziCHLWP4/g/GApN8h6aYE+JvjIuD1ma7K7pskdYugIf7Txtz54Mzi5O8tBU7j7w
9Eh9M42gLGKVJBxjYWPMnF3N21igBnDuiEUa0caBWsAuwxb/A2TwedyXytjVPJ6D
jM7s05ysIMnNp5F83WNqAw5qfmfMP2tXkBqjgoN4Gu2ZfN4rKJKzPZHH/4utbZoa
/4/VTDgDBCw57kX4JgR3PKm6lmf/Z4IoR88N7J8B1kvCSOO5hod2kWrOOsBSv1vR
NyscA+0gy8EX07ODxU0LGQMJSnN8qQR6raVvdNvF68jhHwGFDG36+Wz7JcvIzHrW
uGPuB0ZHDTB0kwlTP7yoHnOy3+nkeiG42TfBP9bzmGnjSmiEf4JVEU/W2wKw5N9M
jCp1bnIRbGwSitBVQ83bcaOJrqiqbFefbDxk7zW9aNnojsLT1wWP+BSQqN7/e4Ns
ziECEBF6+HgoT9LIbuwK4l6EskeraVNvMTqSKGDWHTQCnv/fXYWqr2lFBAMY4AIs
vZy78A/xZY5deGbXq95mMOlafAChzT3KQPvuhdEZR18vWLewSLIofqh74QgyBReW
hT3sP2nqUMCI+4T5DNFh19uRGMj/3UuXNBLIBhlPXJywVsAZsMukM1cmV7XngCbw
iCpbKPK6YBK8FN8bR3rPoMT8S5eDIocgxHzAiRB1ix9NOA2ZViXktth3TXzovbMW
2UB7AcED4CxGtlUJcTpYxWJBiJnV0i16aske0r7TBvoc+3Tl7UZsufDSxOrIWFJ6
9DIcYe6zuiG96t4t5s/A+ILAeVe733od4loGcvNkLtjwpfqLGPcXDqf/lzMVGk5e
mR3iDRSABn2zSErg+VvJkCndT61hxu3Nr5vk8791m9AB2qZK+VkpBHT2BprYBIi5
yy5i0vhO0+DLl0HwawGIQOxKGmWfuGf1mfCt50eUFKbNEmdNm0xsQaXskPuz3uRO
Di8jJWXVZ5Wn8CHf8KC8O84LCX+JpwbwuyYJWQNavgQ5afi5ZtzHdlVwIz+Y2GjX
0Mj6u7LFb5uy0AfQuad4CdHyVf+Hg/SNj0wAzgLwNr3V8v7SdwTxtlSQMZkTAQMV
Jt4EKqf27RPQ7uCqqlu3BVx523C37BqZI9J1gDY3lR4pFPHaPfQT0xFoieZIbBbN
u6nZg6mgO/1kntKN4iWg8DimLpibZVjsPFQmJcuMMG44ctXs/7b3Gf2NPi+A6JAL
Xuo1hM+Ct9eirqizUQC4Wr62Z7mIBxWr6NmpYb9j3PaxIJ/zbu1CD/F25LB5o7nN
uyPTnGbNpmKG+Xxhr+6uH2OYdlownoL8ijNbPhAftjpVP5YDVZTN84eHf0Hz887k
jxFxFbMdY2cDPctMDIJaO8U/SdDg8sI1YgIJO8PJEGTxpSI8Bti1bA0VfxazZbr+
gJusHJ6ju1+7gI3PzQ+s83Xi8RJhl7yfKDjPxISTogszVmI7YCMwM19DONhS3MBN
6etdFEP7osvq7uClzfu4dciZghThDZ6+nXxGzeoVMeKkgJQHoX2pb+MAXWcTJNFo
TABshOQLdtgaLhLJkDaYI8oA/bOm2RiB5/bDDqJO75uLf4ZyI7LrtZaneFj/dDrb
/FV5uTylVXfGZ9QS+JU+lKmg1gARuixetRBjjVo1NeS6vANtQGEGINPHIBpBbPrQ
wtWhZPcapSdTgbK26+XSd4m0iMOIca8ibnjv/9NGQGB8mDC8l7NIo1WkzcP0NEHA
A7sTUp847xc5cWxQDp8VJDVJ1Wxue7ja95a1tCyQCCNtm9rItH8lRWrWtx+1v7uR
NgKfN0swp/wVYHBr0yVqQVJV8GQOtkWMdxOCJGctZVEpBOrj6kITWE2eYb/vNco0
VouH2+DJOweZdOZ05jMslnN+vRYDmj1I8u/ZmLsmWJ3mrRxnW+elnU4hcEJTg4cx
L9tS14mz+EhvDhRo9FtRpKOJnhvZ4g0PoGKIrpQyZop+3rTHiJsiGRkHOzLGXNrr
mmsgYhiVCOqiEdAj0xGe3qBPdW2e6QoPPKPI5syDbDM+UxsbiSbhwPjj4sYLAAzU
P4Bc7t2dFbDLsrqXl8QO7/RQQOC3qVGgAis/XgqtM//5QCiR0gHzduurPHbCGast
B+mwTAcyVhC/BuQ08GeS8OCK2FdIiMT3MvKNZBLAIpng66M8qql00bMn8GznpLB5
Hvu+7rZFGuqDi5eKEAynkMrLD+SMeeQ8391YvDW0PUbhIklFFzKXY06Me0PkApuk
Md2DhNI6DSORAe4uiVQXHNXmKXFnL92bvAHw/Rb//UnjlGZHQBp4t/F6JNEioEPL
RH+M09Zzq2/Lq+ydQVnaPffoOCa/EyyXaPxpTMQ04kOD9XJRWySEI5YnPX39+2vb
nv72Qmk/a5Pieb4n6M0XFStPtI8KXyVjp8tdfY0nR/Q5vyE7+8JmnvmhqHv+n2lD
TeVM6ncjTQT8QOKBPJNLg8OZT/70SY0J/I4uz/ytb9NDTdsxt5Mw/SW8B6663cQf
FA4hVnSemXHtG0hWYd0502b7rNs3GNfV2axXz/sxBTDLYbFAsFAcSuCCzEblgV0M
7R7RSycypWB/oDcRaFUBBJX6HZL/gNN5q3ywPBhuq7CKKL9P/1uIhZT40SDWkNF8
2SNNCje/ZeEdluZzM/mRsINjzN0w/fuXkH/3hFsX+YQ/a/yzuLVbFYhFEEem2cn4
XDTOCf/Zx8CmwuSdYo6bPpt2uQL0kEKh66rJk03F8QG9iEs7sAEezOkbnOcJbueb
+b5eceWatbZU2+9t3HJ7bIUuc42UwFAcIIXEJEU39bkk6WNmtpAjnflmotppgP9G
zEpgjnQlQFPMd5TY8DpSGqUttVkfekTcx76+yA2yCyS/kPnAHAjY3mDEKhy/uJDV
49q4rxUNhDxa7LNuf7C3/FdtIxHxlMEV18u7Z9vAWirDevCOe+oepx7/vICzSLgZ
wgcRgOSi/6PzOYlmDr5wUej4rqmecvDql2R2Qu0El3GZi1uDSXH5aVHj1s7ADx4n
5u2bAyeFSk3P/1CdIYfxxEGqGaIA8GpaQZ6g/VNHsmPRzHxdonz5ZVX0tIQsZvZw
IG7lRe+1uWQvbsljlpMmjufXmO2/Cp/rERefLZRURknji7OqGJcyoG31AroWxKuL
o0mSn3YDcIZqls3PiVtex4fmAE1nDeKf3wOBP1Ljh5gkVs6z7s6H864nQTIJ6mLu
SUDrW9Mv15pnapJC7BhvEHxTxmRJVBkDb9/wJuDFteQrfOsDv1P0IZ2yk+iV8nPx
9rwRoztyw9pfSMnC7YG0vEUfL2AliTYP1OKnbZuCZK/X2fXug6J3iXHHHuvGjdRR
GKIQlFkom1G2IUAR44exJ/ZBOFtKbSzdBdUbPXcpl0WiMs1xFvf2O5201t3JB8ZT
mq/FrxgAsD1lNSNFFmybQZtRAfw3VYqOWzbgfuKKVrn9b3AzkC2eRatMXRFf8BoL
XKf1wBWslPMXmm6IRACtf/J1cPnmhcWQkmidPZQpALqTqiZAoAjVpN9zeECzjt4Y
WPIG3zEsZMGnT71vur9Ar+qWpltpSfZ0hb+YpEyuuWb9Z/k/Hg2FsVagt9ttoG+B
WnUFCTkZOJkm3a6W1rHJiog2T6n6RWaX78m++zAkUE4njrqrvSPtGrphgWzJ+4QF
bHh2ekBywI1odYeRPTy7XBMSy8kuDwAMrKeX1liapBN9xFrJzt5/fdCQ0igPQ0C+
IiSUDSS/Zp7ApPgFK0FigOSSiOKxEqWg/xdRZA6dImJo6e5wuojNwgZ8WgG2MJNm
2VMO1FVsOYMLFafQXtSFRW11RF8Td3/9Qf4CAbyGp+Lc7ywu/OXc4Fxe2TEo3CLf
98vcaoodKwpDEwrwd6jvpMe4IbhLLlpnTaW9CXNYNxTyJ7DARBwc57+3gd1FcI/Y
HbPCFq02BlX+4q7VWvSHRGCxcJLaglkNM5YuOsPYsPUzqjowF8BIN1g0rs1/p44z
Gyn3wgDsYBqm2DXhYVVFq+pXDYLX/GqVeF3Q2IJfzhKqB8zGxkp+TaQX8JS/oppW
ny44uxFeThFNQPcKZraxEDC4MGsH+yrp1lki1yAyak+RntNVuNRF22ZH8rPogI9n
bqdwHQwML6le6rS0M5E/otZAIJw0mIsCvKrkiZjRKFpjgZKDbnssZI5nqrZqMQYy
gDqrz6KkyNISnDqx3KtG3xfC0Cc0cXq+6bzZI+2aCilQPHY/vR//dqoL8h0sbXfM
nPWFB8TTwpRe9hgyYwUvy9cp7N8btiI32ClwtjS52SJUQY8UR6qiEAa3uLb7iBoe
KM7ksJBu1oWqoLgl6Dri0fSb6M4DjKy41ZD9kaarmozVDbxFwkvWETTFe0eKXMZO
FcURcO7PwrABzozua9fY4UzWwB1/kAGQOWxFs9Cuvhrb1hE0Uu8uJNnb5rZ9oF1x
mXU1D0vO7ki598eXp08tdOu6jkSKLZXYp5E4+1AjSdnpei4NZ0W/xQtcbE0Sjorl
6le3HJakNtWY3AcwCzTRdXwgQiNBUINakovOrgHetPf9jOabJOcY/bx93FmgLlt4
T/lOkITiS0aY87wL1q2Vb+UsadngeTx57pLnm93fmGDWnMtT82FSOQ+6tsdObYma
qKuiTITmmKKa3dMc4TL9UYDsD1GXyUFNC4snrWFc8K47IiKUKXwaZZ72083GCqCf
9+NllEnlJJRE1ARnI/SmAbGHxH2dU7M/jFvfSU+xbe1tgvINc39E/u/m3rpZ3STC
FZ0Sak7VqHbgxSRC2nmBdQBoxSg7fBUJ1lMvfvYvWChqAU5GFGYS0DqtrYM9Y9sv
KfGdux6zTNSFZ/1uV8J/3yEodklP2r1Yi+ZykY8ew/n/MSesCS4Y2cQlLSKc0NRC
18BNWTZQLspl3H7Kz/yNcwTTrqvlHI9U0UZqDsHps5P0sunxxfTwB/NjUieHr4gx
wTcMBtDzGJIx842qtYQjcZe5A2sVxTnw1sdXBYRKxWpxxoj/h1bBnYFLyxPe1A/c
um8bpZzfRyc0+B+lzH6xqN+FQFZoO6CyIRjBHuWzjtFYixYAcCrWTNgjKAWDE+6O
Toaot/Wl1g0DTXAR5/1++x8BUdJs1TCMJYCWGFx8yHPqmEMuMvs5J/diTPBZfjh7
C3tcLtdlmw8WGVJNCejZHDEh1wBcdIxa8SbCbucV1O5luyhFScvo0oE/srqo+x2l
xg6oiVrp5AxmUhuewo3Ch3y3eJd8zk6DTvM6JB4zqrKhJMy8tGVK39AoDkGFWeOA
6LLeycqrf4pabde+sCN8r6YMGuYR++DB4xFzEdTkzo7kD5qdu/QQo5mSrwTTOvG2
Rdxz8N27KEPH5XML+9lAjmyGqddpzQ1SBfg0Ho6r7kk/DeV/LUSp57d6zJ6iTHdf
rSxSrcomfMpJCkkzlxZ8TOeWZE8zWVTfe6hF6nxYooBzmg0NKRQYzdt8zSzgFG8N
wFLaZYmArBh7wH5BrVrxl1JKx5AfBqV9iCP3ndwUzLk26wqTCHOx3aRcQPD/d8ah
ANkMCsjglHQCzIpUMLTyJ31PsZ+LVP3ZuEPlp6UwjfeJW7asepIZuDJI9F3JFINF
iTMGpHcrMNmIuHsTDDMX8L3tCCWH0doZa6MuCgcMLCHY0vYTLAD58kmDpgAkwXF7
gVmdG59nJFET5ZpWtqQfJNoOSaXT4oA9VrOF2hTi4OoKQtAg7X+n6iWF0GKR4vgp
7TpxunwdG45oZNPk3rS7knC7xdQtRQaY/D4UrNKNly3eEF9Uv84qDf37TIOaM8/x
w7j5AytxH16PQVG1KmaeioCADMGU+QQqWTQMFZJ+296rgt9YhpvXBpw6DE7t/2qX
vN79kb4+l5fUz3TQ8qu1Hw6vccuMF51rfntdImtWzqP3Pyyt6BInikY2KSaMVbt1
jSEiu6sYYfsNEmGLxizdiUwZ2x+MsoosbpxVSB4oSZAYUdv046KHNCVSM468wSJW
WKlivYINeGM4Gh+5jXsuFBpaF+hIPeGimkufqjiYK6wmgYgq3HFX0SPZU9fdanNK
eFGsV7fTDDA+NMJb8yLa6QEk11IJKaCjKCyPtSmq8lTFoEoPqfKro2YkUl3mBSTz
ZYqRoNhRMR/vtTBKWJefPhwxc9rrRDjbbFvKoljZFNmpNtaCWDozPh/mdvqjjyaV
xoRsOIKrWyA/ne34+BjTVKSQWMbUdFFC8hsiHrrUt3CGXCqFqWqgNSxqy4b9E/Wo
DtAKyD4HywJ9/Egu7yn/61bKMgmQZUSnhdQ4CP9j4Mdqy7WOwiXzA2Q+T6FJNH1e
mUrOsEIO/gpRSCU6ckS19q7Ud2bv6bjfSUfWMOsfleVJnnd1K22inavcUK7/Zt56
gL0qB15UktnWGrAJdnvBTvYeVyCI4IXoNDBhWXQt32WP57GWCFTg6L9bhvpJ1LcS
TMJ1uTSc+WCLAFODVzaRaAphlb8XERY0PlIDY+dNHEeN1V6uS0g30jJuir3pLDop
R0354raEwK8yb6ZzqbB4Ok2xN8JNidUo5zxjxfVIjMcXZs1iYFQ9p0GLO3qL/zS0
xeEoM3nGPl8Hb0wYLXq9SvWsP4zw7iUpqLpOkWSqg6WP1ZlpxYflLyK+8yD0wI3n
TP9oNIJjOc9zJbnjEH33vgK8WRspRq3IweAQZ32hE9BwC8rkeS0Rjm7VFIpskrGL
JpnSpgqR8FFdJyFGwLcB0yIaRKlxZnmrrizDxnHLIdBuW2m56Oxuj8zhBJ/fJ/tU
aHLCARQJMKFcx5P7f/8op7QMtzdvaFU5o5NGRVc4A4whl20qb/bsW1xJCCi5LZ3V
ZZBzfiJL13zv48/Cl3NHglyHH1rvCRe1kpcAdAuyFCR3n1igB0bYtKZz8DQK6wCk
0/8Tpg2xAUhmV2DiOZuG1ALxCNL02Lv8v93CcghFdJJXNUtuql5dmnypKNXr+nW/
kNNOKtXuikiPvOMSSgR+A+MBtDUUVHI1rBqt6NL331impDX6dQortEVPwfMUsb8e
/82oyHsvyJvDdzPz+S9KF7kiv5epkGWXMcmFa2DUd3EwgqK2VHOqtMcTSsLOx87z
Q7o1gxvLDgQeWims/4snT0L3XjTDUlZq2943nBxTdrAoUxu79gqIPQ5CLFlh66sa
eVyR62LumnX6TbrRCEtjnM0b3Lyx4ADQO7ock6y3RlS1lkCF7vQ5qH0cB+tz5wWi
xSFF5uqMBK1VzPLipR0VnFCUfSY3iRV3L/TfgPszSAe1V5Q0HqGwy0J1OyLdnXjC
aDwzIOmZ9IWN7XEWkuXY39XF10Df7C/XStV6pggSqKLOBTSmE0VkMit9w53mThTd
5AJ3JiosoL8LD1kz6fj2vRukcerY9Q3pX/iDgS98VAIPVWOZ+SQM+lwO8/7Srafz
LKaABtgP2mY+1NQ+JoXhjzaS3BtPJ2i/GxvGlQsX91DD93WTSL1JsPDqgFSLW2wC
pcH+bau11MiDyGdljP8elVUjlOXgY2QkiD27tNn3DRZN2c5mBCk8tXRIJsrOSN6u
8OQiRZw/tj7mv7C++VnUeG5M6k+rShdiP47hhIAbnfpg4lstIwbvLMcMsQsuyt9J
e1PES/pReClh6mdLseTYt1JkupTg2WBmIvy9iLUWxvz1xSSf3JGktYAY/tFWLHRo
aoAknTBXD7hYHZ4FcP3WlzB8egbQVkeKWLoSBure3SejqcnFZUGcSWfTCYibfyco
MVvAMccjQgcYrd24WvfpteNJgIDS+z/XdWiWJHBns6m8brDVkbW1vNLVP9cryKMH
bVPidGyahIdPZDVg4dZIG6KMCqvwglWqkzxbbDUJ4j4pnBUZq0AFJswEINZ9vMvc
8NIG3YYmBBtgqEC0oDt87n+VcKBWXqx4S4vX3lo+DqZGC6pQ5wY3zeYbUsF+71Ds
rxl/co+lWPn63tcOC7D9oMrqRmfkfF8kSVNPpNGXl4clhG6PfaMECMNmKt1iNXq8
rZcnoW2t93SLIaE5qg9ZupLx+2yac/YrBHnXNDKpbfdrGLGL9D0hhmDN71AjJ3Xy
XJwdotQ3pPvhAEoGXVyQvTOfKWlgMI4Uz+o0Yao23Mht4+Ynqj/Xh4bpzRLY5Yg8
9/1sEMgkSLjN1rLSCBjCMZ297gGY4J4rF3zegASr4VfuvFWGKqr2oEoQYPc+PoAe
lUx/poyulnDVspkbtCPcqeNS+q85vEUQTDYeKyTqH1JrgouZO3W43tNZyzJ9SQ3w
6qyMgWc6vfB/5QVtuxWI/XJKqet9mXWNuX/UUVf/+1wQz8bMl7PvYPbWPTJHcesT
WV3OyQ8xBMVsW2mFBCMnpCNQOD3Hib5AXxUOfTowMkjGOU+swBN8bRse+N62E3NZ
7xutRPrHOEM/nThdmWIIiEHubl9YMq6chZtQAc/kEEBzphxehMcfuUQvpI89C+IO
07618Hj97XQWd8Sm1CqsNHpwgGFIDCg1BGN4PPUfEDTmI0OyAIyLaJv40p5er2jv
iiHJp8kYKFV3aNds7jU5JcxrtY6s3JtkOQfYodBx9i/NbE8zQs9T1wZDuAdArONc
AcnvXmrrgk782eRytFz+0ou86CdfMSxj8JzPn6GORcVJWj7AO9xZSxE8Uy41Bw1P
u3BiDo+eWVeL4k57ZMf9kqYnAx5W1LZ741Dg9/cE43BqRn6tbS0yyonhAfUtoU9S
uYZczNyE+kMP9Vldvo1kJgKdF2IQM0QzbiNAkp1KxIdNDRPO3ucRK6fsfR6ybgkO
bppkcLQy8EogrQIb2I5jZlHWy7BCwxmWhTR0IkcSv9PevgL1qvf1uUmLFt127cYN
I6WPTkkeTF7RYbZLM4TpTzHnKfPQ+zBhlmUOVJEUG1iEmOsIfiW6xiWbSiX6pNcT
7717cEr5i/erdJEeFrTVcVEjDfVXzFvXHkqrA9HHhLID0oZ4gCyGIdeJPbrbnMI7
iA2bko5WdktAr2JMutpj7+bV/berhIvCnDy4aAiXRGp3nAsM4WDcHNuzQOMxTt06
u9IpPKMdFNqRlSMJp4lJBuDh3C/vLYpJggXoRkJMDgDUVh4PhcKl2C7X0BuorC+u
XU05e3C4gMReJYie31MxdJxV5VdyHXvaz2HClzmoJgPHsd1SUYkkm6u1tDbAO/tw
ph78PtsvfYXRytghxUHYswCExUouUCx/wjgw0Fs+KKQfe1AE6WCfVIKRaGZU7iAI
m5dkmyyHbDpw7tLFHeUj6e+0MFNLoRfdAev2VlYwgBbPhJbUv7DNfiXaY7SV/JfM
0Sy4suNAcTjZ9kgt7hvJI2g+Oc0+SNWREIn4jOldiB7EeJsNA3VQAE1DWrXzc1SA
NvcWTJTfMu/QEDM7ggKnFDCTuv9Pt7KG9MpNkKFIkkz2KKoTavDktLmlL5GX74KP
gtcGUuVViNcc4FjEavDA+j9Pvtyl/ZE7ERb4LHYgDcofIMC6F7yV1rErQTDaipDR
jzpY72WzF1bcdZ59KB4rA1RVWeaTkUNmzt2bwhV5BQ8Wks5GwMmn+rmF2z/Ia02m
z877XlFG4DAPDg43/ya9P+O6EUPqvhzCJ9+0IsG6SnYjt3jMOTzL8ogxJ7zLON7n
d/8xaeQm1qEYCI8xZZg4On+YaRgojqpjieQVcosN4kgOgRLu6WUI1wzsrs9NrwJz
jNW0yc4mchYCEqejN0P9FrcacR1NdLrHDHgqyiXGFsj9diBFSr+CwTDx49p5Rbvf
bmw9oWLNeZRvn858sZbyoin4cRNP//jCf0MIOD9ZAWRCQuowotI6ve63DCudQRo5
K6TxzW0gAlEYxnOdidQHX8JsMky2WNYVl7+rki9pcHV+ytAafsCN5lBq7uxgheY9
JF2R7anGSC10bTAeB4kSLintgpDV8DuRW/wBtI7MfbYAdSJBYkxZkz8FYl48vdl6
sPF8xOqh/f6x9XoiG0n68cefByz8TXoGFgH9Wp6RY8ObG+pQkiVsJErML7hOqIXW
upKHlTaqb24QkpEOgCJmgKW8UINnZlXtsbd/fN3jMLy/vHZt/ZHAsJaQ5PJ0qLJA
VtTrQA6iS7KYC5Kqo3Gq2vH8RcXcNVXDeMFuAqrWbdf33JA3nyPjo/4HBFX1yJMF
zaA9x9vLQaI07mOrj0dcRASwOSG/GscIEzzRi66yyf9d051rojuol5OUEocaIr4N
gdzFN5UlDC5Nu4RatgayUN+KTvgCSg1+5afjphGG3HqQ3vB4IaJvTZBm6fjP09ix
mv0ksAuh30OWnodL1ezIAmXnh6w0Gj25wtbw7Uw/m3CzOglQna3w8BFlylylabaR
g9yDFSbnLSmGXSvRSD4PcY59cVjAw7WOFXDNphU/XKwET5nk6t0BRBiOHy+TB51Z
kSLKeOJSN0lobe6ddzGdf2WZ3kbBWYcHB9OSq3dsUxlrewbQwYFnWc6T5SDT+XaM
/pCgSPWlkeGlRorGfctU1hRo9xSa64vijerkSN0IDEoDvCLiz2rFT8nHZcC59hmK
0hA+qSfiStOSDkNxHzMSWM/HEwUZiuTdRQZXUf8UdXKSwDqKgOTlS9iienL/L+ek
QuFBk3yiOhs/AxMCOOL6WkdOGh1dLe34pf1AD7Xj2+dp3nfkt94+IEnyeIyOV7JT
Ybn6LKJF3/ICQOqBbA4Kk9hDD5ABrrJdRgqtgLLGkgPldJpBjopBjdFMg7p0tFHx
YU+vtTZvYkhjJfxznlFHqH6WIU4MkE2RkBJDHKJnEwXkLy/2AoinWX3/WHMiJvF4
VYDOb+QSZBNwpkLStA/kV2dGK0WLe3hEZP8Dxawg2s8t0mpLKpN4032znHvGok0b
XdOW476+UcJud/CxroFIdgvT11Oj/B3qT79FSJx5EAKHVy5gd3bOMe7krctz1hkC
esIFc6xnFW5Y5qt2g5UBFylhpLSMukfV6zWzxRa3+NBC59IPq1FbbF1yJyJVMnS0
jKC5FQ7b1INSUQcZO8y4k7eGvgzgPhymWcZkX3X/VNpI099QgIXDLL6LGy0vO2+X
gmkPp/gBUcn6Nr57bUEZP8/Kut62B9BsLq0s0FU+dzYR6QKHzO+7yNfSoJthNTni
IiCXI3HRYg4amMYncnU2aOA6Fieep1U2iQGRpZQ7vslB5VnNI0Z7V5Yz9kYdKVVN
Ew7T2LL5qLDFFCvLCA7ukCi5ObdJTMrzJ0yP+R+4rit+NVTEUb1+tuv6ohJTHfZ/
vLKlvSqH/tTxwwOgNUOxP5f7s/ArWPVaAK6Gfg7xO3IFtu4z4pZrVKT5NY/GhllD
fGtpbgkaXmvBHh7CYIfjihA1DaHK/v0bSGnxwolefvZY83NG6UONzDfG4Quvx+Pr
srHH0JpKe3rbtuvo3lpzVHRv3O57LHjvblsvD9YNR9lT/W0YafM3zKWSWrr3ecgt
B2dDCogRhDvTg5y596mmrghqvpI/vqmkqZNHIWI69y/bPSxf01RGK/ZEvov1a8JM
MbB1OuYhyfCEQilwGXDvBvFS0SFLrezJSZBVXwBHYNWkGBHEzTv41mzttG0+hceA
fccBo7XmdWiGU4X30SzKgv0CKNSFhMIse8a4ZN29fitW8ord7KknApSPWflalTsM
/DrR52evBK0PYzbnPytWJtI337hN/SCRXj2c1sUn4ElayxqBqNmD+hmOsU+qeXCy
eenNBzNpvrAaT/ceaEh8CAkBXZcI4bwDmqyh5/WQT+O7ygp5FDZknwYHK8EWvzO8
gmxxo8LW9WjrkjGZa8dMqi1zH8YftiqBiPmk8f7yOhRZh9yq+FqGaybaDqjl0/NA
CcyywMzIhiaOhXhKOgdwUNgxw3UKLu/ruFjacMTtzpAMETAbL6nbY2mG3CC6mKRF
RpRLEtXQFQVf9MOWvNZ5CC1noxJUIY1HAZtcWi2Obt9pNZYzF+uIsLCyJv/pEwkO
I0xTqJkDnYEqyetrlxwTw8mFCak2o9HPmgcY2oid5vRaP9B80rTCKyu9W3+OFpeI
40Gbk0efHwpSK9yRS402LyVsd6JoEcGdclhQAz8IFuvGMGqUhgBY6fHgvxpvkylE
g34WmpWRUvaoLAATJeogB2OQXyfgtPrjzDm9UYm2+BE/Y/GPXAFV3KPgVBMyhc+p
ck3VqtQP7DZ9O2I0Moq0oxW5Ktuc/Ha1R0lfy0VhQn+GJDIa53n57tbP561SnENI
YzF4QR8XCrhWHCU4zLcs28anJpuPQUNa7i2Mq21zpJoeLFZD9PdMno11MCwy4FM1
XbmFt7JQWEepKnuejDelquPonI8/Q/Vr7jSMZAPfZn5YBxGzKMr9flaMkdCqX0wK
32aOnvUObNq2VvcuzbaKBPSO/X4VylPuFdh6Bg6pP7THgyANe+baZ5DxSlKxz1nu
ghRuT5N1N7l7alk7JTbkiYDdnm66WAp1SEn1k/e3eE03uEHf6KF+t7z/P2aWqqXT
4IrAUHEKsHaoMUrPqG0jWUOIY83cL4tLZuN49xHawVqBuC6bhJ6PjFvT63U3PGbd
oyiR94kwNxyzc7hO2QriV7ROU+RgUPb3xi9M+corVsEfBwQjyLcR9606JUtPZfra
IiCMLPiNuzlQamF2Gkvw8FUiOZOMN+23CAN1vqQAHN0KQoRtcayf032tM9ulE0aN
5kLInOXXVHspCJuE8/NHTTIaCVrzmUj5Fzi9u3kw4GCHPQrFUOJRYYffTPD6AfQv
MbEakdqGp8zG0HQhvlT5BGUssz87k7d7BhEHf234z1PJeiMG3YfWMZFjmowEB9um
QoSO0KJiwYZoedWhOw/PGRZrWNR9GVhquOLc1QKDkVMprlrlGV2F5Rla2lGcJEwe
X75AfbWzhN5SFQjalId4zct9Dqw9oQUGtYAdhke0auX9nFGN1vuKZIN/D2gZ+0DM
/YMJd5mPibd9iEx5Z5qPlJrShY48c+8hp2Ez5OrWYvK69/YxUDbfyv0mDvtU9j10
mAXarXYvTwM0HWMCoAL1ZvMC2xVAoh+UkoQmqnIcDKboVZ228glpdJB9Gx69tsz7
DF7ZQE+Uca0yuclG5G5CZ3ZwkZ2d9sDSHMy3PiuN5JnXPLB19kv7MpVE7vLhZ+wJ
l1O38+Rr0QNiXyH02hp/DA5A8BLjm2E4jQoO5/HwjAE+sRFUiRvOKcS2c6Hdvvey
pXDTAKqGgWrl53dw+BTP2CsTUobhYUjCNAPIL8exfVjrIoM2TSjIxkYEvwWUwlqK
1GgWcJF2FwIBLHf5VMkbSNUPH8ywo5mylHgRmspBEEWLShknFNHr7rlJnMD06voD
GXoyOT9M18ScJV7ml9qNtjljFPZU5xrQnlREzLEP4xJDdMnDFmMx3X0odDaY+URV
fKRDSj4BYjjht5c1QYmKzwa+W7/TJV/bkXZu3gm+hynmvp1hdPLjFib8fglkvZYq
K8KNVosgEhow3i3ocEB5jhFec8mfw5NtPqEMu5ExAXzi1FU7wTr2etg+nMFWkaD3
/+NJmgC8Np6vtKWjBXbz7ZBgLz3roLqkoG2t0t6wj+AFunBaJwbf8Y3+E0YychX2
sRa37WsRM44G+Tpateo0trCTAPOF0bSnBtEcX9ga/qgbw8+pm7I5B59jUS81x4k6
tHzLelq+whtbxuvjxQ1JPW1y0VjMOC9Rzcp/0J3MCIWEZ+cZZKUVb2jQj5+q7Q3W
ag9SkeFB4v4RNMW9X2JhGDYho4/52pCvyZBnrcujLATVlsEPbyk1pt2r88D9XXIL
bDeOY04pnDvIhUzZ6IzxZ4XD3DuRVBvy4eZva0IYfbMiitwCRyib/PFrq9ZL5Auk
wpC5FXlaorb02wRkvi/RxA5fx92UjXEmLOhkVd6X9dsC5FQts5XuVUZZt4+CGYgN
5378hPWLk52i+YkjVA6Nzo0Kx3rpND0S63RHfLUUEXjJrN63frObjf7Puj//k4Ci
S6lQoMzY439wOPbkgZszIYgLwvLulZfupYJbdGFXtSyOwjjtWLiMTmkD5Uzd3at1
4bPxg47YYt3tqvVst32LgCEeDgistHOqHDubEmliPR3ojAjXJzlrhZLOPASApHen
s8N9gLQBlyck6dJf08ttAV/Ko17JlhR7CNg8VC17X2uabv7sZrnLEHJcBXvLODsk
sOFMC8cCFl2esk36R2IyDrHd182n4puj3j/UFSRiMWeWvpPMiEKiiBA5Gsp0nx9u
AUa2zIiscAAjtwmPdaLGgTM4dmDVVK0MDJHOHXS011/n3y6mOmb8UGBsLA0EIdUd
w52dAH4gL1WzBQ3T0CBlddl5J42UrxXWVRddA4D+hJPSrje4REw5f2qtJ7Dwgehf
XIEoXrCT27ghoRv234c45vioMm/PNe4Ki6r7kqQAgBRWGWS8yeK1QCUcwQdun8dC
MYtQzkr9jxEHpCu94x0wG25LaV5ZZD7JtdUdh2TXcQTMzYRTx1DAe5C8AMutGkSE
dP/MnLsezVjwNYzgwm6Ogbqoq552Ka9SJmas1Oq24FW3RSEmuR2Ml5xNB9OWtNoB
bCNdFTedMMfkKGtWFpJI7S+0yYB0If2+Nc+jD9oFELaNhbi00Op/tN8P4LLU4bZR
Xv1L0t8CDXpJYsCgQMjhz5N2+C1EJJ4NHOseyO7TeL1W/1i66uIw/WtMllNf616c
k+RczzV8uVBOo5JOASKJ4ZGuBE8efO6HVAUU5eKhG3vBi85xCGw9wZHrnMh+77LZ
ZY2hBouAtXezJ7TAwMRCOUVkWUzNBA71oAQ4tz19IdCrck+OivjGgdws0Vdp9rD1
jGShxZvY+KyunwHZad8ZHAnCTWtqEhfptcLItabu9ksdO87X1HUCt5Ki+UNZm0ds
iKfz8mnz7jjTKXAaGI1SkI3ArzMhrK75nDV96LHY9GfEDdi6zTpwB35fcLawyzxm
Er4aE0T+OjSP40Mh6fjpSCVcXwycERaU/VodLM4szrr77vjE/kpUfnI+op5Eq5zo
b81lI1AeoZlZ405vcbXf9yZpdKMZZE5mrQcxo2duCOhh7U6qJXj2urkY/x3DDHWx
9KY5micBTxaoh10LwR71vc1O+GLvQDtz2kB7D+hEPChovOFWzF9EhPJMdT5DvogY
KKrp1IkxD6O1xQPs/sfElWv8PkrDSpHsd5FiabBZp7unnYZCKTWGZdu+zMxg4POc
p8iC971OKpv+pccmaGn+9D+1opNegB57z8ZjfIHhG610ZMwJs/eVTKs5NkkJ8G60
r7rSL47txCL0bcVs2HvZW92i4hX8/O1UVRQ1g1AgbYWfh9dOlBco10bVf3BkIKrP
Ql0QSli0iOljnHlw8dNl22fiy5DeIZRRgrPFQfBgOWO8aG61+acvxpD5D6GKp/hF
IpO72A3OXQp0ZIB1Ky3dUE6+9k+pcVCJ5aftQcaf6mTpLG3gdwROZXOjxgvZI428
uVMhn9eCg1CbavIf9MLksnZI6+P8/NXDQO1dNyQ4lGG5M52NJfVnsy/IAo0vVANf
QZp9VuECqMhSWqCWmbc7hdNni4wAuz711dJ9za+WEEKGLTqjJPxymHt03x4QcaEQ
WIpMn6iCjJ0+xcqv8Pcg9XMMjDwyijYdADeDC+XxLYeyUeCTTY8fCa+7S4Yks2ZZ
8pAaR0EJS15N+9+6J5tBP8dLwTi6DgzrfCFRgS4apHzLEFFS1vpkWwIesTWRxBJw
iHPA2JcCydkFtOwS5QeMjbuf0zG580vP5MuNC2zla2rcJQKiU2AvhO7KH93k1p+k
3nwrCaFmvE8yDYMDOitOF6mOch8M7FQkdLOIWZ+wvM0tfcaQQI1qTd6zYn4j8ha/
om7fJ2KBGgR+zo7RBecBnDwHHFLfik7ox3bEbW3f2Mg3sMPT0bdZP8tJz0mhN1dW
CacEM78kpi7rgS0IXHWzCtG8ZkbUseMIdhcgrZBmRT6NR0++2TyDRLUK3ke9lAP1
Ju+40bBf2bpS8xWEe7Ogqbvi1MtJ1eI8hl/KXImZDm7FlaHo/hqsOLx5V5jFi9HS
LzpFO1RtN30RXsbhtpkeJAbcrpg3fdNuOtQceRXYfIzbMLcROi3ca9ZtSWO2/b4f
CgHNbk1yboRcXcEhLpV0kcPX4v08YEy4nYuYmQfklzjikqYv81qCFa45NTnN+AlR
U5cx9/wtcBIStOIe3mJABUE9WLN5si09Ht9FxWs8tFMXU6oSMSgkkJCaRaZ16LxN
Z2c528YOW8rqS3ZBkzYUigb/uh+BeZ7/zm3xBSV2aeVdYmO0uT6Vwpn7uRHAucRA
sJGQVW7SXKgJoakEKwdi+2zIm8J+4JN8dUlR51LBpCzk7aeJMJcf8Wb1ASIKCP2P
WEJfFDjuXNysTYDkONbY/5M9gjxJNuIhvVYkXWw4uZwr9H9YnaoyjmNk0OLRM7Ig
suQMGBih4MYv/cCsRYJuji9zd9xj9i29DnRzBi/JVSS9yGKcnXSiFnLgfChNdAYY
FO2XAViyzzII2emZ7n9X34D8/enbtrlxAUr+TOu4fKTucsSOINtJ8jx61EVqM4UE
HzHmwDsGTjEYYkkhRHlcxUkCFo1xmEIT54jRlWi6yrmCCwhe+wNLBeqlFGr2aFwl
wDdTh/TtCDY3GAiTUaoYjyhYgyQnhxNYu1hQwDD2VH2OfIThCTLwhSf8fSo14FGQ
AXJcZMPuzhumhv48htXS53sZTihwfEO7t4mYkOO3Wmc0hQ+nMU4Buzw5nIVmJ3xN
M5t25hF/Fm1MOqJwrKK4T7TDodtdGx+DVO4z7/4RcGrAOTCtF3U0WKnhdBkqv/qF
AsEsUKEe6OA/vm/aTFvBhVbesdHZqDz+4pAIjAnasLvzZP6uNA05Kzv6NkbWwYeB
BO1g5xAlyZZteRaImTgz/IVQMWyXn9yZ2KpqbZFp8fgvA3q2rBnfKNDpPggZO5MD
yXb/+UnCGJnBnu98zoRr7dkeuJbjqCM5UP0mylLG5+jH2iPt+ksf3wK28duY4Y4s
m0Nay5ZhgbuCaLnKpLfvm+/1xvVcmxzZQwgZ63J+jB0LUFCjCF8onrolxDbu1HaY
xD9DZ3egvglL4YRYk+xeuL3BBbS2ewawVFQ0tHk4tJr/wzZZ5+pDJEb3pfzUvuwu
szmzxHQpRBqGnfSuV4CFx/p8Vpz5A5o06lDGe/haUjAmdEDfpO7uP+ZTPg9x63nX
Wz2oXl0TPDTYI3Vleq+mIotM93gQHeYujBzjJOSQAC+PJuwlZSBz+MGXCzP8b2jr
maHxXtNBXPkPN5Uuyyi0P46VYfzikNF3PdkXrPWQhdgfoDYrrUMKvCD/F44lHDSs
zsByjhkcli+EyR/+84e8hLCB4XSn0W6SHkFsZ3rDrC5jVYuRQPrIxSGcwMGedYBb
nX1uTl1TUxchNk2ozF6mLBCaU5+Hx4C/Yb7JBEFixiBVVwQSgGjqkWIjvOELhm+j
iBx1qUMcHoqD/nF0twc79j8Tx7RpDlo4xBoiCJr1D6Xsdfu7Cf1cYJN4B4/wT8dq
lxVVabLQWZCRaKfIUGiV6cWI6X/iAIifSbVW2Md/TYW/DA2iCjctvDDaurunqMiW
Kg+8QV+nZzxaKdcjxE0fTjB3YKLAbLOyWWmMmT9yEqFs3nFjt3K9wVh84w67oUbc
BHJYafkkDa1buv6M+5RFeNp3UXCszEBussrn6MRpCVMQr/fB5Et2XTuPjXQEz22u
ZZ4KwEovKyNVKjzgL2PcgjLcTjFoJ9tUUOh+3gQEXKeRk5fQyhxudse82N9FoZqy
DlHIei+oKsL2qgnEgPWoLaCmoZl5/yF3GrFwdBFcGPNfVG8ukxltUh8c3Omwmwpr
+71iE3x3cG+sRi5GgPOT3Gue/3KG6oCP22fowOveXKR81bQIA1+KJngqAxqcJ5Q8
JdrxfDGo00bzoNinet02Pjf4eSJriOa3nqUgPb+LicnQINAiYw/lj+YPbraeHAfC
JVWsW49wCdKYrzhM16qEMCWUwspOXSdYVCfMbBhYIwhlcc4Im9r3hdJnMixn6btu
UOOwL+oKNuPMy376v/0XtMpTW9GMfkwPhVRIa6MvQeA8aQlYhUTxxSVnO4Mfd1va
xdbDq1AG0r7aqeQY6FmVxu60Fuoyd+w9sptBuGfgW+qOsdSVzcy1/F+GUWMNKH4H
UcEU8PcmN6MRuA+4pekrWTu5y3f23sqt51lJt6fUxT9olkV75P6qJoysMOnl0HMa
iaMpiu7/hzLLHcgyYpjcCU1wcmmbWwDt2q6Y1NmVLu/eTiwuW3dzfVLiXP+ySKp5
4tga6vlWn4OPrBG7KkrDzV0byvwVXSkWj1hSyGkZrGaNHCcBb9sXQ9RGRdTqegEq
mkcORNgjE5kU2ybYpyl8VMl+dk3MtD324NoYqxeQRNiB3Rd8wuXEc8Z7yohwUS2U
7TqnrK2pEjX2u5jxprKZAfT7+etMqIwb+wXb+zk2wxroQO8gaqGBaM5AlQNpm+dE
ZIUq3VXTXwNTnDJiBo9EOmlU8/iwOQRzsErSQk2WWvuo/gpep3kGHjRYuv2dmv+9
okeGc3N8/HExuK0VBitbnlTTdZ8AlmZsnS/Qya9dAapjKMOQLoun0d6oR0zkHFwS
KSKeMZZCj9TLAT2HjlUU0OHAMY0MBVTNB9rGmyNKSo8HrF+h1f8Xatzm+B84WwA2
Bbvc1tM8zy6Sz8S/V7iqW4hBamnuWj97a9h0gGLzjbXUC/tAokv2L5gEEBwgdBDZ
FnX73eYFI3eTDxh6NTp8286bLYoR5iJP9mmv4uo6cRm7Oh7ouMO/ZyVoar2Bmy6t
/Z/qqMiEb4EIU5RAnc7vn0yBbRFuQ+M9cq0wGsQjq3tJjpaJtgByrubqMKdFamSu
gWVWezzevM+hm0ix3xi84GOm3B2348WLiQbWCQ0bzt7yG54S031tArV8FQZGcs/q
HfcD2aVeIDigGlC2Lmfj8xtTeyOo3zEk4RzDg8h8HjXfrUbugLdLcR8Euweron3u
n0clbqj3Hvh3DwSaFVTybPRadvtsLlY7U4z4v8PorBlTVXLW0XtIsHYfi6L3a0Km
3ewWZpid+KLGMaXO2ru2THnXhbJ1xoBxWPKV4aTdA0MhMzaBUVG5nUMK+ZmjsoMh
s6CQg5MXeb1LfkdQ2OM7jhBsIZra63bP3eogjje4+SRuWRah1ycu0J+eE5SE//Xs
ePYEyFjnnEQ6ycaZWTCkN974xJw2JzOeRU0iD96/IYDIKZ5EDlaXmfrHW7kf9BfS
V39xSCdmz3P5sJYhm8it3R+l08CX9NdYAh02mrGsXSZrMHP3QS7tbXGRU4kQBKnM
LwjAiHVrzzIa5lgdieDvoOLWLRLLBCogubun+Gge5DMcvJeYs0CP8C93o9mMpmm1
4vg/XIXCltOvRVWhVMQjhSQGXhLhu5LUIY3OwNA8nh1BhqyRcbrEMRi38U/fqTom
LL0BlDsKttR+R2D4yoO+731utjsNxifxZyNf8Flms+kKv2jfsaMHRcD6qypSdgys
1HMl97m8NFG+bK37H0ujNr9PuBu5THk6YrFheKIV97UTqdIn5RiNxhHP+CNdb2UY
sWRvzMeV8qCtRXMyZ9LRfLPZQTOtGl08bbTtx+1tlDprkO2QXraBmIqM3BpXqIh+
TdVJZGRV2smeNK2UquuSBhJl0mppVo0Ni9s8f/9wDCoctaS6gOQqhsbj0vv1j4iZ
JDbmGC4HgMriRyzZR3T/SwuflYwtCKV6O0IDJ/rseEqaPP/KMu2AjT5d52g7QjFV
VCTT8XemQKKFX8rmaW4QjuFoIX0ZoPORpPTjwggVYmLjqnWqG8faXUqKJkIhy91C
/rUISabdTzG3g9YJaQkEyUWRxk45wlZ0PiltBYPweDpNxQ3MFQn1AixS5C1AFNRf
8BpcDjB/zeXFCns5p7S0CacLJXRdYaaLTL+1orqo9wioJnLX78NDkIUhVvqxnSNf
xyl/IqT90Hyl/+7Dv5hcjWsys/uZBaHCtWW180UtGUEwyV8HrWsyou/QQuRAhtYg
7k2ZvU2Tq3VsuttuxfgSCFzA79Yf7OPESSBI4B4EOP11bdtDaniN4/8tUlHpyQoe
VWE10QCxEfiSxv/K5eSzioO46oQe5CXHU8LPPfPlB8ouzlH9eWddgoA5F6sR9kRC
7xnJoZr48kfPT/p/GxT3FPsOx/XGRawE9grCjGHb8KFcKUbL/7tVnHClz+Uo03QE
hDDzL3udMuwksMIJP6g/4CaKam+gWLA9bLwwSkytnrOW9+lXNXmYZUpTMCB+cFWd
A17ckjRBpRPyrcvPzEgzb3MgHBX6/u7qV4G9pUpT6EB67HD8XoJ95R8jSU5ZEZed
1eu/Of+TDuhSAp7GsGMWuxXxUslw+SJ0bEL/aRkl4abhk/Oqb3dA2RmcnyITzl7j
ULTPnuS2LvUJJcTEPzEAOeiIlmjOxhOlEs/+0ggCfZ7RDDkwzZEQjLbtdMISQdzs
QGwP1t4Iss8IbuuNY1uYzeG8hQv21YIZzmSuhUp7ucG9a624+ShmoGuHBeXFJ03a
ZG5HOCrtTym+V/7YBsLsB5yfokxh53NQKIeIY902+VtL+ZmipnaDOvGhVAZzZVAW
OqQRDafh3cf29XaFCmUCbZstviB2qT1JlMm8RlcOYYrdFc1pgizl8GekL238QVG/
uWoxaMYwBlgfyKHcY6r+rdjrIDHksVSTfkiRphloaNhRCQ3v8jY8dNrAvyypKGuY
3fr1YpeOfjmFHITi45nQBwePQPvGNxW0c+wRrXLsHmyb3GP6dHaYcjZdTNYvxTCX
rdcW19vmfDNQI8RtSdvp3JgQDqDt7yQn6fTp+r9CJuqKBzLixHMNHi2+AqajDCKq
pgXLV5S5XMxtfGBLpbNR+zig7R9WN8zU3du3qm2hpRpbe523V/huqGvbYzHod5lG
cZojnrpqLYz9cyLUfScrDKNHfP7DXBN6bZMdadf2KiCFqEFc+WKEXwhfkYpKsW5d
/yWBkGf3PFpwzBvgeVMeKyHoyHLIpVMB/TstmOZ+RvJNN+w8Nzrza6CBQvgt0Pyw
qy2l92jKYKIzKSxticL8Drr0Rt7SOkTnDZupBhLv/L7eQaXRZceiVIjarGjEXYKO
5ZQEIBiPVSJa2N0UzX2S+6IybGYDW5fhiiyc3iYaAHPB9I8AlW1FoW/uvEyAjwO5
OI1a1OiVslHEZd8RoXb40uT4Hk6ZbN/gK7j9PUijpsTjFx71ko8f1u/NUu16gr/L
NiGFqspm4SDzYR9al3Reebbxto1dC1rAk+O5vHH2Obb4sF/OEn971APEwMC5nESE
1F+IMoknSM73LCREglMYIlFWMrGru7tKImyeEcf35GW9RIcbOBAulzQGXlZpcE1U
SmVWqfdCJBbcBgst9ztgZS/iFoTtWWo8CUAGF7/oKE0HKV2s1uOHiPfVZJM8OBPo
Hv4of6ob3bj/54QRs9MtZuWBDZWfEmgfQi/3vhmh388IzxxGUjxkZ3jQcXh2AZLZ
fRi7E611XVb4I6nnZUssmRSFW+gcgEUL3pebORbAqN/kV93fpFiuh4HTkdEOxCbR
o5mNCLLw40cfBAG8ld+9qTLd3zw59eFbk2n70I0LFjL8mP612kf8aMF4YUnRzyB4
7726SM2W/O/yfvUoDeprW8xe9n6FYcmsuIHyy6Zjpp7MWlzy1oIVrHBy0gX49Y5B
QixNDRQC0QQCa1v61zZUPV14lSNCE+uNp+XuBaflbmF80YkTBLeHoWKq7qO1p5L9
uxUJbfxvOZYYyVTDF37qEKZQgYkh2Nf4kQhxVsXJU57DFcMWvaLJboqL3+nj5Hiu
2SzcHZvDMUzbTA5fxwJslpfKsvd7jkWcOImucJ7rTs3GQOC2Zr3RXKF5hW/IV0xj
91FMANtz3UwxgnTebW6UkXzJCx34S7S3HIGEVz7YEkivCoWfDZGpmiwEvaXkTL6O
EpAG6re6QqtAKe4L3vdDAn+gjlZzC6ZA/8jBHeGvY05SXA3DgFZMZgIR8CI6Ez03
/tp2ha8/w0pKTS6ghK1BEG08fMwn9hsg4MltYHcfWQh17U+qBqVZXy3CNOydWCHJ
S8MNQKwYOh1K9dnU07xlfysDsXbN0rWbCYeoEMU8rDRHpWWgtVO02MSyIDJHf3oH
jXPcUMpjyTLYm7uQaE+ENXSPyY/tBp9byb4P66TeFpTx2YXPSnm7hX6ESHVvtiAg
gahaEe7JRUB0rShn3qQJ6p2VaBzMevRmSHm6YPHFVFe5ZXTzbabb7ITMa2VAOi5F
O9YbLTQgFIPOrUrVxtCqwtT2o7O1oETjURjXrQqA5jGXMTUSh7S2mV24nAj2gt0m
06bAyg4ykPNdkm6rfKPV1ONxRIqLA6dWHV4PQ10ce9Tp2UjbawPGPEanZpjuPMmi
fOXr3pskD9taWoidgVcYD/KN6hGj4M2XMApqexRNr5hFGmlEsZlFM2WzJmf4WVJt
JxAYrAR0GBvItsUw1L2uDIWFi4mUaMgrbC71xR3V1bEpAq0C7ChxsCtWucTiv+iY
AMWMGXyOlWbWpExsyihc9QogVSeK4uMpFH2dvPKACZkG9VYxdmY9akDvkd5+NrNX
/6Cu6Hlob/Xil1eaY/HwBnsYt5UZh13MMAMMI5qLydeY1wouP4EXjLWKWCDbL8Et
KOUqgqNp2r7+1KHaLglOlHiMrqD6UDZsXM53j/mPpdRi1VZD+zd9Ij3TIukR24oO
atwfWPl1ncaqnmazH3+AS5k9Pn4Q8h3ePqn0dOiGHs2fpp4eX88fYK4ZfHnJKItm
KWgQKj5uPsQCd2DAfB/Hd6YEwBCklNG6yI6O5HhLB72pdMFLWfI9TU0cZ1h42/o3
8xzgPguEpL3mlZGS+RBQWwU52sNvBEOoZnAM90wUw0h2nPpJapUC1iup6FZZ2Ehx
zjR13zMxqyrRfhB2Ej9+2k8BsNDW166BdjJ8wxDmIPLIamF8AEBfVBfKEtriFP3D
ZniQaYjmaLWRYbR/K5lofbDp4lXfrfLBw6hfpPMCUc3paY1WkH5Bsjb5arpVhZAh
+Yc8X8QQWuBS4QFvof0ethoc91yzLRu/PhX9AAQBrbDffbEDw5nBxEQbIcp1jWsg
a+O64q04mquPauh2qixeHhQ3g113hcNocxwHve3KXspc2bWcKzY9qppcrWrNwf0T
pv9Rabq4HQa7AwMhnyIoX1LR5MzvdltmuLGaiI0IcQ18NuBtaudCEijpzCVSn2eg
azNL2C+KgsbFvgOD+7xIRGKERS8+0sRMESXj2FlFCsxG8OuSmJlBf6ilJWJTFJ/O
kYAlvLFDA3heukT90kzT1HZyagvXK/5oepfBtL5H0ZywYl+Pgo0bsMu8TEgM8Vqx
Gd2AMpSCoDk7TVuufej7SC/0kA/BfblB5ohK4/6BOeA81Eomdt+/5gJMB8YywK2J
Qzi5VDC+6xiywdhL5Y+pdscavvitEkJyQ9YUrHk50Tic1Vppe9GZLsakHXiTPP7p
6KiyWGC+/4vIrBSa8yT6ewVHdLaBio5p7Z+BJeCOdg2SAgE4YlxZLo1zdKfWY2a7
I9ibReK1aHB/A3qFHA3MRxsOtuKxmc+douEpnEMOigg9uxDI65lE+WNfXwaYpo++
6JdeaeYtNUZw1GiH9p0tzH4qwQRv3f2qq1JgsJH0Ln6Cn7jmudRJlDHkV9VPkwqq
iro3rzhuEqLUHeGeQjxv7Hd4MM5/3+tS/pwXTMcuo7UqdSzWngfJMAnDlZCvhrPE
xyyUcG3KQSNt10A50X/nqcFHzgx5BTU3CqPJ9eROFaBm8Vknf+I6AWRG7rRW2yeu
GpvPuRQJDqIpOvqSC4hHgVC4+thIokqT/xyKvednxp6oydc8FF+aWINzMr7MsfzD
JuJIv+CU2LE+ih09Qgb/xxeTdBpLo2wUjoBPr/jMQ9Fvpou3qE9km4apNeFhlM2Q
PlpKCWb7j20inLlVaf9TvS2FAPDowjwEjuOsXZJoAqmOOssveI7sLQPlEWBj1qlb
eDWCPxA2RCnf2m5ZfexlA08R16Jor+7gQOxWwaUNw368U9fnoGyZHHcr92OW7pqD
MTD281jj/+IzuzB96SnNLyjHjY7kAZlCq6c3scF8tvLSlLIMBVJC5xV7VvDplWFa
tD1rdxfwClSnT7uTKYNaB58Zp5tYRcpWJpqit1motwVX1b3H0Cg5kk1UpVkpJGE4
kk1i65n8+PDbR5N3eXmXmMwCcm6OLxx/65kwsv93/kjs2dE9SuR0XlMDFFpGLfgV
/TdQ8TOHuHjn9TIqlCDidexWTQ0Rt1KIxummUPhmVpgLFOFtNKMUf9QlbtZxvMU4
PvL0UkI6SfGFJVSW6l7WmC9DitV5XBRF0Dl6F0L5WZAE9poufFASRVybFugjilYC
Z5J6RXQZBERz7NFX28Nkqe6I8uuXYwnqd3z01E03/tTG9LA+MFEqhtORf6GG+brs
+/DB77rfm36/Vm6hVEhUKRyOFxRFV0fEvY4eGXQwdy17YGtgBDhfk3+tt+emii+b
xtdnbbTGaSNeeP/1NDmGMFMIcXtnS2iMxLjZnwN9260V2+QtP1yamu8cK0UXxWZW
jyQrIxd2xfWZPaQcLkNlvgVtbysndgMQhotpGN1w8PlBEmg3Ae89jYaUDJ7ezUT2
/WmlaNBQmRjvmBaoLqdUhomhS/6Xq7o2g7eYhr+FUEwwpU1cAWPt2pJnTCG50UnK
CPRe8GD7q1l+ilYzC7kJEcn4cotuSSiOJML8YUsrwhmPr7v88EEbqKGyEtSW+YWp
Sot47WatwkR6rxk6GzDCGfjxAPNrsng/GvbNMVPU6bim8JdR7JNmGqhnp+PYeDnA
Dii333jokEtz1XV3lKpA1klcBILgMyiIsly1AsvrGFhsexr+xTyt9T+RRqKlH5ox
qlau0uRV2MCUkYz5CgFi0n9/ElxAzM6LI+tRZVQ6E43j4Mci7xPamVW7vkH+Paqq
h1nZDSmDte4zjj7JSg5wpeVLYWTX+e4j2RHIGcsXfgZmQcLrxZr054YVvLre4s57
2w3os+RmVekz1K6PSPsATlwhzhEhQTlp3+ZblEi9n5kgYkIW5Fw20pDDIVFvYQyk
S62J/cvGVgCiZ0HlImMC6oNLrcCDwWVjFmHeiGLA0bz/5viXEv8IIU3qRU9/Kc73
0CTzYSiT3E2zfaiIGB7daOJuZblE3pa9zugyEIOcojDtJSdRCL9QLw7tMxsvrcai
vQmBnA7qapFj4cS07Wqp1g8l41UA2PBNU9AjueYCzNO8Fca7fXQ/pNSieD5gpcjd
P4N8tXjWcQ7Oypi4/Niul6qpMIbYdV/Qi1vzLtBIK/q6KpFKaJifFhp/Yottq/2X
cqfjmaimSa0nFMzncMh1RhBuF5w/4OUGBhAVTmKQp69n+m6CM+GuX4eb4ZJGWms+
eok7Q6hcbuLEcgiQzIJV19CzhR9OhHTJ3X+W4Gk/oXFUlUqCctDlSceKIRaZNGBw
ZR4epnfWhF5BLyRohX/ildGitv0WXC5gAilZczf6p5VUyDymTCxi6Z5gMr9iws4u
pGtphsPJSH3N86T1sDin1HsPu87OrRj0brIch4dJ8aazFAZe8x+cI5QguN0KSzy3
u0kvQW+Wir7G1Vc7RPxSod8sIkfPBfrLwmnbjdpbbbA5xXXB7Q2PDofEkLGg6k8s
3cUH9v260rDoz1LZiKETMAlWKnreM9UGNM5xmMBoE2qRSCmfErTjrutJOq8p5Bmw
T6kVYuwPegiMEu5TqJzY9e/Y+2VXyp7jQy5Ik3rOaTo9HF38q3GWDmmWAm36lBZH
2CSub8axy4VVnBtSTPM/4PAwzW7Grt1q+8P06DvwhCuQozk1bYG9I3xFp2AoTGcj
hWFp1V/fh9mUWCxRfiR6Ze49UMuXqELz6+0Ik8lu75OSUs7agA1uqdtqa82X5ZC5
0gIQUICw89MNmJ6mrrUUnk6qPSnSkoyFK8fXNZXOJ7wrmoqM9yCRWptfs7Kc2w+K
g2Wu60SCuh2CGeQR903hWQ0RROl+0KDt9flz0XL2UMWWc+6vlLY4ypeSuPOi0Gss
DU7AM0x+UAqCwp4jwVnJnCBoKFXoPG6wtrQgRD28h0rN1bOCICJTfQ7qKRxGeEr/
J5HjdbAPTRKjTS45mlkCj7lxFJ1sE2BJTZ/uvsqOB91f1cZYUQ6+6W4zG+oKwDrC
Tsu06bwAyP+opxFM4sN2JjJ+XgrPpC1uinse0Fss9pFSWj3e3pljeRU30dsE3A+r
Zs3MxrJc36JmenpTs7tbDIXRtyngC5sNGntHPKOCzdiopmHwFhuB49urC0XHWn6W
LDpuZVS9u932Gdc7w6vmQg7QJwmiN2HvAxJ+052ltSAQrqapVn2sCabAG0vU2EU2
+dLoATL8lh/FqySrwfexCsyjGleuY6svVCuVyyHrfREPyDkz1E/zBH0Ib7df19+u
Y7Exx/oUTVdPuypvARW/mleXU40Z0O1n3jgrhpg+K6QjlP3yue8ZlB0h80wPhPpU
eUgMAgxBbkDZXBI2M0SxIX6VUi1zqKbOaKMDLfeCqbe2DaDws5zBzozs64UhH0Ge
k0uuhja6WCc4QUuGtt68T1MwytRCtUPxHTDwsV3XkRth3sAsQdoSYGqXD5MTbUaW
uOfCLI+fHX5RFOnI5EvIYDa3SRlD/4P0c+Feip259ljKsYkH9DJ82WEXLOgkZDBR
1okccVGGRGngtLWxn8TQBsu6pb6hsn8bKESJIbZ3DYpipF8c85rZ/iYpicZo/4zS
9lBmns+JWENqkz1wZZ4UvqDG2y+tn+xdIwadO1atL799y5M0DWI+Yyf8HdqtL4N/
baQynsBEsd5fE94hRS++k4+gHTt7IjPxFqEQKClfmiCA1BmcnAApShShabmAuUJn
OQEwfqde9tFuNxCY0QwSdkH/bPs3SpDdea/zBaL6FDO1Oq1+rwdJApUlbaomatVZ
rlMir9+RCHOl0zDqbzXBXAyQNm24BBKfBUa5epE7hKn9ojjRLmemEy7I3aPCS/hO
gghFuznV2WTCwLoOJkAFxmSksIKQDnDyaTXmuUv8ZBTPtC54/ExfaJOp3QToXlvd
9uYXPFEC+KbowYwmEbZI/csSWK1n4aI/P0/wUFO4nh+ZORG1aQSElW0gAMS29F5I
L6ImED5I83byQS2sRiUU1vIVsD3EAXfuw3KWgLxzrKMzWOjXNlTHeiF6b56qT9uc
b4EMIse06NcJpoZptJ1/oWiVN1R3pp3vttt6A609Y5IxFInHqVVULuhLSp6dWzWO
IyaNwHWkU6XRKlkOnIollHIytpm+8pU34hV5j+gxlIHUhun5yM7w+aYaltgjabnC
XDYc1TgIj4XdqwEGOsP5UkMX3QknDfsoa9PL7MsExW/Hj2cPmfoIPUASIplEcs0C
7FltrGKXNH5xU4dQls3CToJbLV3i9PWXEV+aS7OC1FAxP1xb7L+Y4qcPYH1r8HPv
z0SPaXuJoqFPiXahBfquqyG3r9/FTSmJeibNXR6/WdjXNGJRO4moWEBUdAa7Aez+
BrOEOC0GMgo/P5xIaNcQgnx09yeKZPBcyWJlx93ZnyLMZLJznIsiLjcNPcLcV7Sy
NqnpZzpFhRNNQvNVtOWR/Ab0u4iTfgxortwGckI03/jEOefBnsJJBOMji59PYObP
M10lrM5BRpFifDaf+W6dVL3IzO4KffO/Tlp6OXCuwFa0A/pMtye53LLo5HfDNQab
lHKkMY3c3qtQn3MeZYsJp9ZzSR3cg8KZbT+7ZclRX8fyswmcTM0mlzTyRdBEaauA
mifB7+AGnNg5QzXDiC52U2DUykuGHbLOr+S3fne74x6mgm3qH1q3O50/TzUUHpky
FPdQuyYNXIgTLA/TJ5STm2RSJ0NYlfBUMTfliOdz7cbl6jRE0cDqJFz81K1ybft1
mw9UpbZ/ET1MowgqojM7bW46Roqw8/AmSq5P4OSwoceSTpsK7pWCuKAQwk6yU29d
gLFMJreLSyxEXTK3qwVDzlKznUcidh5Le66g8hV9jSQo1fO6FcOOnJsfSRXAqo5L
UIF9gug+omxAI6t04t8Op4d4H7tjA/gt+Z+Y1VlzDFILZ5QOy+fi71iu9V0ZFco4
kzfwovycDO1ixz9/aSYMjPtLS7tq7rR/ZRNCus04OKn1p1OP05Mv+K1TqAdCcPWi
wIN0A/RWEECTMUIQq1TXmLAAhy2EHUTM0+tm7hq+RXO3wY9Rk6ZAastzCfm5I1JG
iVFkZUvJBV5oeYgxZ2bTowVm1JiJVAuimoEAZWqTOLRymyCsf07kCMyWE42BTVg3
oTHPeemJyz427ynp6yDRV1pCF7Ovc4iIHzM5vFJZtMkjXFF9Ezjgw2monMSNMPor
dr2Hs9rIJm28+IUP4Mmy7LbrQUMop+yDRYUUCg4G+gXiknl+LsAH5J58uhVJlaLA
uUn3Q6cTdhKGvJaFf7FrvbGuQTiaGBvZg3E8+OsGr1ckdVVztiM7E0i7zSe/QwpO
1YPwKrYkpyrn+quOXYOi0OFcRjszAGGmIyq6egBOlTz5U85DG2uNNwe31+EN34f5
WXz4Rlqk1pB347u/Y0k00re+hjJE8yHeBONMR5KpPSLojdHwH0/aWxLZb+jKJcA6
wmcNbbp4Qyed5MDZpMbO9en7JcQlbnfr5wpF8wFpQiF6ez6e545Pz5oPIy5eRK+K
T94Mz+420p03r14aAIDtj8c0noe0JcIej4joGrjwBsvK9KW6PyzuI6xOvPc8+UK6
ebtTmL2Fr10HYyv28R2r+YbDbwJhO6SwzauUC3qxzSRrUR56mvuyW6/sVvwoVL7b
qJcTH7FJtZlE3iWHPwpDORArXEwrlDGW6KgpXTP5BpcQ/wPPe01tu1dVe9C+ACSZ
wxhO/JcuZhkaqmPuVzlOtCq/aNOH3mUSMjWDA39AGnr0ab/x2CPowHs18JL0q0U6
E7UHBzm6zsEPDCuHWLW543WBc2VDd6MyF6fQPhPROYnRQdFOzz2HQ1T5Vx/oAwD/
v8x6Mosuw+CFtTIZyg9Xq5kZyRcy4K90uNLhmcF1xO2Db+P2ZqMi2lN+A1laAde5
eLTQD1vek0qNbyxKE3wwkMWnJd7iBj7PRMJEj8lsfE1NGDvnQPBMQYKOspf/hpFT
DZASyntLq/owrvhkYMlXQglFGUe9W4U2lkgVCJB5sg2p4azYdMtFHLU1CeJuI6lA
mG5xzI8BFFbakr0Y8OkXn1aPaoepi9l4+j+ejhGfCAqP4fmYXYVrteeBgMDNv7Vf
4u8C4M6EMLzqJVyirreasuAAJWyftMHe7As+w2zPakr6GLSTg+aQWpN+gb1r/mLf
R/uIEQj9YpP1ijfplJdfqPZLbbt9tUcYIbUW4+sOylkprpMl9HRabsA9CPXNCbEF
y+2n7huyDRVEUPyX26T3BPWNfzU3ioqFgEFUcKkYiK94WNMZkLDyOivNsCS231Gw
GfSXqaPORn1upC2wr/aGHP1cM+gm7G55eD3vD/69AKzg6dvTJkOROkQ3aUDMQLiz
gKQREiuG8eBd2WK1Zv2Zp4dtQS9OfuRtQN/9Bxa8CGlNrFQdIju/esDuIrF5GBAq
dQBV4zGXWaueJDWSoq9/LhahPNxukFRotZYtviDzcYh1Kpq1qtM13vN6yJj4kZET
+pZwoCyVDVKmrZA1n0KaRH3CLbx/uNo3NzDXO+ot3mD1YaxhGlTWO1agvAAfFnz3
+DpX34/Kr065g0kfVgyfIjMeB4FCOy/O5SaY3YxoT6TRaZHn5qwp6D9/YRuQkHUo
5C1DtDKjxhiIX/2GRGJ5dtUplsYEql85h+6ndYipK1eTQ+NTsEzl4Of7X6iMi442
g9JW1IyU1YqHETqKNV1ihAr/DmVhF5T11/5mzP/p0TzObqBv62mW22p6AFi60qUN
39oDsSz6NGKiR45vxZt0WAa7b+pL7yEvHTs0Ck+3oAZ6z06Q8MzDYDNeYbliy6eA
UA9k91q8UYNk+v2XgSRjx3AvARzr3EGCHjMJi3MHNKtH/4zUoT9m417dsc46DV48
rfnbNurxIk4D4J4bRXLwYX3q+ecBFqs/O0PylUH5b4vdpCP1DvGz0QbAQmKBEXOT
F+j4gBUNhuWKyyT+hL/Vf0gh1YNBmpYgJfJ5MUtLw9eMJRoL+R06x/QRp3ezI7TS
Ufb0ApFJHdOc5xAoqHu1Htwk2Re20GaZdHUGBwRBLvGiVaTXb2fsXb0tcWqA9hhK
C+f9F6DHzvqvRcbGNpdfEztuu+GxOcnYFFaWNRj0LFDyCfx6Dq6mzgOqMl34SucR
TUO0dkS2bXVryaeggPysoMPgWcXuZeT+KmQt1GuwRaacQVzMPWeCBn5Ru1q6+FHr
o1dJpUpddJu25GbtQBkO4v/LpMJsJIt5kMX42v625n2kTE5kP2GlkFkIuphXbA2w
NjHmpRzAcQWM7JCTxDm7GjT+nDyd8Z7dzbGHxD+wFw4e7BFUmOHeCcD6izzAYnSu
jAvwH2amMpN2UzR8lLoCnHfHBvbAg40clJ99L+Ek9yF/IjZhJXd6E8auEwXfnK0G
2L1g4zEooHHKwVxuBUmCSCVQAuPApjRh7jeMwh1v9zGxXxwFmo9adQEB/ueAH6+X
T1wScC/p2835gv0r3mwBcM6IBvS5ko1INiZ9dzs1tdNENe6orFhfN7jL/1pnVMlp
EK6q7IedshAcoFb5CHLBFcKO1fFts8RxkurmSulcDHApnQMzYI4G1N5hRNex7dST
uC01CLgFmZJMJTzFtd3lRwutKEOY5GyTyi8l0xqgXevoYU8ty+xmoEExP2Il2Wpj
rTI16RnT4q424kz2txITgeDsOznN+ln8f/836TVFRF1j30Af4ETVRq1pqv50OUe+
zYnk7JkKqDB4DnUUy+bHbBLeiU28RGEQ6iu1nm4XXmtb2mcuERPDvfuTKNZMqE36
MeEk8O+sHZubEdMqDB+icHcLIysq4Gq6sgbszHi/2VhJODBn6qCT9Wv3NGOhsZQU
Xj0sYLA6IfU5rkr0TGykM8pJ/TULDNng2jtXG5K+xkaHYoXc5XQESUFFm8oanT4D
64XsUjTeL8r7jTzUswkJ2gyE6iTnmtyhtWtDZFFjXNHFzHLtNIN+P0vtEtBZYSBt
gKs9oY877KncgehlhWiVUvI49yhPtNBZ0mbCx64BVZ+BAw0AwVZ46wKDdozEq6cm
0Cn1sNk67UTiuc4VYFf9p2yJqoM/cBFvjGDCzjHTNZGhlaImuoSbq4NyMQZ1u1vx
urp9qA3SIjDVcxzGWvHFGzkmYEXqbPa01qME1BDAT9OO4ftcCdSlsgPCtaYS9kX+
40QpuNzvI2aOMsH0f3/z2Z6WWSrfvR+KSKGYok4Lda0+N+T+LiB/fBnFCdSHK0QW
Vl8tbDVc6wV7c1mElSeuht1b9c3KrtC5FL3kFx0IombMjgfDy38jzX2fZjpPyggT
YikivBar8zZGuIN6AQ3Euj+w+82wnZ+Euo0x3q6DrHZ+te/ztghLGIV58v8UXXhI
ZcmrNujW3PW+22KqYKD//L63CNeUDkdLxjaituFj7UGHUBaTGNsFzhhOtPojOErJ
7bIucgIAXvpt1Wm8851wEysJk1p/LxjGnazCt4MlSxOqERfmyT0B3SBElfsiAWVJ
X2NugwQPJKJwkT9ViZoAv4iZH2T6ExqWtGMWCMzMRhAbCM6sNAUbVvHIwzuwHP8K
05Cmbc3HRS++Gszqio9YDYsVhAPio94CfbPZ64QfJh7jWDxl2EgyEZlvkINtlAGE
ikyzmWxn3YGOFdu1hgydi6VvLHJta5C8TCNWG0UOlZYIzdcEs3ufHY48CyQBO1io
jDrkpBCcqGLxgGiJoNCw15e0smlkO6tc/cx3lYh0UQ6QZEop4Y1Lqw2BhelRZia8
DpftmAbPY2cKQ2VqUlLd/ivQjhjdA/WMlFlYyC+vMmift4K9D+EqWxmTbEjn9Apu
EpoulmGMPNuazOPS9IqRBhpvnBM1Kk15+0zqhPUkYYW9k0H1RYo6QJWYjINXZDWw
c2QMNEURRGhfsHkCBH1SO/qrWC83PfxMtRUD5wt8eVB8uXbn4ysHZdeYqzIjnleT
YJmLeOIxjG2OhwilS+WM16quHYMPuOMPdIeiZL/IB9Ud1PNd4l+blrYIHy9LmVcK
KJPyZfM28jburFE5sP/wDl8iMdSzhyQnrSdw8ZrD91avqocf6EMOzdVXGPi0sqgN
DYBOfc/67538HixCxDJFgvNbwoGSUGdzQJYXBmMDHNdm4HfaCs9k5vBKxF7Px1uu
gOQBlDtpWJI8BcGr45R4uqiHlBJvu28LLW054ztXBifG8aOzBw5wVug0MFZw3XgZ
MH9OuUBD/7Imv5BXl6saszPQe2lRZll2zsmvHvTG4BABOFLUtwDgfOaWmZpWzryB
xe3JltZzMyx/kAyDskIU4NTyT0tGQs+Pw6yxiYVIcEoy5MPUJsI+IZSPSqQr5jS5
iyIYm+iyuPwpCZ/sUn5LWdKfwqvXzIW/q5rSUy2KreKeTSLW20YHjj8EeLBxuJk3
EP/QwolUWZYyOIIXJrRt+UriPyudkdpORCWpML1brtRGx/NyQ4IqFOVuPhquS0nH
siiZGz3FiFhBsxdGAZRnh0Z+8fcKmm8O+xehMdq61HER7l8BCwmFsw78qR/rGYyA
oQyZUNLbg8B/llIL26c/BDoXe+BzYarfduv/7g4RvkoU0434RpnKtCefF34pSXM8
15igCntCKnyDRW+afuHP8S1tWrbJ3hZ+kMUaAzZ6mVPpf5kR0Z1dDdTz842seRRb
YzNrOxXldT8i6ZQ2Wgp/74fMM98UJi6GplRl/mTTqYCD8c8mEIZem6Gw3qfX0xdJ
sEllkDyJcZ+MFila01CsIpsevukKDhuZ04Krp5OQFvHFyAYOQmUfRIcO5cMip1ml
dtH0ah2v0RDM3rabvteW4uqTTK9xOW2UTMCCwyMiaYaf0wk4N6ikUeO5IXPz/3Qi
LcYGNrZ6XcBv3IWTaCslZ5nXo6H5goRFIfacaXFHNCgwvzu2K/1+gF1wzPfnvuMF
kqsaziA15qKC8zmUD/OL8na5yLhazH/6U0wWL6J9TpqZI8ln/Unkne4AM0DJrLAq
mVZrHYRfxd/4enk55nLnEwepVtxY0GLvi38Iu8kSbaXfJtNV3KCTUVynJo3+Dyed
KySvo6CvY9ydME4P19wbAm+MOn5Aj2ASFN/+jRP5VIjD5S+QdRjKed3SN23apvXH
Hvdpzr+ITKxTUJWxHOjyJsV8vyIL7Dmk7hSwUPxfjlqpqo/TFhr1qqxahZ+jrrUj
L9JiGKB46dNdL6D0ZP1Oea1ozi+/4wkYYSU1DiMoEHKzkM0pIhFmSnzAz4EE34PT
oN2dCPH/atDgJ4fSA7nctDuy3Q7hw+Xf0a2X0loWAYCAUbYcpAQdCK360FavSXkv
jLrtKZI/OMHMQez1YQ5/CALBbnnpu+NMUNt+WPhho4mApqzdLXaFXN/fRpmMQ4SP
OBmx0HzZlCZEpbBOoHrA4Ajw3nFU3he5L9Qw5eDniZ3wf8w0t8e1jhOVU2xkE2Iz
JIhQZe+ItZ9DgRCkpgHpPSzQvxQkBBUlLrP968SKwtymGPqzLaNlXtexIbxSKPqp
N19cHPFRmMHstgh1KuH9XfX7BQQNhaeH5Dc/enPLGAO7Gph5/U8oDjNkRSBMwA30
5xW5vcl0dYfPKSE6AV9yI6japEUqkY9Z0TNplDSirds/icNmTX4bRBlIGwmJmnX/
XufS8HScTf9DZHR2AWFfaR/Wxh1Zx8bHL2vUkc48bQ4RCzmnMggad3LWJ6jRE4wn
WOECZdsSUavhbtCQPA/rDvIjzXXwqg58UTNmbfuQw2gpYfoOPlABnd1y5dxfI+6n
Ea/nVxnV9RujlLNnWop7Jbv0VPNfWIzOeG1YD6HCp4MyukHZtTXFBzVV0BxEU+A3
CNHLcEtIoX0mr7sWv7lGyfOnjPjZBz0TzlBynVTJzZq6ocTuSSljXPylp9xgw5OL
Df7nc11cIty/jWnJhMGxNxrktmZBN/0fCTUvnxfFz+oF3XHo7Hb1VNFbLssS+bBW
0wGj91nbMaCK9M0PL/Sw3JEpbBWEAhdOgcR2p7ZYCJCm6AldaCkdldbTiJhOrW6k
p/lgiUBBXqTrkFZrV0Qc5NyuqT/rdqdp90QdfIXco/a5IX91KC/+ovr20UpKQg43
Pqngn7ukykNOJdPXfHoBisc9Sct8NgsiJtBqAF3CuCS+348tANJBzovfiiMqH7BS
ZeOhQVfTd1A9WOl8tN5GHZXflS0RhqYqE+Yyhl8Gu9w0MOGvAypULS2jlD6O5h6p
jbsli+Exo1LQl46WbmzUXWpoOZceyVu+flVQu8kVwYdBBOKdiWckd8by8IHiAV71
t1uLk83BQD7zw6zjigADb36/uBXAANxmfdrt4ipSu9V8v4lS2lkPNE2FjJz88ph6
e8S0gVnhFRdipwIZaP9fwemIucBtHSOCj1ZO4WkSoucnJhlXSNWn3cPUxzDBaC7l
dQiTTAlIBeORs65vqJzSZZxMkU6bcKio8PQkJXRCNLgnM9aEIk5yYoDtZtT9UOaZ
9AHdm26/Pnr698x9nynucNgqwr58gZJF/bkUWXnSgv7991v40qhq45JGy4ZhvpHG
xU3BWl1szsWL+7khe1Nl+2Y0I3uVgVb4kqataXNOj6AFE5xS6xYs13yDGk7S2spU
8gdAc8Z0PhBVa9q1T0cZ64J8yJp9LuFl/M82ONKXD+nW8+OdysOhqD9XTYnLzZLw
Z7NIysadeAGxTS0l5KQxhCpAVqSQ/BrUuB1xdLWpQTzI0MJTu9MgrmZTznLTnzPK
mcVw9ZG49qCjBEqyF7YMpQWlxuCZSgfZrubDCEaaBSFLOAV/ypR7MKaHj2ivg7Kk
pbddlKnKfx5FLfwQM96mZbX6oC5kvm6zDsQXsxBAXE6d8qiEx5oCVOMDELs+njwr
vATX7KL3hXEpNGhOvGYINpqrRUmLZ8EaQ9MNKlysNUXWm7Py/JrFKWpQ8i+5SoLF
bCMvC8p+TvU6XXK7+Q7TIr1YslyXcPWGnq8VVS6MRd0tJ0Ai7o4diTkusAnslxYh
QdVLB7m9DuhKDP+NdA5YRLqfGXZgmPrOR0nYjH6DCqKiKhRL41BXj0mZ4F4HTThz
O5HxHb/nT4RIBog1Mc+1u0qe+Zvc32a6DL5SYOf+h36QIA487OujH+mWt/pYg9Q1
sR+WBwR+xVRS44PYqrK4WK3+s1BHmdfncGkp59ORZ6C9kVsCipwgFEUQJk+7OncE
T+483Z0MMABlWQPBfVWbuw5RmNwmm/r+HGjYKw08eYm1pBDpVaehbL6sIcyabXKm
8HAE/Z9/yUd4EbgDPJUXMiCEr+rvsLFY8Xbmq9KCP3Q2rigyPepLxQzasYPro/eo
/BcwV64XcfwY5vjWHK/12IxtNvdBmvFjcF8qTu4bPzPMxVg8WZ0y1pc4xt0x95J/
9UMMmov2h8KHn/wu+mGMmY8BrV3DjLyXz2625ONm91LhlM++fIxN7gq95boRmltC
AEnIKd0AigKOoMYx8Gjn65pZDzgIpQGExaZxukw4YB0w12Q8Vc86amX48jHHjVyZ
mLYTfCYE84Tx+AhbPlYjVKKqU6+9x21e22iyVZss/Y4BO3vAr7ccTnxX1oBKMA3X
gZxQYwvrEEBJTHC3Z/iaRUffcIFz3exnCBMh4RwMko8Nm7z2SADw+EDXkCLd/rMa
ArIEj5VPxYdcepdr7gOddiJ5CP/MQJR/Jf8+rNaqrm8QDfDIcIrw//w3LBn3ZOb6
7nhFoA+lOMg436AqRVc7LlUBlL7Q0Q1qpIxOHSjIGyWqJh1CIcf7fdCAOnhVBKdY
Jyq87PhnC8OOTonlzC3wfFXfTbS/NaoMkcyBlKjWlrAYdIEm7v17ApbccMoGaxxJ
dRjuFX5Y4BF9AUswZCrbJR2nzCf6Bms8uZATguhm0Lf5A8qN1nQbwFpeu5Rwf5P8
K0NvyBkJZx57lwCcR2f2lfL6RqGN5her1WBTUZ8/DXtmD2e9UVpC0olItO2FKP1t
LqjDSucIVaEXLvC3BWoSTIT77hQVQXev703B28T9NkPbJWKr7htAbGcu7us0qCL1
6RJ1fl586433NmvmroFFiX/tQVOOZgTQVePE6BO0xh6khyA7QJkfVzuKXK5tRCSD
5xY/qKYGLLsTy1i/ot/mUJuR7ELdJzUs4E4z8yjAc8YozyXsQKhqGc3oEt17HOkj
GTIqn0Ncw6KVr8oS/RlqBxNrXe/nbnOo5EEZ1hyYn8RAococetYM5ony/iHyAiEu
x/8kzkXe1Y5pGgad5AHxXwEXM1WZcE7ANzUu7IDdRrzVlbPCrWCJ6zqMKJMjSjSd
/UwGQr/pKP1GnTufk37BVrfA22yFfO/esTioAc1x8ckD2YpAJ4Ngh32A2pdmmoBA
8rqk7hgo1UqtvSZ5+vqB3CYHKUn2PieOJ6B7VIhpkK+Wf5mIUFG3WURhpNbqfD/s
1v9PjcrM0iUNRLPGtHWEjuez2/MfAUMsuvRMx48OGjj2MkCEDDoBDENxzRoV7+r/
vh9NwBRE6ZwvvCtp/mUCU6LkYfwSRq1E+pK16iJZyHwfAfeYh4+X7SC7lWJc+O4t
9gDY3BhIKciUxprBhvxY9fm5C01ZcrTI5YyS91ebNStiqZpA3quoXYvQGuHkp9hg
ZeFkEWLI+fOepUv/Rh3Nn2bth6UFX1uMaHF0/o4zcD8wvKSXot0hTRtHfNA7xEZZ
QPjScul2QJiErZyJFZTdNpHXD5+RC17Lis8NXROz5uvt8WCyR2n9WtqVt+gmAQqn
+/tRuwT/MXNspyH8C9T2jlnz8W20We0HmrGsBEGO/5fuIrqPCGNtzY5/sT+n6Wow
/Iei0eXbkERVPqdDsrqjmMCvMZQF6kQjTXUz4M2YGcjWpyItFxysVhXmAv1QPG7U
z0vyA7cQi662Jn4qWxiCeTjrSAnTKGo67c6Y2Kzx1sE12i7qMRVTtcBhe6EbLBro
vEQx2NptuDiDEJIcQ3adY5AcVpQvZLUV8tQCNwwk44Ol1i1KGr3rGz6i7QfIZTAN
jX95rI6MsEWkchmkETmX3mgi6kMJiW6B/8qsPQ6CRx3K5JSaDjYecWru2jh/tHGn
BqPuNm5QvP13FA1s2b8ZisZ84K+2+EfeoH+FrjZNMRnN1xKLgzP7kTb94kqI0BkN
4UNd4VGHUxk9gglkswG33MN2PWZy9WOuYEnu8APBpxgkMLSsY8ckCK90l2NDp/Yh
uApZxTYoErrjnLCaU7jcDwR7L0eWSeKsFPMTuR72LGWXmJlQSi2MmNNqB7JqWzUq
kXOb0GAhHlhjh8A8Whc9v23eUjBUuaGQP/CoGPPXZxpe8j2wgrP5EJCowQaqstZD
dKUzMVxPD5hCm27kFJt1oxzjpQWiFHwmS7rBPkI1jPwuF2yiQ5ANd+5uRCbsoyLj
Vytv0Rl3XAzsbh4+H2iJnBLY5gSrAtzr35WDz9Dc0evwrmMMp6fcMxHJgfYYUD+O
wRTcRNmASF+CprLGO94/xCbSg/yzp2oZbr3T75QO2RrmsPVPo2HxNHn9OHDUtsYP
iRHuWYGokpwMIEgAR2/rqsrnnKz70DuZO9E4RrNdQ6bG03vD2opM7bEZ+qB9vghI
21xVmHnOUddyWCNex09DMPIkXhb8djBTHMldKvsAclB7d/fgeGIoXoDlYjAENqpZ
p//ljGhjPzv2ODMIczFGTjnLpmXVML19T39H1Hpgv83WKqKjBixOKnuef+lYD8Sq
SMtxTAk7dOYR5kxDeBdLq6QthNEMJkOAikibOY/hSHNNCj3J0vC69AgcXovzUvD/
DRZFOwuDpsND5u47O6tRh0aJ/TyeT+0QEix2cSKW5KOsXv0oTDVNIl98UMo2iXNM
N8NGdmgVcVffPRjI+NtMPkgk2SIJIM7X6YeZw8zF0O8OSznntM27W04swkOnKBQp
ffSqh6fVubVeja7wrgRrVt5UHsle6u6zyvb3TDKY6FsX0JH7r3i+F9s5FJk/UvhG
L47EkdtuqmAFafKQjN1cgCilojuo8vVfEwqy00Hu9q4ncPA9C8mLJbEzZ3booHtl
YbXTF3tlqRaKTg6gyzkJRq+nO2V2/qUYZHxaxxBMxRSvOq4BoaCxCPWGvqdnxXK1
9PaYsYWdaoq91YFLlRfvx3gZs/U37r267kZ+P+pboPs+QbAFbl0Sj+Ruwaq1P8QV
YRpbRa7vBliZuhtBW3/yAO4m706TP8QBfqha8Qr+t1rOGB75yYnqV0VUlyQEQlix
FszmG50DFSoMosM/4j2ffhyDouXSe+UEx+hfSvlHeDcALg51Bcg+01ooqCuMHsps
dUVeDpdXh1XrlxUjJMEWZb/GwVBYVvye1bmx9QWV9N7MIj9wj+xOJAwh9gxKOiQl
YT9Jx3AsqAWRJs63fuOxcxI2+Weg3RHilJZHZzfCkVgI1NqJV5JsYIHFh04I5qiZ
4MnR5VGuxI9CMZGOKPf3rG6aUDkDwu77VVLobfp2OE7xPyZtH2VOABSmDe2/61Yj
fuIKHJ3MTHUqBIT44G2CjJE5vmkJbCiDzAgKX4bdSXj2udHieonqsoHSkqIXYHYv
wrd/sW0msQqcwLWjKtRc7oWyxgnx/RRL0l1QUyPxxWcphM3s5+ueBIFn8t9KPWVm
22k7qhWWwOdObVhVXuDzwG5Gpm0AFHO1ZOLRbH+Eqv0ocman/cLoCKUX41vJDOpA
b9nOsyeAM4fyMX4QjPX/Aq9NqNoTXKuKNHxN2oSkGh9ZJiy4DTsD5PrqtoPTkuIc
gegUwSeN6XrGiAAxH4U81tfNqyPtcL3ZzTz9IbvzMM4b1dtBGJ0LGyI+kGwXvemX
cOpgvke1G19tIHVemoUiDGu2idFD3iR+YGgwb2rzA8UwU7LRkd16rUAZ29Lu9Te1
F79LgZuMPH8JqRGyCvgYbKQu9hSIlUHp2kdvHSFpznQS/niBT6sviWZzCMHTNDEf
bKdz9O7J8zvhrGe8M+HRwelFzCHm/RHQJKzKijeum9sW9T+a872b6OTgUtXoWXLL
5nev0tEaIOOY7q1/Sk5YCbyUHBFJoxhO1nw10aPD8Wxr5vFMJc6nEmdvgQcVBHfu
XiY1y8ofdVGZOXIYhT7aekuoUCyTNPPsSwgYagPcQ3pHWZqHB0wjKCAxohJkuOd8
7I1Gmdx9Ogmdz3Y9XL1Dz79MIj+EUmHKpFGo1945jggbsufrblA6qsQF3fOLbA2w
AOip8LoxO3Y3QZLoWWES3/F1uuqAQQ5ELbtS4Y6q+jUz9mCwf193H9W8xDKu2X2C
9M/w3lTrd0or1cRFraEYkoFFYAYakG7hon1b1ScORbcaxTdofXaVgSHchsvBysnw
sAllosOEooMff7MWzZMGCceGGb9nUxMdrPvXAdML+pniprBYTuKF3uWyd07qAs/W
zd6GRGwA91++WoB98jku6DkgGlIQc1eriUfvYrrpboeR+5m9v0bsvbhFW7oMkbw6
U9pNI3FWDWgspOi2eu4hfNU/5dG1dEFU7l7C42oAYPuOfbuRk/KV47rG3oS5tZhh
iQQ2+iQyhrNjEkcBRDG4OSMntW4MEvsvcGnWDkIkU94IqBkHRYvLbkadq6ox+5bf
2+rsuDG16nknRwn6uFAQlNQ477uodKHOwX2SDSoHc6AhQnYhBsGyWjiEeu0tcPVF
//n5o2aePQUX9tTwLxStUVB81nbvlgkcy4Y5rdPt+NquXLDAVqaLtnlBEbYNKX0C
MW1Z2tHldnNdTmUsg6fqv+GasuO6Jx+C4NwD3KRoe2EIsl/OVieMK9GWBWmpfzyd
pSTFVSyE7JS+7L7eTY1fDRK9TzziY8KuESjqjnJ2BFspULR+//geJ5rwW2nNZLKK
I8GPDGK7eRCGkWmj9Eru/jh9AaNd7O9EcvDsvMMh11aUdVAoot01VVpX8jn7aA3k
vzquseWjSlfG39QURDT7moQ/N9nosgDA9DXI/kDBpN471sUPChA3RNGoNmC2ldZZ
WWLZjY2w84/JLVg3MsT4FnznYAd6jRy9ysGJ70I5Iovu6Ex2jkhuDJ7bMdQv0VPw
D5/pvq9shBGdN92hUMH8BorItBSP9nqdBXMqfxpMy776h0+V9qVhq64iBHtxeO5I
Yh/T6v5kQuYvd+UvwvWRv/SBWlTav8DWFn3hchygeaXojkalgGPz0IkFQsasp3N1
IwyeZ06yd10JSX10T5djYsLMSRctKGq0orBTSj6NTI5OHxUJkGHmjQ6f4XdW9Ubx
HXxf9x4dgeukOnUXNTCi2lDQ2oy27vy8rJtlAi4k56weiYzFyag/b6gUxg8l3bdc
YWXbsPNEPRImqo6wOLsy8oZ8ymzpkBFWHnJyOxzWiyLr0JxCrgeTYpAvVPM7Vrnt
f0zGRQGg19yNpXuYzSEihgaDTHESpCxeYDs9PmRhYiVI1tfvpqEuARkp68g2JMfo
fP5uksAhm37yIJ09tc6FTQhIIomD9nXd/zHbS5QbTW6cDjb0HYMGvs0LDYdly8rN
DejpXYrvbmdLu4uVHoimkeJU7wExfvrVIA6mriPgHWXk0qyH/iZ9uO1QWlGrcr/5
Yov1WojEf9+OsTR4/ov7N/o/1jQp24M0CyZgJBeuQYwfDonw7LMplGkkpOhFlLRC
myTyABMNzlUaYVESNAU4vduDTAyxA419ERO7DpC2NjHbP2/38h91NGHIcfg3ebQf
FUErNYBRRdOR/Yqtp3g4vE3kKKpAjB8Ik4t1NvBz8cSH+CB667SQR8g9KmWcEhvo
PGoxGKPxRh9YKVCqawXOk1kzMVFOGZZ7JKsmmZJIHrRXklo1/7/FogpO5m2BEIem
qnP2fDBR7zin7/jVw/9XuBNsbQJnu0oBZJLrrndaDg1On1vhtA4HSp/eTez/gS/l
YI25tV4LaVqnxa1K3rf4tXHcHnaoQmugqMcfxVPu6P+ota4kHsteOraafmelLJ/T
mqbUaP7ujzbvFa1NOm5Bi9ixLPnEdE09PKIL6zbRZdYCHnQ52jyC3t009vQS9SCF
2evC+SLP6SJoHAW8Tai2NT2xqPjJLbx/THioIuHpc2FACHpPex/0LbwUOiV5tEd6
Ye0wX9Am4k/GpTN4Vhc0nMwldlgSUXWXQ7faO4RsaHP3rwLFGpsYYc2VjtZR5ufY
GtyfCsdUXnSUskjwzkugPV6xDs1qdFf3oWkchUtckoDsU6j7mlVrroSVUuL+r1Rv
0VX49tOkPBO5RUPtUSLwPK0yFEmVwGAWejZqKbSPRsloZkRd0o6ueQBWDSGfLui/
xe6YUG1pAoqvhBhH8wwQucdpzffZbONn69ELFeL+tqLs7bxdC1URHl88bVZQol7e
KcXm87iREVXg6g1Vl5szL3JtoNx7nDo7aJVzgBYubHQ7f17o7kblsy9TPrBRoHU3
82dBEi0BAmF5SZMfhD7+DeRPkp3typKQ3C7mr/Y1kRPB1+9Fpj0NUTnU1w9PVT0o
75e0UigqWxu7VbNEJ1SAQPJRDty+Za/OEsgGd6PoSo028XPLGRhnJskL7YPgxE+b
e1SKBCwqYjTqEqmxaBrbRLfS54a9x8XcyFtUBvoaB9TSGVXfn3Z4Uc3GFOtKcGvN
j3nZgp4FIKhUA0OJBfXPayvcSLyA/OyBBG3FOEYVkgz7Dj8EbSMUwxktQwfpamJq
seV+JeEl/DgTqZeEcfusj/ZH0fw2NP7cnV2rdlzwyr06/a7yxGr9qKk+vH2yyJEL
iYJgNdwGzXiGAOwCSVtxyaEd7ORNkxZGTjXhXkLvMyqHajXEVfwOpLDu/VwzmyOk
0I7R60LaOlF+1M7sBr00Pq9HRmEgEsy471EgyTIRnT7Bbkfi0DcoL3d6Hk01bhkM
vVbpoc+oGCKSUZme5AawnWaS/pIrDC16nGZR2DMMkOxAvZ+aaRMrUciAzCqGTCfj
Cta4P6JcDhwx/wp2TiGfnlR6PRM4EJ+/h6+ze2rDDlZxFwRdoZE7Iv2I7WiFwCCp
ZJopQXFDqD/EYcyPPCE+rebyaxFmfBa8Hrc9FGOrxE6Boi4MWjECLoavRG8oFjVu
atGeWiEx7kLDwdzXQVjOKgfQUBuxKYhWqxCykEo+fzBqe/zpSeX0w7rduCzaYKxd
Z1NlaJMuJgjprwJHSTBFmM42/oEZnzVhVoE/e0sfb2Z8aMSP2x45RZ6th6c+BCWw
homIz/aQO4/w4xYE2Qz23nxVtmiLKrLjVU67IXW18VdyugSO9pv+TChGntoUrZXK
6+44UBhOXc3hRbFqwUgesYMpKo9AvMvRKFQLBQ4ykSqok48gvV+d70YTM+4+kHqL
IYgBu3UGvHbk7UCdAJi/RLHCGeEADyRItsL2AmU9Ihh5050TxfCLJg0hvmrGZTjp
UFo5R69Ooimsj+pmr7VoCpMM7ndeUQuKunEKLPWUfUUsu38eW/78mPyJDdjS0XmL
7tkRc5PNqdfEJgjbINhTQtHQnj/ww2PFQlLxuNmOiqLqMAK5VtLSzYu1NiBlGb9/
FerCchrScNLDOYyAqXxDMRtBK3IougCFKpVeTEAyIE9QdxHGQW6u28a6j/A9NwBC
Kif/BQHyNgDvsV1hVxkbEpukxxHyZgUgwiF27bePh8Pm1u/QnorlWy5aV7lyxETU
0WvKiYX9jEm4nQuKSEY+cbyPtBldIRzAFcMAZD9R10aDyS1/XfEmzcLMDMmVaMZw
ixurOFlOFNB/14X7xq9Wjm3QV1nzITpr5HgvJ9i0Rg/LaJ5dFLlSoUPDgwHyZbih
9IS3py1XFfKOHT0teJ3H66STP9zbBsBrxoUEroJAGh4aYJmeoP6fGMU/JYgEEFBr
Xj3uJgAlT8o65cUmKzERlSqtYU19yvbFoY5HEN7hbQbJSyJUFMvmLwAVaVIN6/g/
r3QmPpfX+r5DvzjzSQX/Ww7eZqGDpJ0BuSM44hIMmwPLanNLz1ulkZIT4uLeLA6K
wz3/rLbdAEHCsAEG9bbrUSjXIbxKcRxnPY01TLWcWpyUqKRgMihxHkgV86U3JD02
GIbuT7UKDdsUysijiodC+cvExGGKMxMXOxOe4NPEXmplhFWsmdEwBwz5k/qXuagu
RcE4F8/5iD9XA3maEgDqa8z7tv/vwDtGk1aQBks7OmSxkMRqHQcfnVFJ4jlImq7r
r7TH3HJj/0O0LfRhlIoWLqaYR8WTboyrZZK1igWoSMnu1jteoUPUrQR1N0HmJLBt
dCHeVFCu+VfUNuinxpS4Ou5rjV7dqN37NtZyDkdN6GAxWJAKKRqdiFDfwj7jvmj0
fbAX1b0KfIy4jr7fNNSukhQTjlwM4Qev5wBG6C6OM6TY6bCRNLNvRiz9Fu8NzcU2
1uzf6PjYQCUdOZDQa8ZBBSD+P8tZLX4cJO1ILTjrk2FEPVfaom/ldrZ52LMtXZAy
aZ40AxacvOfKxPk3FW8vWiL61T/qUT5Spfn3HOeeqWBQWTss2L9DaysveEw7solM
YNxB0MmvOgRFnU4pm5cPm0CjpB+UiA41SQqYDkPx6LLHzQUBu/b2mpprl6xJxMG1
RLWbYULlGtt+7BDLzDfwW5NPYAQ2PTwgmKqJTgRtM738URTa/s8WVGtZSueOjgse
mSKYngS/+JWn7mIMnnzx56R4yIkspELxLssXdzFcb5rIB153vuPZgkhAV2FM1Eth
ynSm/73pVVkZp7gRLmvY1kwNu1zDAvwofLvnGrDcASUaXV5eSlidcYwztlAqQgbu
GRsJF/BeA6TEWNTXKgXo1aPJbO/tyeb26yIpT97Ro9m5CG9J7ezW3A6JMP9DuNXJ
XgvoCuKHzZL/M7RPANEMlkJ0bNDx5YqaVUuYYAamGY2MueFL9ppYj4LqY8MHSfkE
LigN4P5rGMbNvVMcbYCdbHnc3F3OG5Zf3nvwjh9iLPUzwPH98CQo+OAMPabjHjGQ
LBNs3xfMwTnsg5tlx17riIDkrnuvcO+LkgHchNhiQPQJqp6uYdu4Docr0DTExHT1
hQqEFOn5ayPdeXvhbG4Lh5QDCDVfgL6+mvaT6xJJqTgVEd4HzIhWesKmYWxkC9h7
+iq+7euLzBkAaeDVP1zmzvd6ebA0LoPW5gWTqaS9ZO2hlORYhueNYuy+jkUFmIiq
MMf4hhpQO/MBXt1gvpM5dgCqjaIx2uqLKyzojBL5m+PWUXGwfZZijRXkkt4S0ZCN
wLfEy/mqe2NXZ9F55745fvu70tGl1xkguAA9NZI3bkF2wSspVBB35AVbzBCLSWrt
wqZ3ZjnLeameJa8Tmp2duxNHHAYrW538OAQMT/DZ6XgkhIt2WRH03pR1zmgunOZn
+wFjwCgFSL8rMou15sCfxZB3cVXk23IHRXrpHvjzs7nhvOoXy5jXDhI8+WaEdTaO
z2cf1dN+VbSBFXF4PB8jBh9oP/vtJB+I35V8XjHAKH36Oya4NrLdzvGzTF1Rzehg
3dYaYkpxJHIdSBtKw7m0wt+yr4LJsLvoMPJCo3B7WPwCB9pRc7weI0+T0D33TGVu
OiumkfZyVuVFQCwy2D1TXCBSHTQglwJjBsNKEiKgZJxckyJpapLZDqgUrYSjqAgv
iCuSBf9uPLg0ESYurrfyHTCGm6hDYSpgizkd/T2hZ2xLio7h6gteoNbbwJZggSPB
MjNd3bJyGNWJfLp99qoN9IDHAidxppbRm8sfAUrSrF+Ua7/SGOJ/nszohUYAV34w
QINBJemh83Ezcm+1y7kMxTRZ2kYbEedWbK9C1Sqk847+ruSl7HHDe3QmKtQn0G6y
ZvxrIINj5GB1P8VBCAMNJrdQ34yYzmoo8Esq5bZW2VprVIip8pVXQmh6K9ajPAEP
FCm9EpiS4Ij24S+7Yj5jDDx8o6t+2cHKkeGdFHmB5R+xLb/4ArZyMTttmG8Ou6MY
kPNTsixjbUYGRWiegZE6zIxiKx9CCdjS6Vob25VTOCvf4+NQZQ2WQwKidVYDbSpY
RUjUvndVLS2B7L+iexLtoXTsrSfobe7nu8cTPrJHybiRSy4FF/9tYEwgvaMw8rp3
3s1z5jD6N2YPQmezOo/lrt6tPH4YBUQahN4x+xWjW3onNHiMpYGTXMW4aeROXdU7
ViIfiZDXzsl4TLmtrpMhGxvFIglPf1hfcC9RO6s0arc+oXO98vbj5XGlN4KiSoCN
XjXen7stlUCnnsqBiqj6efJP2sVoP6ZP/Ag2JFGptNcv0Cy8/sRnSL7Wqi3yWQLy
HuF9nGHymDMFKWiyh81xQPu0km1IotJiYIF4ZEXIMhxzpwmPAJHZ+JP9W29efk0q
tOrLi8IrXSBXz30u1vz8CPM3NETsoXwbDNzcy9TPoAdglJzurrmPyKRbAfhbl0RA
rBHPAEOI22FH1qwl8i7NPeCVbUFqkVCMuHXiYgdrYSHmbP/3Y0QraNQPR5011dKF
XngHJGHvApS1r7I+/UVOvR3kxQCQN1hGh3KMK0eAYE2SpfkQlK7mFTiY0gyE+VFz
hKh+/xAsdOR+Q1sNZI7EFsPaigxWHLAmp8qPHaNgNhLpDjpNO27ItWOpBehhl64h
iRpzs6rkzRTk38rWf5h+lQ85RC6UKq5WFhPxywrnQSwNjo9BZzb1cYpBRaIUraUl
ptmtG55/Hasly1ygY7jozJ3G4jsG7ew/D15YrW1u0sQuLAnB15Uo5HLITQJg3+EI
KHHS5wBshZ/6Geg4YsVX9KETv65vWhZeN2p2gKTFwioA3wxtqd4HWHP/T+a0H82x
uMPIRHO6n2X7e7LpFoTylVO52CELl9CrZEZIWesHhSsqTXlPhXvSVvHnkmh9kiJh
TAzotSHxiG83TrcR8wpEjdq8/wR61wgvJdRFd9I2Lk7LhMowcwKYaQ3m+dAhowxG
Amls6Hk/Tjpge2rYYI2ox+q1zmyRi7pTN1AqK+wfqMLAEYCOkShqq3scP7+q6RzZ
cnZYo3FTQ1Eoye/GY4fDZ0iisX2ccgy0V189EcooflhbtjNIzFhc+e/vgwbRhAeK
AOOOEAnRBdhRVsAKwVp+L1edW541wyORHSMMQ3exoE3RKrLfuOS9WC/VPTzUOh4H
oR0qkln3ei5ha/JYDydiwFto3tOSglbs3tnrZEnXuOS4X3gWXenKMW4hRe8MXIAa
9V2qhMZBdw5j9Dveuwg8XygToygCDMhGZm1jByp6I54+J0UbEGVowpEKCMJm6gFD
A3gHO0lGcoVy16A2J6a9sRFHNVuEXcTe9XDCL8xX2A/kVUNuDtukU1kFJO1UNLUe
UnmvAuTTqaAYAiYrkikaKejLzWdRxq8s1q1rRwfU9AQNAfSiNmXjrwPev8rlyyx/
gXcggG2+e8EtEQUpRxrQZVoyGf5hRUygM6cok4Q55+2e+thiBqHiqrYS+pAhWpd5
eKTjsXRirOerlNYfqBgt3zcLQWntYgfMZFTYgXwzlWy3yVxhEjZGJrJv1UGMO2L9
+E7UP8b1cUT91/Fgd3D+YIa4l8KAPpKxa3n9kngk2DxyB3/XsbR97kIgxcSC46ql
OlmLU0X9OCEs2fIuAtA4B1DoHuEu9EVVIf+qSqMD0STssysLZkqgNYZ1gizrV1Kx
coL0DxLslgNIQhhs4HkYNYwcD+CtjmI+EMo///U87/q5CtcafOOhNJ/+QT420ghZ
3DFHDuntGAT9SIIQ7VQ2ZJc4GHyA9oHnTM4286l7nCOHHf5hhuj4p0R0JdPDjr8h
fwCqNJMQfi4nNs3Bq+sKA3eifOlS55rNwT/gFvwzPJTDeMazD+DqzJKpJxU+B5Js
9HgOxrdMks9uTFAowj0KqOtAa4rgSphSBF/nurCCaD+5Dalwd3Ykv80jnBtQyoW5
1P3/3d0B7Islo95+IDSIdhuDVg8JdkvbC9fEuPGQvrC52pUF5ie1Sdx2/0/QvNUk
B/rAPgHB97C5B58INESMeSbtuwMgELpfKYJiMsoEf9CgeMThBSbXq6oatUJ+AMFs
BOwCpNoZdmOymAZzJXc+zCheb4LrHdS2GQbbmM+k4W2RYr32g0YzFgzXMeaNMuni
ImKuK62/MwLLhFsVEX4C7jEHb9KKPAUtWVuUnzjYSZU8UXCeAUvGUJ0OIqw07+vi
WKcuInhNMTnouQtTTONwdUaR+H07yygHSA9c0p7HGJ0Qri5l80UPIDoutuXF+sHO
rqXeY64g7VUsQvExNt27ARJgtU2oA6OmoWLQVT7xRNMXj8/PsSKd3iC+FIQ0yTZH
cukjdU7aYwQPXhHNZOlShEwC3J09NpAYrgRPkz/43lGkT40kb7GyzJ4XC4yhp7n1
95p4yRC0MBhKeFub4MPBdL5rzNq8+tOkwV3s3iEVqsCGYP7o1ajSRikSBykhybLj
ruttUuXRTRfyNqtdUjM+/UQVSbneyj86txJSfZQLTqRx84dQP0p30UKMIFgxvMfy
WIkLz5IZJ25MCAQb1zykBlxy/WOy0zcyRLQnJ2aOhrGOogS3XoaZDLeomK5yIgRO
kPvZMdTiTdPnUT2GeivcSjFxA7QCOzsuNwqaF1bTsD6DpUazlzq5UzmKHwszsVyw
mUe3ZR4WHVHONJ1IV1g1KEqCp+MmweXlGKfzbVXRQmoc+aOTiw7ZX9kyPObKDmS4
dMfGw5Bc+y14eJO+QqvIHqNjYxomlSrLeYog8VPi6fUtJ/m6CYmXLeVL1mVL5f+l
Vx1A+1IKIQntuj14E4TnivPueQHGCbAqD3tQZaWM/AXtuA26RY7vEo6wChJq0cAR
gsJxYNV8WAw5UsPJ1Zlj43xlyjDNQk7v0y2Z652zIxBhIF/DyteI5BLvrTytUzTJ
/ie1M8UlaIlhK+LHWwMhVCeveoslaFInbfXMOUOkQd6dbhttA49vqtfCFgJ1edgk
vZBB3dnN++/xrqLReagfW5kmAY8ptdQB2LIWlpPOVfI5PmHJ9ZR/p70TAi0ZHlyS
KFgTFJ+0BJn7YjEe4uEmbsnmxEscwhAJois5sAddfYLhQlNZ38ivPeL7KH0BHE0v
6i7phwEzRIZh92BTLNqj/afcSPTNatdEGlX2RKZ/xxKaizWW3nEVp7saxZozK6V7
CdCJp/+GyYFTfzabBO9WCzhjdpSWF+2krMFQBiYZ+RwGrUT2zLEi3membUB8LNMV
68NYc3WjwLD/RUEZ1Z45PDAnP5ou54/SvLjNuord2Coz13B5DJYLTXEAKYNLMQSH
ZyHHVqS15FKvykp/yUzdf85ylM9cppGfV8Vzi0KaJ3J/xqSDItnaZ99fA1NTxzjk
kVE+0f2DHqHAtibUUL4HmFvm74dmw5cHOhD1ojkZVzd5Uyt4kunSnSKPzAVwq70c
wTOAG+TFiBYFkDEFikqLO0JE6aZQUwI2CJzAujV45j/j3e6qdYohWXOWEXh0mVm/
1OFgbrUVAlicdZ/zGOsS1L2Q08HmmiAIBk7xgM3x6/0lxB+3yTggEUGfo/bBbtJ5
LWeT95JHpDPi7IwbJZCmyJiAF7YHYGqPDREoRzPoRcMlx/729qRw6fdrPOCyv9vw
gnkIXrfGChWKzsPchX2AB1ldZpPpw3Bh1oXQEPZhOKEgNWZk/A/TV+NSj2yYJAeQ
DrL6ngY7HTJhLexFJozYnBxpezbgkgDgOhZ3XGhBYAe3irCZN0QckJng/czHVKls
nt2AUW2kzlcns9lgLhl4/3ENSCLRFS0/FYM3TNAZ/YZCJWu8tVb2tyx0sCeLvYID
KWESBbOQu+2wYJ2fXvV5/PjKj6A4k3ElM8ro1il3CF9vm4JHPS4ttw02KLXeKbiX
O/wXBlMuPgHi/WqyALparBsy7NSrBYfbSTM+4qot+METWluRo6qwrCBUoGPgt57V
AvKbhcnNXYSCzwJdnE9TtqRL9qEWLG/bKR1uznh7s73++XKEEF76Q/TsdbX8uSFf
FwehD2x9VRFmj8lgw71CXll2TUdvqIfoDcHg1yvHlgK1zqecZZTKWJeG63ZYt5CH
JKQ+ChaJF1jV0COWM7aeHYRq+jpS0LGsYtP2yYf5/B5TG3Z8X1vPUo8shfRaOr0a
jE6wCfMKTgyrpwThWvO5rNPBmamvyGeaQSmYamzGKhAXjEKH8lum8ZwKt5rei/tC
tq+wqCuWMvm65BpGjykdm5Lk7ns13BnFMrLG/Pk1kSSsAkuKxl6w2pEXZcNjndR4
KQOcqgJdgwTdkXwcOkm4r7RXyv6IjTv5EA42rWoETTo3d345LyQNXo2XicwLq3Ki
bH6trPv2h+nfPAmKrkgg03x6iomRy3kvmu0b2gQI6qA4VDW3JbeDE5MTcanQaDzw
7cABBkBzHdo7tKKXo3TZe+WGh8wkwQNh+oBaHsYYWEQ2CmSvd7NuZD6TX9Y6Lz1F
K6e8ryM0wVaUx/gf9hu0IDTUFSueyNSBogqWHff3bEVXu3kjlMtEPbPhXAuenKrC
qt2L5W3akKxCr4UKg7Qb1POvi1N6cR+X5Vn8SqnPHYe1KMi8kUK05JStlePkceS0
6+KFNACWhJM+EUjfYNgO0CdVsDW7UfgkXMNlracR2hS3UpA+iIU0RooxXIUpozgS
axGqvTVg2CWX5SWeqBtvU/hqiR2mnU+/hr6pFrggYX4J+Yk7apSiJ6aVNIXrLjjO
CZ6w5v9t73lXAGmRIHxx+P7U3qTLPQJkqL5dR96zEKcaOkq+Vn8AFX0/O7gRau/0
L00lmwWeny3527RuuXvBVfI1JxejMvSZcyKz0ywHu6AlpwcvrJnanyWu7H0K/ztv
2Y1AL7AZocxkQ3jmTBAIW2MllUIhe7Lf4jmGQJxIW5U9M23QYovVHSdk4oePCCNo
FIbf59x7iGJJjn6BAViD8QpXDtESXvjPM/2KfkrdstrgmiKBcbCAYiSMc8TSu0mp
+hJiRyhLgHpbw+HwmnAqoC80SrP66YgIwf+l8vdH1QUKV69EYIstMnGF0wTtj+U4
LrhD353xBabTNoPuDUwEMcunKO7LOn5SxifmaF2vx3fmxPqZFR/j7Whf/e5/LXWS
FHBjxovaqv1Ejtd4uQzQgc3EIF2YmjWXKsEqwYTEEBbsXf2aivXMkdjrWFvwHAHC
e1w5+NSyXDDNh6lUDdycDfQ7F06+DHeL0DnTfkNfGrZVie3dwdmIWLNEEwU92LNN
O7eAl6FVo2pbrNZ/f5i+Gad2CelhRWH4Jj+qI36kDivN0gzBhdZfgi9VUcbtWzn7
rGZ5Pe3IvIX/DCgceZgXwAcWXvQRkHLpUVX53VbCBczE+2JT5f2U627aMoZrQkLo
tyVoxz1z3WnoDHabg3csufYccpJ97Hp0thhZhhEcjRgPsC58MRKAvPHqW8g+tco6
9OCNXwczgyaZuY/GGM+R41II5tR3QGyZOdWVNJrJhk7SG50rWwuiWlsllMr80TAi
4TLZyXROXJZhep7l/JYhB7nf+AoEys/9jMkSqwtUSk81XBThwfcZq2oJEwezLoJl
IkpHDNJhCTAocrsjExFQtkKw7NyrYlJJcgW2FbnlRX6mzsqg6OfW3B6P5BT3daWu
UgwY25BBN47GPOWaD1opxuwBwDjOySTrENeWJqSp8WEEQs/j6TFY5GWvUaWznw3e
CsobEsa+wbxGbzb36XVTp+Z0oRgLYGEQwJjjsjDuWp4V08Tb6YEcQCUryYP0RwDG
FOm6Uf/vL4+lXotGs68UBzyiODXIG9Mry0IRjNLAofanQcBghZYVmSozVIjQOrHA
WduQy0461p13WYaL+SIRV3cWeiHNr3kKV0Ii/qUxdhrClESq7jvOOrQw7bB/eRMd
4YbhGIgG3T91LGnLX5WasnEfyzViTPsbyC5M92FBkoL8OtHbnIw0gGHxUzOVXExK
d6ESNdErpwO1I6D+gsc0SoaeyJ1uKuboeDkazRfBqt8oRj1BwC3PBN9knpoNFZvd
kgLFGROzQCpipFQ/415NHGxf6nNS8sXtYHHD4tyuQRCC6ELyuLbf3igxKqtIZbV1
ReI9A+8E1kr8Kz1F1OwnnRH0SGRIqDm+hZl6uUe7TubrbMSivdUdLQIzgElsl0bL
QsCzGHdAGI+2OCgP4PyFhIRfzLWQUhsuEECg1tYdvgVc8SaUn7YZlQLackypDkD2
kVH9S49pS4YeR29Dhjf0WiuOc7SyCjnt1o4TQDw6SKWwBTE1v66pJVfJxHDrJtsj
IrGy1XBgfLGaw0sL6lq2PgegieMOVpN6Le9YUMmazCx4yeiuX0pB8DO8FCbycyDQ
oZWYUaahZh0H8Dj1WbwfnPiG2Bl/prvsS2A0SzMbzIxzirPScnYHzX7vgQK6bRR7
4ZfC36WYOH4//kMGQfitWKwudsxfOeeRh2xIY2MICZKk5eGIeNshl5cmCO26ECcN
zZ4Pi9VwZsg9TgoOjuty8YJozr2N4hkX4te+9NUfvhMobHVrgFMPY2ykd8uPVvMg
Rap+aYp5+bTHGbOkoacCQF8mRo+g6znUjtj9AxLCIS2JiV8ZftYzx9pkBcu6XcRe
3mN6xxDrRtVRkEndU7O0QQV8xR/XgptZ08bTBRHa+5dk8ChItnDSpWVGn52DxyLg
n036hVFD+2B+yuywWrFmAxVC7Hbxtjy7lo7QHJD562r1IUMcZFx79ju3E1fr0wlR
4af6PiI5yFuHviiJYznNqRb3lNGFksZc8rM7vfIz2MAD6hvx6eq2ZRENU7DjnKle
XI2LF0/dOne2SdgCp9jszSWYnBCgaqhqxkTew8L8z7sVJ80fHeykcakGM4dsQmwE
bOCZYbfREt/Kv0xDZ3yNvME2EJVHM12mYPMkpCNF+ghykrcQA5jk3cwWfvq67/TK
pVJJiGMVGs6b2IqT/L6mMSAF+Cb8qqOWz+UZSjr0AAAdy8DFlaREqYwBGUyuJyji
NHWl2Ai9H2VLxrAW+DelU22IcNyirpZdsF6rEm8vHnNHgQCg6SToWu5ugNnYLk8R
/+SLGvYGYLl5WIYE1l2P+Y+0w1PgyKcdCyfsjnZZ717JbvDMtGpJLmNRbpNEtwOF
K4KZauVF5KLsZKCZPRieY3Z2vkyv2A3OPmgFPBfpQhn4mVIX34E6js5JnjIfFhYZ
jBf1xDloMlq2Yo+r25tF+J8lVCxWe0e4td/6Tz81dhCbozBWu1H6+odnFFWoLo5l
glgS6E4qZ5UOWB8eTznGK0YG3Gt0e9UvNBQaVnTIVbJG95Y7COpEfjC6ZfsBCx74
9oesivLdO21cnnGgr0j4j8oFpAztRJrDGcr+G8KVLJqLpPZe9LAFssVRWCr12rq+
9xc/FzjMGZH2uGwu6mYYkHtZXVHFQA/kVO9ZIo4nlt3amosIDWtF3S1s82XzNeIE
GaHa1SqOz5Ksc5EC976hCWh8cvWpTIkml3KjoK/bcogrq8lfRu1fGy9kS3j4Lq3m
30WlsmmrYOExmSUnzpP2IlO4L1PRNLG3dbP0SclzjjV3iJ63eeo6CHH+ODYjbo0w
yxPjWNKZV5TDokeHLa2sx0jHX007IBovKBlbfww9jYY6f2D5BuPbSh6f3aixjNcO
twNC33dMpRHSJA83t/KG/qDFanbqH6m2tAx53vZG3kfP5ipUCZPtvd8dAOGbJRq+
39qcjRxbm80Ifmx+ODIRlsNCyDx4gvqg9+cLYfEuY2a7IYxcoiSIGfv8CLz2Qstx
pmmJ0aCcnCh2pAXhdLSWOvXGfQ3FbKgDbeXG5f20qSvOGC2lLzDjusrHyTMDxT3h
XreduC0qtBKXNExTi8d22CiUTmw6yvGqFmXgVLhojxXL4ZRdU9GVfLvV5vxYQyor
J9dBgqfs71nEg1GPyJKwvnoc/j+lTMDR4LzLpeRfnNCx1fsjw5v9GbytpZvfSDn2
xuipcLxlRP9Jd7KJBBpzwgUFi1tTRRYqUU4liLeqTpi5VTse97q97hqlM0iZnhPj
PJMBaVMiFZaG/mhrpuh7Mbp5muCaQmJOlHDWQpcgpacKHsY6UIJVU62X6BaNOoRK
lnFpXLGcBCG42cD7JR4xcYaRQSi9eykNVuD6XWCD5eU4YArnArcSgEOFCa5dhE3y
HKRNFeogcTi2tlwd2fSNhs3DtwSSI75HYZgwWGx54iNlx4571r2BbCvbFnJMK2n9
iLwlMlDtnwGQxWu8Hjcw3hfN1uzJHTsbCePrGxcjY1Rid9cJWPFleEuSJc3UK7q3
3ZRVMAgmBmjzQhYNUHC4Pp5HBbC5F8U/8hWIqpPF26Jyf0I3JyeIVS2L/5SGKYjV
m65GSpMwa3sR3avj2FkfVoiLweM5WvF8d8bkOWgdt5157o4ec6aotdCOfIzd14w8
kDFwlNQlyJ3JM/m+BWAm/IQ/ciZuHM8cynmU55ULj2QlmKKlrrZ9YP/NIGnZGGzw
LLZoZz5TNn4Z+P5Q563P3ZPe3SJ+spnQnxXMCX0rgP9iYACojGOoMi9ftHPifO6U
mARtljyFY5noGQla4pVRcm9ajBYWd6uvI1vRGmrEKIkTHD9sLhaubBSQ4Jyz6S5I
mrMzrNyn6RXhkSmdBRZ3qk48YQdz4Mn5xQbXAtMeOW/sk+TuGtTFvzgC2vpDpGKS
2ckOD9hGE9VwLZcYbXk0I9Wu0qQVJ58i37tkuPVuAHv6oVlKFHO4Hs9Dy6U8BmJw
j+3c5Pm8ngAEDvnEVjx0//8DNrE+TFdKwxNMuuQpiwWtp7nNLaa0XiCpUAgvHeHt
yVtYvbQ3chlyfX8w5WpfsFHOqJ9tzNSKgFv0wbUk/KK6cZKj1+ifsLTkRF8qkVb/
9dB/nbAYrtsyEyOIxm43jIipj/1ifQiPJ7wfMOzpnTv9I7rwwHEeBTQzRape2dT7
Np2oMzPefbmTCn2ZkAjvXVA51He9lf19N1bwt2AbBEh96fUPMlT0gSSA6KntqxYr
8Pe/aUiJzdP1KRVxXf4CZYnWk39sDQKRGtnv1BUCZtFwSg7xXgCe0/24zE82QtyX
a9bJX2Z1MKw8ABcwzkHfoYCPHQQfFuLVIxmSaI80TiQK8I+tgFoIqsC3lghN61xD
Bdc6cu6j/v8a03TyAeGjeUZDC++DAMWCErQuLLT38ebXPKf3vlcb17Ev4aVPyiLC
rOU97ixPy2OlSY0z3ItnKclZ5MV2yETU0fdcwXap6zlY6xgVD7SyjEZnEv6q3rCI
L4u81qNE1VSaUApJXQ35fBiPM7TpAuw54kZNjJsyskvw/SEONds4uy+HzgxjU9DN
VknJ/4zmS4TH32IyegwU7UfshLFs8UYQDosrW5mg2W9gUbJukgBS9NglSl25fk9N
/sPCxsn3QvhtTBdkmQHdymtND8rUc1hQFv0CBnBxKewJBekH+9pH6rzFKocwIHUm
R3r/J+G0b78xXX/wXkhjjvRrSjQ4a163iIPHVPdDAyyC1RpouSxtaXPXrzqhWsIO
yg1LNC0d8imwu59uSggdDgTPY8aoJMYCGnno9Ia6NSNnbM1nCF7/W7whqG5mutCi
2V8UGeo6JMRwnHA7gAEWvOW3YZDReaahXaT7IqZVHO6FA+NjxCFdgfGgddI1hbQs
L1FJvP//bQ3o5dMP8GSsjfr1Eb0WwxZAmwzDs9hCJB8RuQEK1NirjojUGmwrU9GG
W4I/e5u7BL5ffUShy+mqn07IViz2W4a7d3HGN07Evuv8XP1e0NDQW2hELEMuT8hc
CKUjBlOiZeQ9vRkOthtZDv9gOkAAbpbbSCEwPZNfBSQJE6ogUO9VH2tPREaQ6gR3
wIpXhB4mwp/5Qal2b+26Jyob4hKuuyGxU1lxkoX5MKqVlpe3VNSm0pN9lWKk8Jax
0ug2AJF6lgyMNhsEeDvENWTW/84icBr3t+vmQID7xW5YUYXnQakBlzPodlcsZGKE
YsKhOAxsuqm8kKRQs1aCuUtzbhHBvz7QY+puNY/jMLMpDPrN7wipEUX9TfRqYz0Q
LSvcAtWW3HlX6sIIwMLd5rAk94CbJD117m4rGOTDzmyXNkKDOQ5K64cFSxk2m52q
sm9V5FX9hpjxGg9VJjcUb1eJTMJXnHdtyVgGtD2KaIX0E17t3nAJ8RD0TkDiDEXW
J4VQZwkJvk6CvJlUj32XLGQZepDZe6nAJe6cGtDuJ0xBNtvpLX0y6EcjXyaidqYR
3lv0ylVHeILo+CiEAKgBhElTDq5LmW4QkEw4B64Oq/FXAN+ZzGz5FZ6sifdZqZqX
P28kFbwOZ3RM03yc0k2IQMfyNU0Ktr0+n+FKHQK7DJVAeThLq31w+4NFNeSVf6Ep
E76UXXHh2sG/RqcXQBnlEJIftqTeUmGCCltFn2lq01JdBIie+hZqkCtSLMfN41zq
7WadGPMthjUPHXF8yNanOVjc8QFK6nalVo+Mu91uumOtxd9fCbjr201oTgoI2ma8
pL9pPvSmb6+XSVda5VYwtS75VIF9zGSxCpGzbqvE0h3QwmunCoquq+N8VK1TmPOC
bv9u4rQjCiMF2mJDIlAddDEdB0sh6QobyNN+aWg0sOvFsbGt4wwFQnVAo/tEViNP
+lYvbC+uwK2e7pWn/NX4Qruh9JQvg41IFaVti5jNYixZ6ajQR1UZVx3E59e3BqqQ
wwmgfNxu/x2TfLMUZ4D2dHDUCuldoIcqDXIO53KFUejP1uT61r+caP3bG9Lp8s0o
YAvBqlgGrwgc/R3fkTw0fDfPy2iDJglb4YXg1xBRKAHqL2qe/dgL6tErPctRaS+p
sOBjrNux1QEctnsrMacQhi1sR9YLv3HtkW1yufZBfis/b3yDUr1uDIJdfMJqkk5Q
3NgHzmHX1InVAu1wxE1lgw38060JkniDks92/vJdCkdQPOS4NLsn9NbkQ745qGXy
yGwYKVFZsaIQh1mTUpHsbhy658hq7qf/O7fC6dXfx5o37PKbJceqdVOH17vIakDF
x3eStpAadskLEEivLzISJJvkODU0118W6eo8S5DZW8D7L+tTPhLKQmFiftRkgHfE
3RHx2hiztma5ZsccGLcZhC49dbpfy6qdxb4haJUTs8r2Px9no9ibY71V4b0Ldgxb
fuIwZBrdFxAk6m2r4LHUhsZJu1vWUlbYMKOxYNDJtx26654o/0zqkuPOv5Bh1BOM
eq+DueupNPOhudXlL1Qw4jTOPD7drY5xbYpLuhi00EUd6ov1SX8rDt/lVLxMu553
T4qa7FEpvkHYLANtUl1jxhV4Ic+shPLBgBklDjMsuHyjB2zcs+GnmsAOyFWSoi6b
4ALv3Lx5hpsKDDNlTp0tFs8ww3EWoyAXlH9d5dwQNP5fy11mAd00J6A1xODzk6mP
2OVNi0oCOJ/0Ptw6yVFU7AOmie92kIyR+8Pm65N8fS1vGYvnRgf4WFSz4tMDfEkh
cYcQd7lvrRGGabAfkBamtxT686xBmEkG4XYDJ9qhQj/NxblBKrqlmWNWnRi3M8fm
H7LC03bUC6aRSDQN0ZZ3kU6/dtX6Qj8/N/oRvWTQxWF28maGq4KgEYMuIawCu98C
A541l6KUIqdt4Qbjm1vI0Mu9R0R8FM5pL+ijPUUYBJTqGuh13iMgM5INY3H/EAJl
n24IIX9TQcQYhpQ6Fi1pKs+xSnGUES/Dya0UoJJvkdNlqiS0bbLT5ULUOhB/DeRc
pW5h3QIInERIoH0/eWSWeALgaoVfLiKKP5ZfaIEa/wZT3X1+GRhaXHDTl8khMtUl
AiqCowNOLrfmNNMwg26e2r4x/vdAyVWCtW5cAI32GaVXivKkADpo/V+NEchlxG8c
oSeJTGCrmis1OZOr07rrLmh9vQChXGmvBZ2vnw5rFizDFVtdjRivYVg5dLjTRIFs
UhLVcM1WQa5t6bCIw/PE3kCJvQK+Uopp87Bia6znSJOHNWqehSueGhdlC+l7K8cY
J/1N7C/0nO9V4BSGz+wG+ruKylYjwIaBPVXEOuVWSPaLEtKKXhRJrhjss3jPXT1H
nmwQXT8xWqs/nLcURFN7//ZQbYEQw5jgnn9teiMAY/p35VayYPVvYUHbpfmDwPQ2
NWSRZBnualBScoEEcPlo2H+7eW1eVKmTx1fxvzCzryTYmfplz9Pr1NwgdahrJNK9
ZfaawpBfqKzcldJrAtHfyZIPg1KD96upFFltb+4uYZdyvgHoLo04GadpU1t7cigp
FvUqhjIW+2ne0TMVZE2KJpzr7LosliuKVQu4ywScajU5vtX6/1a4dNSR735q7w7j
R2wrFVR+54PYJ1zISIl7w3NUyeif/NwBn68Gc9WDPB+qObrJ5QrOaBvH8SNl2UJF
cqN2qIOmBDbnQlfkDxzU1Y+PVZLOyq7M/+6UW5baIOXK38QjTd4OuybR0Ms7eOIt
jgfnQUxBHzsfgd/5+EvO9VOJJ9NvcigpQVoQ4osDIFnWATwaMzR1Au3Yk7McwDnD
ByNTVK4DF5KIbhR2Z+nPwJa+BHN8tKvWppyGdsaHd56xKjZ571Nhm+pmHeF7vC7h
MOj1yuyZIcKkgYK4Jozq51Bfo0HAgAzXAaxs3PEiKom3ZT07PJTBuYEFdNN07hQ7
nb+ttpd1SkAeQJSX+lLiu9W9iXrbyFpTtzlxT7Ihhy6ajulzHB8xs1h9Iiyc4MT7
VrHcuuQV5m6Lk8ugTe2l1nN+1Im+XZ56MBQ330kKUi/SPqQ0N3pzWXqlccR+ovPM
oaEas2KBrgdzoTjngb7NCWnzqjuyfntlzMAjtvF0rgTVPiZ1XdSF6FME0w4X+1dh
KbnOSh9JjKKiXd1Wb/B1ObH0SKr1y3wGvQnj1L6BvanKVrxa0JZPTK4Zp80iu2y1
ESu8mQcaeScGbyzXMksAke2Jm3A9mAm3Bdi1Mk3KdIg5xPZrbuYfFJBHiSBnm0+U
q243C/OBLpptBjJBkFzJTUKj2Dvr+cRVdk+2edS4eY/aSNC8P6ptR75W/DWFjQVQ
BRSPbJ5eR+wQy+tqHFywdI+U/fzyu1V2UFl3scdlQNq+brvyf8Xz/3n35uoZKLF2
zNMxRl7PZaDM/si/E/uZAYdkeCIc0BDn+sdvpBj5fXBv0wqfgWFOo4OKvBFdAhki
hC44xda+/pm+Kky+5tEL8JXPdHl1Ox4xES75oQsKURyiyCjWRWfovo6YRLTPBpbx
qU2nlaTbAXEVlffgpJXPBfKt4y7/SLZktT7FWOy0V9ZCl4Ys6NwdQ+16Y88I+ri2
5cTvPHbnjeoFsXJVbbuMcbh+cVk5oZDg9MPTzZp5Fb/1fpViSM4W4Tl0ESHIUT69
UmqlBw9wVYhJRZpRdOavN20PV2kbe1oirlWEpw1PJAdFlTDYd+LqBlIzJn3cj2qr
16wdUYqLOa+cSm5oJ9tOOk+cW/9Dgz41t0VDuPP3Y/bzdhR6+u4+TNCFvAhKfIDi
gB02xtSrGHKmcYbKey7MdGVgY+htim9OmgQP5kE4euRgamY7aDf9SI3EKaSXavEI
+/W/PIGZ6RadiLIijNk8C/ITVJsLf/eVW7jHc0IsjTvQq+21XX6IyQnt6MBKQ8ln
+Qo6Q5FYTe9SVnHucuPofJxPr0ri+iRQ7eIl15IBi1oUZuq3EuaXFc3AU8/nLxV3
Q0PsLBwrUCTn02qtVIvI7Ny4aAWY9D65HB3rCa8mg+aV2ZXJqKfuu2yQ/fXDrkgk
nm80/JgagkR8WT+Lq+bckg7yc1NAdsEmuiZDZtES/mAnf6NtRrkhEWMQKVOAtv/6
GlmnjpcRIZLQs4E7AJu7qo4TO0WsKkeQny5lRq9f+Vh6EeWNUr7pdTLaKgJ00nH6
CYcZSsds4b+Zg5ds6kABSpXoIRxbm8yIf2XRV85dWN+gYhIj26b47T7HjnZUfRtT
oulgS8fMePclaz/h6dSP5JmTFTydXrWSe4V5B7KZ5qnACVwsUZW+ywtenUJ679oS
V0hb8L4BubVhsQ2MbIqhehafzbcOlfBHRnwbMrJzxC+DoDBzUsNlOyF6ykQ33On1
2y3CYqCdO4/gHVAWs6dLDWk0uTt6QsPGQ2itnzj9e3qwMnpYIiSQkFEmSRpBSdR1
a7tWOfMV1rWsqNuM1G0wFd9ZROybPd1oXGfbKA63egTmZRRjozFwVbSe5WsNfAnw
pXXKXo67KeCyRVEg0klksXz/3/Ubx/V3hKvcpielnxCtHioLNAkzXYmFWOjPFa6K
83jl8I4C/mip45t7L7tYCj/AurFE2rMafDN75MlJgRty0TcGwwZyzucyBcFR3y9X
qqTF+THIKBRZleWEKlrVPSH8gKUk/Wnxu3s/5c4NCaF++1sUd+bNj5XMa0e1ZnNo
b2xC9Wqo/BHJVWzHP9rwhxPsxlL0FcN8sSAdrZ1+gTfU5piBT2RGQyAjupowkumq
xYQK39MEo6KrzaFYEOOL58sGCu23KTPCPfmFGXgpwY84+R1sI6jNEUsNgNACTuxO
uOFC7B8RfsVYCDaS7LGZ2Z6eyj9dllCkIw7iSrTK6gOIx2GrbTrLAJxpoFoNum3U
uylgz1SLizXH0oNWUUQN4hIgF1tX+2ITKuWxl76tcaKisH7VUU/gTMaJxwp8NHLx
WF960mI7dPQel5pRJDWEaehi8TtCJBhLlClqDfCIZVYG838ozznYUhX5rZLPYMLP
exZAIugQWM+0+OZ8EDuh3fyeaoNVEYvzqEMgVLqD612NpIpoIKOeEH2COCAyetXk
QN120xlGzL5gR6ad0NvgHRwZ0mR023DSoIwshw0a/1Iw6GLEH2QxZ+2gnJlTZFry
/E/mF3TnY/ZQqiPOkhFTreREeTc0Em1HmETMEOjyd8wBb+IGNN+NCFC3PhE9e17+
+8T7TCOkI53MMHISEVl8KJDSZjhn6yV5H36TH5+LgRPlP5TQckbBjoP1MFM7JV5a
FpNZZpP8P5lg4Ge3Wjw2Bz8Xu516IOzz3g70YOlseXUvmUUbVLhlTAikOFmZsViR
iFBm6f4zfF+jsQNt0O/8Q5ytMWqIir4rmxityBXI8V6Kd+tnBEPdbcL/qdDMM/QA
Ocz8kmdTXnDPbxH/rp/WQIzBqlTa0wm5FtryBMI8JWoUziMkDec8XTd1mtIUlu8j
MUssSRAzy0+IZ+1QrXgVzz5N2CLrTLwqFSX3lNAPeUqhJhaz1ZeWhgsKxyWeeFAd
9z8ZuHx5yFt2Ig1m//z2XylGHqGeE6TaGEkgbTYgfghxIDHekCUhrBAuwSRnnmVs
421eUElBfvyWnb6WdKZYvwmCtgo2L8q1d57q2LrKrZCdiD6YyMg3csWw+z57+AR/
YmyYXhF51Sr+sJQobDLU2IaqgZgF71/MxKC3uQSffuz69hqa7eKli4eMk1Bn4x8C
cMG9FyqGZrWa/mYo8mj9PULdn4FR/a65Hh6+4+L8+Yp6IeigrmJEMEtzD/6ipeQ/
vquCR9TUOl9ec9EfmQcdgvRYc6YQ90foxTO9f3guDkmMAlsUaILhUzg9IruLvqgH
GDsQIl2IwtiG3G21KzWzGLkFxDwMsYGfz6e22Xq/fOgmENTYGBn0jCWQsfjhZI/6
sQ/uRdvXMikeQn4dyCkNpCwhutAiOcniuHNI7M2oF8uo698HBCSsBhRO3NxAfxoJ
NmWO25VtlWcWj55b3GDLjMd1W4Ok5KbFDGp0BpS0dvH4JJx4k1W57BE7dY7Fs+H9
AhHzM4CdBPawenMxH/TS8W8qxtmTej7SSrq1oQrZNrSnPStsLZpdXeplEJZOY6ii
8Nmtcc20Y/Vzfx2i+LfK08qwUiBRd0Vv9+1DN2xPR8zx0dbxnSwS1bfCQzs4MDoA
kHkJstDcl9GWI/EUsTrmfJpdonA66CZyVXxaLkUjGx7R/O9PfspsUZjWWoUoH1HA
xWVUWt14zm6dErdVAUGxe1IOVNMOiZs4TBkS2ZCNmmUwy5lY4dn5gVdhEs02Xsu6
v9OlvoVKyfTLobAnmi2GpGCQVG1Gst1Lhk94veyxtvzqdWjrdoJYXpaJefnEqdyZ
VMTKtcKd+/hnDNiiPccEOK+9U+cEoVrjXPdlSku0lb3ZKMsxz4zGtf5TnqtSlqv+
pBqPXDrv/IC5Cl9c3/FM3s//QIMjq8jboMQ6770mtwKQsW4cWGEDRJzRJ50+uy/H
L3chyZhhNbnpm11zdNlydep89CjPG2RTzIagYSGBydLoJyKNNr2Y8MvYwEjj1If1
0T/d986W38KWOIBxJP9T12+pxbKsTtOrskQ5pvdKfroCSMRO94zv+0g8t7glUEYw
qZW0uyHvLu2AWko2c/6F5gQ+oVQyMUwE0XakZzRbY6FS+bNT3ftn6xwrDgUoo308
99CWdcl1bV8yzPB/bfB+a6UBj+OKBvmqGfGbCvhiC7XO2SmA3nrTib6vliPvSykK
jXVEyysn0JyFODvS3xL0FNfGjVOaG6ocq/4zSfSJWh5vtmXCSLN1ItI6iYSZAxrn
xTp/dHwHX4+d3Ay7vVN9AHAxmgJ8A12r/xT5+UCPamf1RZojcix659RyOQtPLV20
H3h7PCnCQuajvO18Gnl1pbuphOPtypR9hLfvfxj5zKnP2Q0KuUqioe8SXHSVFq+k
5kOQJ3YD1vkd4luzsRO+sXoSeMFOYR1FBqB0+pNpN3Lme3RM5Xbebh2xWgfzVLWH
YHKRUJN+3qKlgxciYrHLe6BY2klM0GDtbp8bbcaJcmQvYrgmszK0S11pk5LTvGHD
drh6YI+cys/LNA8iObfT1H+ba6ouSVYW0gdtyLGgeVvRfe4OWR9lSNOJYsujB6NH
xNmnbttXktAUpNawgeDlcJwaEBPT/fbaq5XCqckglEC3VBQ/ciMy6t96masrlmDs
MzUbf7QMnplZn/hyPGemkddtsdUxUv/UiCrI4JfkQolLkETYr+2k3hMzV4J/gHL0
m0kfI526uFL5Vr1tD2QW0BAM96IuY3qvTvWJCP6oGxg+MO46aE+S0skkepvGDDMS
wqKCaH/9lUzJE8JfrooOnKP+zu5v4gvES1b6HzVElufM+LWU0riW/bA5oMlw5L/c
CdoCkSo9EAKaA0E+kfW4WnS9pz7ex7NRupK0kZ8JHDNSpl2u2QMCuNatkqPFsXa4
xssl5YpZNYdm7tvzUqjd9w1jlQd5aHfoiTGyLmfGfBZE/tSfVbL5Zk24l0HcgOQs
4XlSNy8izfbQVKiBo1CHerbpv5kuo+954fsBnWr2mwjYMXd90ff6n7yqPsNKy1Ev
BYz5hJASmtLXQRl4D5tX5gbltdEJPWuEJY7Uig7nRmQLoYfYqlStksH3T3P11z/5
VL26VDrCkUzyTi1HeP9l8lPlA+niUg7WWHio8aZBe2IAppP0a35xMofJxIZSzUr4
kchODodUpZWYVt3U2u+UXCgOCWXeFh1DMFI6WCkO7IdpWaogiuYUhhG9LXvwI11o
Deqtw1skFIfVNIuTfUP5DY8paNgYyb1/RvhdAcZ8MojL0IY2l9JBN3s5PpqdSM92
kObZ3FEjsixir1a4Qp5vPcZfEoJfBxWjVWVd5kWP9bMQKJgGkRO8eWQJ7IyPdN7T
bpCbVHUwMwj0a6ZoFNJLr1xGs183mxJD/J5bA3P/s8CNF09OBY/aDx3IfEIDDSat
Qa5docTpBKGe8IcmocEZl3aUcqQKk7EgPpoAVxosH5TmavPO9SVYtwzWx86QsjQF
f4IvsIA7pBZwp7rSJWwyxIn1b3h/FzLe5hj7ukl4DYFXnuDP4rBmuubOSRMmXxcK
Qk10awklBHJuhQDNVgIL9oy4F/nzZeNp1HF4sbIbIaMn05leTG2DPInlkBVfePzs
y0pQ5TYlM6FFYIN8Jh4OStaVdmKAX4RMW3A/354jFW5BWs+tudf5loQ0oZA4ln6J
ODwprAprpcB3brBbzQbhn/v9ckat9CYZ5Bjw6JIZP79r2QbBDXVNpBqBYJlpbDbd
GnE/cN4TZuAfsSDx3HExcjvwlpD/l9drhhues+fRPTh5YNgICbW94MmSfybNgAtn
q3uxeMAeaxVRrEX+O3XEvDRGkyq+G2AElVP8IAAXvhCf0xD/wmMPsd9u/Y0ZO/US
VpsmbR9qEXnQLsPHPLx9rpm9iUY9U+9wy2uZC66sWDyNZ5qY9IEEgUQmg+Zo+SZO
NcbHAIHTIHrCrtk+Dr7+4601mhaarRXhxJfEZYVwpFnR+XvfHL39S0z/xw8K6JBI
MFHGHgbh4e1/pwf5qeHBCwfaMm3ETNOKV7DQJpq04aGfwwsrGEoBePCU68yzUqIf
NBgh2lpJn1cJEL5kuCIGhlrP/DTyruBHCPRGjeiViXOD8x6i2OdzyiTh5lvajGFj
8R05ykHZ8dlccx6/h6dHAbjid1gKGBMWGT/hHeynqqitoiazwCSVbwiYP172CgMf
4GR+BJBvWKJVxVcl3MqO20E9IO/2911kkUJXZMveSPVES5EQed0k7lxKVh/AH0Hu
vS6aprANTZJtMlEH2z3IvDItTODfFUTqEb9og8tyjOQ27hR+JE73evNJY6Aac3BE
E3GoBuP1ddolwAABDBY0MWYbBDl/KWqhGpKBV0pBTQ2mnpO1giBceRttx7mFsgnP
BZ6RxwkXzeLd/Yyp9UnU6+Sy1pWmfvhEg+YliNaCk6jsQd0TvlHKN1RGzR9IS5Na
QG6Nf/0IiFk4EN+KDWfgkYabdHIH+XUQrImYVHjdz4O7I+MNQHKtnXaxJoVINHPX
Jr2DK+0Q9wKwNBxobiO+wrNQCXH4jX6VI2Yq8Q40afDlzGoMuU4HYXkpAHQn165k
x5G5M2EkxwQpDj/LlvMh7JpWa9YCvea0yrirlnV73dJ5KYV6tQ7cdrpqo0P+TXYD
7L8hlctiIDNv3rrpXkPTELOdWebdrKgX/4TJWDYyOAuMwZh9AmvRFzPIv4+vDoy+
RJ/mPz/a/4U4girQIo15fHG49IBExEdUOxZbY4oPjwZlK5KGFgPH2eaxq7edNHmY
oeFoZQ6oJ+Jd5E1uRTcgdFOpV00wxBlDHNEEsdvYdnc8D5OivybuBvf8iy4VdMWE
ww6WjLEKx9HNSE6qfAIRA26XG3N1YtiJ4OLLJK80qYfw+KzsB4sefdzR8ACc0HhV
b9XJKl7u5If27VlDPzqrFAZX4jW07V6teMPidDna9jO12DBTGFoGE818+TGUKhCy
RNTrURRT0bMNlIY4lP/icccYoENJtppakJahiFHQbJuVhS/G/OxMI5LNDC3uvGJ/
6bdcctZ+f8KdhTncLbrWjGrCqJI9PKK/4cs02+cLGDWq0wtspKJi4D4S8b4k32BL
AxXVKNsECU5XqadFRQbpF8LqW/bpqP/5gsySx//945ZrsSj5ooFm3KuULFiufO+J
pJXvbXykJSepGcjxavfFTqyf/8S/cfIxrh6hQ3ByONUWd8e7C2CVYhXM8ijsYBGT
PB8DQBkny02CiapZnaL2WnYKv/agP/LLAFMcHPHBwFhVc1I9QJFe8XjmPuOGblRZ
P2UUyc6mhCTNBIfuwQlCMR3PGKHQC7pxSFl7PcF1nzWzCkgjqHD0UrkzGmJC89Am
sJCIanP1DJqshh/LAYu3nwItV6AwtwwLb9yd5RfMHjTFtCafHYTxaJW/TTVoTCJU
OgxP0WlRZBo9XV5MQeWvYH6Z6Bro5A5d1lR+q0VXe3kcp840V3l0MBEGM/9jsU9Z
wmQsES8LQXrTf6WWKpbkxN/5WcYpaQhTXJvWbWwI3dVC6aA1hjBHsZBcBAFy8u/S
zYWuLaZh80fw6fLhWHM1THgGL+NHOP/w98gqWaMccTv8dArN1MlNGxa0o8DtohkP
mUl4Zowm8U9sEl5laSwN//Wa+cy2tIGMhId8aPM1qGXnWJUbQ/oQUfWsD3P7rEu5
4cFSDKu4OQCNxpH5jfMQrOYbHtEEQq9AB9A32wM5pj4RYPARGLwHRSjQViIR5113
k5miw1TDJZlo1pQehMOdEige2aN7/zAJbQ4zHFTFQ5wmP0XzNs+8wVDSLCA/5zji
cfeGzqB7j/HVo/Tfr2+HCDHgLG8DQczQPRPDNZGhqil856yFWM7JNa4+qErhnGU7
tWRCoaactseHmz190NJ/9dbYHaqvwG+Uj+hpMBBkOrGWFRxW3A6APm4G+Kh/c0qx
mcjL5NC7zrCdx+jKQ8dgws8WI+kDB8Cr36AQ/t5M20610edIk/SVIIq4AqS4AQuD
j4MHomiBXHwJALkawishayx2+sbFcxnTsH/8NqfxluRTOYLszT8cZwFRuwYgX0JJ
PleDByg3quurYyojq6rkWe6hg4N51c5skyePwyCrKvT0lE3rnEcnziqsZ/DEnIww
WvvMpQlTGdczyPXmv35SbWyIZJ2QrX5Xt0pGH1j1HFQhREYQeohTUBvGqarM8rVO
tMl/1HoPCit2iaiJd5/OvifVH6lvofQLN4tUqyjn/nCNvjW1UsRHFKXpXX18giA1
nXNz3hGc7r2FzHAbSHDxCubJP6z5/73NKKuXu7Dd8ShAVAC9I9hWOxvTx6rdWw6O
3ji50Dfs1u+5h1BII58ZKNRuJcr2QphZlcA+KH0/vAy14K+Cp+7lvUnn1WjrSz3S
WsdngvJC1TJDWmXhVWhJClBcvHdzWzhaWjYZmxvv3TAoqSq4lYIytxEWlxBkL6p/
mJ2ig0hvXS8UAD7X/FhdyOSPzsSXyNg0vn4MEzWVMfF7+BH4h9qKwawKSn9uvxgK
yB3YX7kzfspU0NFraDDxIT29lkA6swjdxobTQ3AfZNkfB4peZp18Bvw55ghvpi5l
14tMJ9Q0EdEBGa7RsCc/9v2nMsTOk2drHYMAr72fO4GybHlhf0//5Gj+zVKwxJAg
g+DjcfK4CYiBh2W1fnOe4uPLDCWZqczkYol6ODyk7ywYQjbQ5UR47otLJ7BdHUv5
GBRxHu1yX4/0nJm09Wg3exJmOnnsuGrnKbtQO7Fvxul+Oyu341XcurLavgc+1yIK
Jxc11w0SD/OewlD9b/LMNI9F9W8zpiGBJAnz3AkepVr7OlDqck59AypGMjhy69A/
NGga12IXYaCgzDZ4EpL2FRkxbJwnHFOIXM6UmsN0cjeh+eP8dRmNBZwJG0KDeoS8
pJVqsdbwpURM9sjcSB8LEcUgRY9Q46NRCUoFd0QYYHT6Ry84By/AyZ95lC5VOXww
QrLkKhX5pCwY3zn4Mn85MjfymNobcGcVm2AGkzyFJQmh8lUF9I1hXH9BgmqKg+aC
LsNdVL06iiKHrIyiqHhzNlJwmUWNqRDMMVBr08IuuO2ii3/ewzE6hYh0byoLUgru
cky48q6RVV6DncFBdVIX8AS2v8d0wFyAeew7X6NzDPTa6AeI0OkVja3D87Gnp3pi
T8yqBbaWOOUt+ArjNlRIvUDE2xYWaSpzR351zDBeF4JQZJTCKzUeG4S6tNcqakQg
VyCykSkVt5yW7gN7iT2n4S3kxx2uvETuPYIM+odpSvp5jzApdb5cdYeJoGXPE6b+
9of8NQ6w9y1Rx7Hn/sSV7gZ/jOuLZ8yLZtuIlXaO/BBWNKqwobzx19x27FQjy4Kt
I/msSW9LfbUhRMIBSBfTJY1M3xBo4GcKu14SJ4yK6DGekVnWOHa6A7/ERW5MUhCC
KRL1c7eLUD0m/ljVFc1LOec4P2WX7xRmlSlwd8J7gKoPv0KPukjWyFA0uB6i0Gr3
a/Bd7i2j5Z8Fcj+rz+x45eCs8u/omRaP2dDUWMM02IpD5kWbHoolYuFssKE3gbrt
mwZ6zc6FuWjJTi/p2uRN8vl2qVtEtjoJuDdyJ0nMmkALcPJo2s5lCOFw3fijydTn
tl97x6aeAkxngOl7PIZv1rrzYGZaz/e5nGGOWN6tkLhtHImI9lfc7aGJzkVtcsee
bOmt6wqQrvjR32DqNwMvujauA7UnQZWMA6XpfLABkzln9tEeg2MYzR862/RfycyX
1CAW7qUbW2DI94OZ7KlOBJzQgGwoN3ym61UW6gF/oo95qIpnhNOLXVcAnDX6y/LQ
VY3jX+WCEF3pPDzGtM65us1H0zsZlcGEj2U+dGcL43i9IQXGlPEtwwhp2Of2ZrM1
+SQkbzlCLyi4/wfl7eQm4hd8hGH5cKkzBmR2LenMynvHcoQ3/fzBghooJSvxFYXy
2/3Fd0dVoANxlN/QIArzhZyunZ+gqxKMyI9CvvNCDsGVKIEo91W7a2Hbv9aJYg5R
IYJnntgXDZ3txDoM5udYctbiiDDH2d/nU58FMbWE6u3wAkVDe8IQVVPdvEJdHUNH
eBVNhrxMQyLw1b+gXyCc3RCgP0MprD4H7Ki3eoJA2VyGOWAF3dCYNzLZZHXHJ89a
ICKc74Ww1JIBhscXdSSWPvuYZX7GiTf4OwvZm9wdHuOpmnUq9C1aSeXSUidpQNsE
lrPw5ynkFcwuKWPRTlL8Pe6uHcEsXrJGyGq44liQTIrL4JN/rhUvGkRvaclmsO4y
2H9YLjCyXMdbsrsurXmxMpAUikj0oMAhUg7a5LJj7s5dfZQ4Z009HCU8BmZg/Jrt
ssmY1peBwqIZQmr+MOfxqyTFGv4j/55LR1SKbLdqkvwcB6X/KecJHq/LSr8C8Lqy
rTdHsuC90YaSAUv2BudIuM8DEhKvW8bdakQQvg0VdrvKRgizr34owYf/T8BBYpxk
yPlmk6d1JqOBtouQXJKFwSao52SyQtUV00eQjZDG1etsE884zjEw5/FRqJ1s/KQ7
EbsAHJLo7pVAVD9pkfzzPKu/UVlUVdrtlAreAD8ujR/vidc4HgLa31dUCAvP5vsM
/HB+PaIscFkIopnglCtG2lxf0joWnRBT3NLegypJVFLWJ6h/cVEqdpeoJs+9tAPj
hvv5C3FMpgjZgWMoYUbBNPhJh6tn6OuiYovycgKKfpJgqpYSPNGn7IgfC1gnfSWj
vEZEg904MoFtJVinOC/ukh243S/Kq8LExEd2k7YNYh1s/RGninkRwpQddbHUmbcQ
PDooxfQ7/VHrAIm7Z8VGStfeElVsqVtSZ1x1fEENX/oi7PcmwfXaPl0NQPCrXqmx
AVy1xb7JijV+o8XQ5c9+ckjena+EC3XPwYNb/SiCe+6/1XDJ0IH+n+O3X37R06Is
7ZgTJ7PBuYHew0wNd71XHvoAqZbf+3Wm9gv9HBE83XkoJQXZ9p4xiB6na/9jVvVZ
qktiKi3Uj2/N+MKiyL2eN3tZzv4NyDr/+zODZzvLQQDVP3fjN74pvum6quBvTQDq
PJ7I7eeLOij7TqF2k9+aM36nTn9GtH2tvAVloyaHLZ2o6HivmywlnKCYng3ew5Kg
FsEg3BCIJXD6mdcBqrDB3SkZLBfRDGEgeN6jhcrqdmijkraDtVtB3APXerUP8nsH
AcsGBnP5BPIVKM6/eNXQ2Aesj433AeqLkTifQSZAZ5VLGmZD0FRuP6ZlU4gSLQ2T
5J6y3G9XomAOgg76TNNMkeQF7mB62300xHPH+72YyZ2EooHJXn6E/fRTPLH8GhWl
gHokGcFo17gifMLsybISTU2T/lJFOcp00Ce68embFMy3RG2JX/MLR7ug+1ufprSy
N17OueqIXYQZSKLQtXDXU4J/xYLSUKWuT/Sz+Mn5A0QcRfzFXfnfL5Hqj9C0Xd2N
nRAPkTC41wkycYbH+GVz4HJ3Ve1BT/SmID2X7dEXnG9MwtzpOM09/FgXkC3sJPRM
Dqzk964Odq4BKBd0G6PiArBUHMcPhm0f/6BQ886hxGtATkqrLBfk9APfDaoBXAl6
JjsBRQHmFXDrH9x3V1Drcnv32L+C4/pwyGYpXSkTqMDnG5Xf4SzVLJW0tN1EU8K0
E9vJgjFOm49OVQ0gmes6336b36vhL7bSe3y2oyYzaqgIQ7EhsTDekpAlSX4vuHG7
O1PNxxKmo+M9HZ5rbi2Hw37CxzyT3tkAaeiktKFny4awgM1J2Lr7LtERkbnTNb/p
u6/ElHrCgHOBKVBzQIpHnUvnh9LkQYnM/s/nWDQZKC0V8q0dWc6SHm0RFa67haX+
oaM9vZYP3uYBOlSGa+quC5psyRUZ07fTfPwR8auol9qg1PuEWTNrY7iBTPO4kjJe
imYfL/R3ZPLnLpvqYILo9lZscebQdKgNUS6cmqwVGzUx6f5CohFF/f41boQCaBWh
womr8kfTbEUxJfcd9wL9naVtFo9QmuDjTzDwviU4gy0G1+awneozBj4DiHHlnHfx
q4DHydLGhJex3nHfHtuimh4w+d7RvBu/eghsnqJAGB+B2gJf7UBSyYks8XrfT/NY
pu9yy7lEU9vggOfr//UthvtKRhJmCLNBk8F1qr6tcObF6Fcdvq1h7XBsWScpr/r8
Vps9KX2Ly/dESW9KPYFWTe97qKwoAS/2HQlqS7Rh9/e9+Vjhhv75ZjkOVzw5OFIr
cIHoNt41zYJxe/N5/hO83sE+euzx3cRwKsaoT0XLWeC7ZbJpX0d8Dxvzj1hwfkji
GISELIPUm+yuaiKYvBc/fnpYfNqPhRqqT19ScXSot629p2aYm0jpLOLULV5rJjBP
Qds0+lRiMRVF2/MparvKWoDbmnfRwFfSYTSCiQ9SaPap/cJf+dJIlO700OBOr0jS
QxZ5SGBfN76Y7RR7q23UJsQ1dKUS/b9d6jxZAz0JojcMWtYpyT9Wu7D6NMJRxLYn
c9JcLqohnYImhPepbER7Us2qERqDc7fTeakiZKx2cUBN9VFILC+6+6oY2sIscZW1
htlKsS7KY14YNadfY8ZfDfStF/bZful0LvUwmIF6IxBdLBskIacFmlX9JlEmyFbV
NKCDTcTj/CYzr1lsTBDinCvKWzB3x0VPJ/YUJqAoBjVdIqFtqyPxQN7tGWfHhb4x
LEjesVC8xLtqiB5ThxzZQEBRdQLzmr6yiD7F8rgQfQHeKlxshFUH0+e2Evj95aTP
D5ykflut6nztmm46bAsyWk9DuN4HG4HPDyIT1CG2979r45T4ShwDsLCL9UiE0utj
+2/Pg8N6e40TWDrTkJDS739X1frGWLjns3njp2nGnrsAz3bavtNAFPxXm6yZO29A
DHg0BSUYTlmFTqVQqBDQfmj6k5pLjYmmt1ybqeVxU3xwYLKbc7FijRfXQxGhKW9x
glbjJ8WHoyyqgQwB5okJXGxiF/hu3hrTt+iU7mt1rx9XhOICJopk34n/z9dKzH5g
bRcJ2FkRnjLTDUriBmZQJCqc+n3YqQaujjxFl9ajQom8KjJOP03Vf1e358urwQTw
DuxmaKAa4edFDcKCJjacK9KAg68L4l+NfvApZ/MjR5xBBzlIbV/8EaLwnrbLo+eA
VTRJjrpGf1h5nnZGhgoPuSIwW9tD6wQ+3//kTNGLuoimcf5BViMQ0tGykaA9c34a
qo9x+hJOS/+BgTk4Nu+fROopvVtb10v8K88/J9c0hmX7BY2OQt55WPomNLLkJvLi
qSTT2OlyIyBP3kf82Z1KwU7KoanRuJmwFEBvspfmw9qlyYsQOpjbv4Kz/g8ZDXVL
BeivtIB7odFGuhTUnAIo8rjDI24PJYQqfJX8jTce4/sKTF+Pf1ufVgIb5f4sVzev
yx6iXWPHxuCRN0hLWG+2/ZS/U3MRzjFSVOPiFG859n7F9smpfJy4+k/XinSg8uek
v2Ldr2sAuUNOTVHLjxzuVQ1NbXUnfI4M61kAgOLVC8PDBQZW41GmqltCYyDDcNYM
cdvV91rVqIDJj2gH0c2Rz0P3hQz9pcYDKaDZvgqNGHeJYwl6TbJcBc9ui7oct3sg
DcMU1QcUqoE8sTAvRyFTpTO5tZgRc9zyGjYM/NGsVReAB2OW7q2ZtdkY5WnNYVbw
o1qx0qEHiHb4Von/mJMTdhIVLB69kr0mQwJAT+yiidy88caZ1kw7UQN+q/ePeWMV
dzfD6+fBNqWSUntKBAfiMkWYq0mlENjkhHlrydr28Ixx4tU3u8B7SFfwNqyt/FOm
wiH5fmmlRlqjl8Hwkfo1jLKLBjFTvb+PT/op/NauXZHuMHfybQifRM3DRMLh3DNl
VhK5OGILHd9pmnZZneullv7eL9Ioo1UD9Unr16N2fHJDIYha90XdfI0LJN84ZObM
SOzfJveY5F9LZh1bjwN45qJw+KI0OwUExtp7fGWP7tSaRAKg1E1nJQ++zDVK37Pu
dPyBVjQpowwoRaE1aGAXtGZ4rRuDdHsGjzGdsnJD1xlzbOIIUWyVfsGGlMjFuQCK
hwQ+axaNCb5hIpS2Vh5RZeaR1Q4pBK5izlc9UwQWVfA+5ZnVYfnW/o7+fnEOi/QP
WMMAcYpVD6uvzqg9nRkq+64Z/jUb9fpqEKsxIjq8gbLh98HeTjmQjbG3PEGRouaG
CNbnAMS4gE8e6pFqvq2smkKYV4QY7IWoXQihdPHxGIRWoIqcqDrcnbyzF9mIRTmS
RB4/9lzY3IPsFkFSu572elt49WWpW7CuXSM9HakhcBkZkPaIk3y6uvtBr6FkSlYI
xem2ZGUQdlPcH1mWYeNOI/WuYnQqGpzPzV67YXoSnMBaqnF58ypBcMR3BVZRtukN
WQ4QXdnnI+TLSdQHCvcZsBNu97XvDNZUk7cgR1wokVAWUhR8QfKPsXGWLxHcpTGA
HwJOITYo3Kf+TRT1pLjLyZcx1kBKuhrGGwdGL2ublG73xLJp+wGhfuXYEU6uHBOn
2U+Z6BQmcsdUFaQAQXt9V8XRQEmhNaTPvVlwLQg7+2fXbObeX2Kx2qPsHnOZkxaZ
2kuSBlB01n9WMH9rQoYw3flKhegq8uYYrsf8qnVoumTEh1Iu9x44iYPksk3RZEhV
aPFJ/CQDNbr1mDfAomUbQiRNv8NHR2FTfXMAMwpDg3v/ugiB65YEsH8zfpIODhrq
jVv8eeRgxpsfmJq81Hbu0/JnM0jM2Rn+nWYaeFnTX801ks6vdq7495O5aVqEeqZt
eKeN3OFPSC+4IzussvCpZ6A2CC/fsHuqD0r52uHN+/Sk0zHEsug5dOWpAkv9VyXl
a1jmS49FVAxLw4A0hS28ty3oyzpjl76GQ5a5V0van/R/Nen98RDBsoDENHUzqKWk
C8Xx9dH5xPSths3P0kVtBSzlytBhOI4ct/3YB4Zt+rXSakKVldKbthsf5Z/9zjy2
LxdF9CYtJ6kaFy9LfJ17fX9DT3pjmxsPWcRJ+onSSOYcElL7Ntx93pakve5zA+hC
d2o0bpWS/+OiVQX/TzTjpwjYGvtnHCVKPtPH9QSUWSz4+DKghCys75nw0V+4xpHv
Ok4m4Yq53GuFKhYIrUMdgF4tJiw/BY9c6/V15STgG8RCYFKJl3pBhoUQ53AwL+o1
tm1AtuQQd4eLu2ntA+blsW2QgyXaWHCHkCVBX3oUzNIg51qzUMMjfAYKuI6VEryf
9HafLCLU3uCuZ+iPWaL6rihD/Xlqir5VEbwukTDqC7MiKUNWgqL+LN6IG8AvcbSN
l9FgeZ3SDsLD1FdaVkDJWf1oXrzefukXRiA45mLvx3H1PHYIajh47cW5gmeRdr6e
wOCcA9j7glOEF1wBk/9DttmQ8BOAXwh3asS7mEFBF4riQf3Bu8p3IkLgQUlbdD0+
CuI6Urav/KSSJxgOc8IiS+hZDzTU2OLdUzNRaWUV0YGsrdqDgZucGk6X5QFARHkU
ZIdadS16JgqJ+HlMI+S49jl6bzfMfLJyeuDA4Ms2/l5207tEnxWZ68M7xVE6109u
ipViqWhof5/UU4i0Rjsb9DixcDiDMJBzDUBIEStWrXpijFro47QLHh93hZQxazTS
hpWYPXfjqzSURvmCEGboeL2SL2eOsSJIlSwqA3xZ9yyYnQ9K8ypiTsvGUWnODw+w
JQmdoJ1FYsBfM7H8PGd4kaQYyZVDjiunMgXAC3yMYMSut3gW4pO04quEvEG9/4Hi
9SB7d0G7T3hL5GCmnh7h+tQh+VCZJPGcIpRqA1GUyrtYwtw9giJbFyN7pvv0v40A
qmzWiwgD7enl3ykKETde99NnzNke+Jzn3EtWi7GpdxLkzr1ReZClQNL8G48wx0lI
xJs0iZxAAATBo/hA1c6QN+YJAUvk366t1phsuEimTW9+BZCULvTd0xZNiktmV5cu
VdadRXPgL+uJnh1LdcGcP5hdaX13UtzpVV8RChq9J/Mk19mh6XiScPAykqRBuu+7
Sp1QdXhYlsBkrs0ELQMQXzm73c94rXAVheuBD8kINAG0yVfaauIemfp46hLgR7jE
kShpTiEYMzCXVD5dO8IeAb6iV2WAmLyODgPkbrgHyds3zFKLMg01u2r4UwfMUYsd
j6yhUdqHWQaUMpiFJGGI8vVUOpNNfHJCb0uZZAGNgzHSy83Fq0lBPLJ2pyoO2JSf
Dr9xYO2d51GSBEIb6XpRbfGwHFXQGyeV5VNw5jErVegsH9rxs5EYbBcyhPnPlDQ5
AVLh2rQR3xkceDdqPc/1AfYvSGi34WfoBpu+qT/TfEOonmjEAQoCfce1qkTHEPCJ
yg5I8NHv+BPBh3Re7Q47KcImrgpSIptBGECgAsNej4dfJBnevbBjqZ5u8XqqH+vY
/BYnjBFbr0OfL118ifRGYklSgpapoR7EsKwVJPg3vYxOJ7IupjqayWNk9Lhl+Csr
Oan7TUkP8aDtWVXvOkiTfNvwSxXLi6dgH+DiBnC+2Pn04zaCC+CqbkCCCjE0kU/W
u6OuAZ6pgMU9OLxYQlTuYSYZUeweMZ0Fydhe32m65rc8ilGIR9f8ZZh0Il3G0I1S
ezxPLXAqS+hB7rZjcRLfEnZQz//+Bcb35Indl9wspxdd6IHSDkeEwpA6q16AU7Dz
jg+gKp+IM8tbnz52r0fSlZ9jk/pVLE9ZwKB1kVA2leWUgp6hHaL2lUJckeeWXuRl
klVTepn9eYkyHoPUtCvSiYL/wsvMGvGWlbMI/Jkjk3XLVKePA7rOqxtuZvF6VBqO
R45fxBd7kMEu3HwmVb3f+ck/audxfDhZSMBth6uj0hbklLsMOl+x2vetfzfdUos7
NGm2FX2PekuoTZjbbReYv+RIFqevbeTzIgcAUJ0J4ze2izEAfDBZ/3DiBB94RHqs
JJYGPBQmPl0OqlLUlNZWn9Bd3ZKGX+cWgo9SCpEP4ZLhchstsVD4Kskhu/J25T/e
Wqpf8v/tt11A2PHwBmqGO4IAQCfeAquDXok5L8gGrGbQXNKt7+zWEc2Ymw6uXJRf
SI5y7ufJ/bNO4RtImaYb567bWhqjojmMlEfXWvgNSrqxjXghtECq/gijlNvef/8M
VYDMygGoxGbsRYiem6D2fJXvoYZeUneQJLuJtbCcrQ6uDBtsf0SczvbRoijAjxLr
GRSnqYq1cYP4lZkuPEauSGjb6/5/ArEge6NYLvwFvVtrN/p1N+JKDvjmAWTSFvKy
zN7QIFOS92lg1BHC1863SOb+S42JpUpQF/oJf6yuvvlfynWt99GhrdeZD9g3PYox
T+1DoDgQWltdLcxcYw15GCYMPJBu+y+4/3RDeQ8jpHAZHKEAha01VufG8f5B5reg
PsAiPsqPXWcVhOUHCLFljlq/FqNsdomQ3kTnwu2XujyY0K8e8mVezwUR/m2x1Yv4
GbosgQY4X7GToNh/w7kcwoQeziBqdEGYasm2xqMwKPGx0zlytt2/qMhwt95/gV95
DvkjbP2hew2NoEOTHSNDRXG8IOKOpUU4DD8VwPEhSjooNrVJI/5d9qAQCrkSB7Tc
/2YfsNf9T1gTQZfm2tLFGFj5FisFKxSJUDnEURWVbKEbGhjigrnIP98Kob6atL6r
BPAuYHupXvfLd6GZpWUycOA560bsRPpp6aFZTtXYGsmwGIsWuESkeOkoACzul00I
Tzm3z9jFhVa5v/tfn8A30HbGa5sWo//CTr4Qn3SlKWGMVaPL2MpR4i6e3phuyyD5
EsTv4aHzPZdz4rCj/rU1xtID8hQJqUxSU8LaOvClKqF0l1nMrFLKcGkH1h5X4l7r
Q4ihq6QTJshPKIg6OrDRVKQLGZIpbSwGviIPCLFA+EA7EFrUvQpq8nE2DHC+yedn
aZByqX7Li7axeXICnQO19FF9yLgdU0WPOCTMBiJTm1t+xGhm9RPeYh4ersI+CNrI
P6atTl0KorBlY7JyRA+Bu0dmm0ymHOsY43zAFzsKQ4a/iyKrMBRFZI8/btSoe9ox
sNi0I4cwlncCHtdGKyqlGHcbJXPKIMZhQCK7MrLwoQbTA6mXpD6d3NbMNtWkF5up
yLKzNygywvBDTNZJlP5EpJTTD2e/cBQpc7eNqXaPGMHnct1t/GQ2Mga6EkaGNIIe
Xf9eCl5TA0nMmVfxwnMzfNOtPrwbUXmxVUd4t8amLAZNyY1Ep8fqdpVpiX9PMH8l
iMlylzxL5BGGcuL46lsLzLT6ZXMaBi2YplikJxZ+jgeX8NCP3f7vU2LIWGPlmsL0
crf6LA3pmMNTRVIAUmFAZ1miqX1QjeXGwlYSVV/1qAdc46OjMWppAfz1CeofwjbI
MY9sQuZShLiHU0sfmKLY/pRHb6rM6ryKju7wsjJTSd5yhfPCi9uDVQesxXNOje9b
JI2Z42V/uTgQghNc5VAwi6+NngcUXE7ESpd5j84OX56p+mwPTeMgJa6NRpabw2gW
hxr1nmHht53V3oz/+QOAK3k5Iq4+bTARVCjNbeU5BYBFAm4X59iljbzXhIRwTa4s
7zRphIeyo5Ambnq2vIKorMoX0jDqzSLT0NC2tZwtV+KgkqLOSQ2UkKCKbWT03xWf
lmPJ7Pq/f8X8vamc6HKIMxMkEQM1HRkpSPyBKv+9Tk/1RGrg1E4A+5Z/xhjRkKEV
tAGmz3wtuwtLc512sfTCTSQO8Xy9rD1DVgEiGA9cu52yNNjVH5/HCG1iZaBgiFgx
MTihNJOzqFOir+84Py5tq7x4TApxhQecYunlilFzn/zJwCc+ZrTTAHwOvvRGfpPu
YB1JjNYNjYN6Pnfktzs7dHRcWE+vG3C+WuHBV+HMRslCfAfPygivoVg5ZYGKGDZN
UU//d68FuKibboyzOiJazpnisjEXzECW9t3b8F6KBid0OZBuedcnAJtR2NUCcxx/
HhtfreEwVsHTFIUWoyXrfPg5yobGgVE2/KOtGq05hcdlKQZ1/AndA7cHFmpoSqGy
zEWPOxGmNskC33OOd5+JFyoCDZ9dFgcgqRKJf9wcFHTN8+OBBr1hbzeftkqcQW6T
od40MC9rdhdIouv/HXw6KgNjb55CkZMo0IT6U4Y7xh7OoE5CcQ6FGyHyGPvPLAH5
qbIU0VFn/NvaNPiNPvZ79C0i2KzzZadbfs38KMqFrcXv9toS/1qsvQsiBI0af5zQ
JcJ1qx8yZ4zy9BTX5pCtD7E+k97wIdXn9/7umoMjSzJJpuC7U207w9R1tbaC46t3
+HoIv7Ipnwe70FdC1NY40MLLpcwmJLjcqlCJRok+mVLXzCpGCeRzZFvrbPmS1npY
tiE31YOh441gNiEnnYPA5UW/2UWAlO7AIJ2CvKFGa5geM+qEQoUQshnww+5vd2kz
npAlh6K8Pw9OYQZMmetQaKyh0lyAU/3DL9zJBNahYa9nsDU1/2GBZ4yxDsDcbQqd
sBb7M1+MEmR/RlywHO5AIHaL72/5sPMYcIu/1EJrWRKbnxjUtv3E74Cx06iW2+FQ
PHCZt342L3+UslJJqdbjBGTVtF2ChFsThVX4Sidc2VExgLW+t/5OG2Ecwd1Toy+P
D9jTFw1ddLBS8mQ38VSFJDFPigVP6tIHroFDnbgVQJn6ExB67dF0vljwIIH87mVU
msPk5m9lOmA6AuPMpP93cyfl5PRPzDlWxVFkjW6iCt0KCh9XOifU4XS+JGZagD9/
TXS9sbNZeIaDifYTENOxlrb2oEYgYxmzrwzgn3J6b4I0LtOReJD0I0yIG+6VGckx
3vRhxjtNt4yGd59R6ZIWSxCnn/oVCd2mkTtHva5p0cGYQuGbFg/dDUHxdz4YBUVw
+SLnk9zjZnJMhN+d5ahDbE07zjRtCamuZMhNbStWWIipTYI0uGwDERCaRlWVZbny
FhGHlvP+3PTKK/Y9IElXlQ7Ay6/MEos8wTKd6jUKDHN54JodemHMIS0PpZJ1EePe
UWoz4dVEqGb/vS4QfJ0dsV1AHhPqzxgsE/rkS/VXMJDQnB3b3dthWGd7sxV+1+kO
4HP783Gtjaf2YilFdo+xI0zOnOPPAgZ05OAIZ7y6A0tiWdzG08IuWgb9VTlxd71U
92srN+4rhi77HiXBzlhUAma3Gj3BRk7gJ3DRVomNPUOCutyveH6aazp374T4OWUM
tieyNzldIUinksWY0hdBLN6TT6y1XdEsIx3rg+AtKRAvLrpkaMntgbCJ7gC8QaxZ
+OfYENBT9BV/bq/NsJ3DrHi/NsDq6BpcCl/BirJUao3KPilJTLfjCl2paBbBzku1
wxXSJ8pK5W3FCnEmjL+yI2+e/2/tnzfTd3YDHNlqKQ/i9SNHhBMpJPnB+6gLG16Q
GqA9VuXr3OQ/llE8hahlBFWkv8LOkaDk9gY6lgMVZWwe2QhiTJu4JcM2nxK5UFSY
2i1URZhF/f7oQy1v4NqOrJr9fGtFvXh0d0a67HDqbI/vJMTDoYL0WphSn7YMtaGl
FYiAWYqRfPz5x9nNjnDv+au2WDNu+Vt71WDhIu7AR7beNBjeFTeTqpHwwDnfpIF6
Fbnh0JXQZaptu5cZPOUldLSdhAg0GXUvqJFTaHMBzRj+eMR/Vd5CpAxQcXPYbb4Z
pAwvI1p+xWORigpTuE87yU2MJoMf9sLchbbmqWsYuSw47U6Ixi2qmUTfzeSMG9Fy
yT4x9AqL3TrvRMinuvUY0625kKG9JXFac2uBVdiLFBZjm7DmOIxdiUXe1409Pm8b
phFwRxtOdHToKL2RAptEFByFU1CN5tf2EzOUGuP5jwt7nI0XNIcpj9SiVQxiHA/3
agYGKy3xToxofkJ4Ph7uNXezrMa/cdzgml78SUVNBKUwpAtONgbr3dzgK/1AAS8T
3a4DtiXG632XDwtYLZWjEsOjz3Teif43SwoZjvvL6pPrd7sbMEGLiPTXYOr8MFdX
BZrhWNnipw9MaifjeWWbJ6f+TVmKolwyn15hz/mUPIBvF0vvQG4GRmtc/RTkIBGU
Z5j+raa6xdYuwkvSRSIS8pYJzmjAqpepjnzv7Q+2dcHqG9OAlJlxfchU2bi9yS2c
fx0ywi/CCw5PsJ+3dG8FRMsS2lee35ucaCpkT8qgoTxP5QeBnxKiVQIJ/ZdG6GUS
My1mJSKB8vX5FcVvqQJKr8EUXdFovbFTCJXZro+ewZ66Isg2EjutU0QGVdHy8Xyr
MMO8OT8hDaFDPrfv5ajU23kUUQmnemWwgK8fz2/WOhR83sol2cMyQwRyqiH+aA+6
lOi5+Wh3XQX1J0wS0S67iVOsl5m4c9UbUf5+pMrAesqYwce63PnYNZg6iYWa9Vch
rw0CXKp5ViEoRTPFeZ6/ZKH5ic5/8yyK5zBMPoSJLj8I9MIEsmrIqRYTEixqkyLn
TtaN1L4gc+ZhgT5Y4yj1ugCjr3t0rdahzAvVuhdK6b+SJKIWTOHFyFy3trpSKwqu
T7dnQd6eFAzCHuiMImssaEoRl1j0e82hOm+HsbE3OtL4vtFcZBLrUMbfnyKaim9E
1wmXhvP5kiwO9apEO1CVKLa5xhpRdiv+BD+Bb2qwFawPjg8jqFB+DxHlOAtksinQ
pkmR/yxBYFypEsnnqkzxKWVk9jooeyMKGdAoGHQo2IyHwMsybPRvUj4MlO9FaDTt
H4+1T7NNIDW0dcxRcWgJr5BmgWq4QdyqtdtOkVTkxnPPBOpQNgICvwM9x3of/tTj
0QQ8/SrHqRh/9cH2xaMca/Vwr0ZVxiyKbM8XnjstvkMdbWaIlQ40iz9fun87tGJQ
VyhP8zWC4XNSikn/wEMaItv3RT7mpZ0HFDLo74twaMtYU4QWjE3ptICmJ9jt97aY
Omo5q1DbwNxgI9mn2+jhIjRQ8Od3GcGUa0XTT4jq8x5vuPzts1as6c1Lsv5Ze6MC
/snIa2LVYc2VXWuwUGTH3ocEEgOHnMpTF2dEgv/32GC3Ya6zq8fm20VcEY5Vf8Zp
+zmu3OmgK1uF2+SOOIcjCZAt4E3WodXi9gurwGdrFCUuvidKPK/CZ62uXQmsyVSa
4w3z+rvIfuAMJvGVF24zp5dJ7XYhUdh1lAixKsHB1t69HoBzXQPgcMc5xCcGWfnY
5H5T5Ovnlv/hpM9G3o1qfDB+URxad2jVW/Z/Nbn9YExvYjJwOai0jbwsTWL/JO3p
eB+1YrdGpQnkg1+xDDjOOfGYSgaeLZYHp+wxm42cI75ct0zwp/g5O64HGhb6z5JK
Q7pvE6sA5CBb/azh2IGWqjHyLMTWjoeucRyPBW9/UW+nNv9iBO56C4i/PDQ5dTvF
qZeVlXHysx1Qm7TpbPiELeyg8SWj7V6q09Wt9iUgJpyh7/dlcXzFK21ygVK/9C+K
Tbqjg+0RoyZepLLnTxuyCYWBrrxIKlt6YZHZUHZXnjHPKbZ2UQJmYbLXF/10vLoO
Hpwiel9EaKMJLZBGljSmbBTBfAHx5+Xoe00CNfSZDv28BQ5kUGu8Zi/yg07MEPH+
wMU1W3J+ImS3n6Nq5FHPOASdZwyhPE55KZ4znFDMueAW3GMB4D6UNv2x0yL5js63
YFU2QjstynTj+WaxREuKfnIir1GcRfcCCtmLjBSnPu8EpM5ixEM7u4Q+W4jgpYam
f1IrSoMyf25K929BDDfj5nhPOOfyZZRS3NE6UQtd9ncILllaiVJnYz8lZ+iWc2us
iam/FJk6XKYX5lkbD976BkMBHKini2KkWEEZV50bXNVJaNNz0MbfmW4C4HDA0b9T
ForPJOnp0zsy06WxiqEXTv0M4zZhuTUxZBIAzuzyedqTaygB7ogxCte5JBd81xDU
/IPG1c1XM1llZK/ujHPaz9SR1KQK4u+gT6uvAPAomE/iYH+XgHGaA1JVSlWeFTVg
+Z28IuLzOQ4WS7jSJsnXXcsTEysuu7aseoeMyDjtlcnUkJOhKgN8QoHlhckyBwT2
YcGKZghoi2EATcc0oze1qHLqFSwYXGWysGvHk06FBWsiSuS5PDsSBwHToSrKTV46
Ay7fpfM7eHJqww9XfzSWodKE8mDo7p+yFI79e1jd3VTIElTMg3mh+u8gzvmPn9++
zEIHrtPEXK8Q0xp8i5eqQ65nyQZ6Xl3pAFCKgOsGXDhrqqf74i5LmMUzqZciUts1
MIyoD8tWoESZrhWYRTHxRAc4/a7n1vKcTavESdGtGsmpuEWQFsYX8IyFzQzzqeYq
MKbJRM0tn4ul1Xe1r1PUybXqESieCUfE1y48MlBG5TKyA7jDDuCNkJ5Wr6bgn5Xa
l48nb9vQQ+mxEGiVQL0M0YvAHkFJVYASxyF6KXcn02tpoeG6kqOUlPE71RHantKk
XITWItFZlLBI3lkSvWqVg7BPEjpabvCorPnH6Ufg0qWfTCrRS76P5dE+Q/wrAX/Q
YrFpdcoWsFnxSKft8kXO9fUA6jvArn5gRUbM32tVBsIRWAgXsDJK4uWwhdG/0480
OqoDQM4KMP+iAMtQDyR6O55Ubt7k1Ek2Y/A4IY/qfvscahwAwscvwjSgPM+JrlS8
JXXryMKNXaX7DgHq/OInaEH8CoDpo1SfeSYQz9tFBKY6ycAlfKPfo4a1JOzyzt8v
Do6T6A0vem28DkzXuPt8Sv8JFoLqOeiz1gLHb4rUussjjRMf12RcVyb9aR1t26VG
E6+/SIT8BXuK5M2UCzGUx1UBe6UnbFLl/BiWTLGrObJKOdZyCekUsSRrkAXNEN4B
z3SDyuvI94fMio0qN3fue/UBGkEYF1teDEO+0yBRCK57B5HWzvvlPCGjL9xz8mrQ
rwePaY6t0ZfdU/UaAkx3ERgPh7updLpyFDL16okuhJQYDYkoeMeST1p2Nswfo3qq
ORwkDxINzkMMgy/44pEoJbCThXhH7pugiTzyC4z35oSZoFzs/+XZZ9jYcLkYCgp4
3bopSK3pXo9sHpuDmFqhL+fI7Gd3hPAhAZ+Nylbzi7roQ89ZF9K1HrWaDjRknGlZ
HagypLxlxlfDlAyswv+72eVr4gRHZxG83DsDAJrcLJyXzqEMSaprqBOgfZZkNVT5
WGVHJ9mf5Tx3ocyPvk4xOZjfQqGIusnR/akl3bgxUMdNvWPSWm+0dmnPR3cUyA+w
pQ8kUEl3odGvJS3JPrb9jjJ6BF7PF+gaQzEvddbjS/4x2hK4Oc7NF+bcH87v73iZ
rCPRzwU0Tlj0rdHWEEhbmhyNIneInDwcxREiY9vjTYSqkLeoE5VY6xCEttyPNMcY
K0+jHClTJn4zQJldhxULn4uiltq91nUszMHBtRmG6rtFvA3UQc+k7wX6RAfKqPgB
YsEGUJvIC2t9Ro8UOWMOryOWNV7sl0W6QFhy4zm+NYJfYFgwVju3QNTDQ6p7+iAM
A95o+X16skZ2cyEasxNw77/eochm1rXHUEWu1/wOTyQ/qBSiu5s1kb0ABe/jpGOV
9HgtzlJ7dyUiWItOKf69Ww0LdP/tWnH02LVLp2wA/ehbiNu6MhL7kcslLB96GFWA
kdN58TQZwe4499h9z8vUidSk51hx03c0h7uSP1GdfdChC2lmn+rd8VbceSUu2mrP
vkX494WXgszk+n550I2ssfTMXncCeCELfWQ6uJkCbROn3tZ7eITl/wcsbpyssGy1
i+bF58LGqiVbPelhNLKiOcNzS7tYzQZpZkmAo/sZ29/wqOycFXZmNilgsjJq16ZE
5KYScu1cn82ISjhvSiEM1onutcD5P5rAhnOu1lZ9EQrqFaDMTA0muK8H3aJ600HM
DLcD3Pfr1k4GoBd0k/qK2ScwPoI4SQIX4gh+e8diW/F9/Sp3sBSW3BKHwUxN7M2Z
stn9WWRSILkpDpliHg9gJY5FWFffEk7oQZDX5ZckmMOc9qLgWfxo5g/hZyeRO2+x
9gsf64FxpqSU2cdjoNnIhjjEE8pOArgITZC7R8b3+xdlBy+cR9vkww/TM7/8/1sv
EFZqaEs9LnY9xMwqCPjMr7oQlYjILqju1Gnu4kehCRCzVkfKHF3m/4XE8n46bIj0
/6KW850IhBfIs12bmafzmNyqMhM3AtdyirbCxxsqFuvvFbTj2qtQ/W+kPh3LDT/w
mR999gru7XQ6djgNSlV2Ktsn4Afit1sIXDXpT1kOzxmr2uUBRdby+x6ltK0DIQf+
02zg20GoA6ALxHC1BMPLy+kBgJ4P4vxPbEwe0gu0tNGAaWK0BUr1tY2TIRqyEetx
7kfB9SO5GXlj8L7h7dq8KKF5mg1Ohh/oIuYW3Pry8zaz+h12dhCL/bOjnArXUlJy
ysY+UGevMDwko9nCddpctHapYxB/BRPGkzzT6Ft+Ic5WGNE9AIQzYyK8qNVrmCgy
7+JtliWwquC+aeggWFQ8ruEvSvOOtdshXzzJKsU6HcwMpndI/JI85Os81XLlvMB7
ye9UJgq4U/TfHFQD7FkVBWaHP+stNNOf1LUL07jj0TvV7maurlqh0juYAeiMISal
60vfT79v3/7okZh2S04xb2xzoF0yjH7gLA2Vfx7zqB1PENSf1Wbu72JQbrl1k29I
sMk/5SwiQFKlqeX5qrWGITyaFUlxyzId9UNKWiPiQ3UHxz4PUq4JWBAsR1fym+bj
8NsiOZaTNwbNIsbvdQlXaf+km/IgMgkrzbWc+6VhGfDX3X6u8REF0e6HwRWwKPID
FLrhacrf1OnsJatlecoR660sd9oa03IJPkCs7iO40g/ZRXnaKLwh0mwuiQWKpeK8
o84TQZrh6LSW5ZjasK+xGO+tPn+jR3S602JmMAZjIsSiDpRYXnxdzyTeWAEbwho8
47ZSRUpI3QkX/r7XFjS+cdCrnUgELX4oNyt3dYP5z4tKfVPpXpew6KGXC8NwGeAc
WkQxyXQznPt89WCIRrjV1wxFGvLT3vxUQ7d8CZgQiPZ0YxyaBSvpQVcyoGYFJgy4
qMhC779AY16uLiouWbFJAzvJUV/6nuDTr4/MESEhlOSvG6bO0JkaAzi02YffEdyX
Y4zx0VtbOTkL/wsF/EPJUc12ojEq6+0Kneo4MmT7XHVnPz9D5O4r+9pChbZiJ6eV
Q5gp2mygjyCk50oimMEW3n9tYlqpUPGRW8iTu7gK+hIo5NZ2finq2g6yIqIEw/Tb
z+9UQ43QUm/BnWTc5TOD7SXbRFIran9l83Im+qh/UuopCXB3lZm2FehrF2+Z7wKE
Yc469C0ykRGhyP84uk+izMIcqQw5k/9fFpEiFAOyn3mfcVMI3MwpIlhoH1vRezzQ
xMmfrVe/PI5Fo6VEA/T3zTOygoGLGmNFfjmw46AXGTaGC9PVpIFUNBIic6mrVStj
6Z+x8kY07sbKoJc1GxmsxPnrUf7IKECTKktbIjwg+zaVmxwVfp540LVbhy/3hZwh
qpWh+o7emeqKfGBpwhyO6KVX0KyH9IuwPLXTmMxmyLq4YlT8XC6ql3egNjQShUeC
3TOJag03qCyj9umXU1H+NznLTN7SQKnJyHMqvdarXUvUAZ5B5KwulN5XkGyGLmVW
KJmfuElWV8DglL/y7InxVg5n1seHCEuqh+rQyCTQ40ogD02o5/WpqZpvUk4q0NlC
LTza+er5eagyWSPPF4oVy7ZlyOn8cbXzvoJJWiz/5h1uB2hwwswv/APzokVWDui2
afwqYgAPQDZaPODMfuAEguHrakRX8Oqyxw8CK9suvzJwhPpB9YivSw1ymlTz9g86
y0FpqFuFhHDRcmwatCJzeDDBKy9r65v6fjp03FRtkEvc5yblGrKewR4aBfl33GxR
jcI5786MZ6PB63RVjE5T+uM7AX2wTMjnEg3ryDoBCJHCRVDrPHjUEolSm8/q09sf
/Pc0YWw/Z7J6K79aTNwgyV6v+pSlSEqjB9aWezm+wEkA/BgxzFczy391RKZMgA13
Qap74jed1ESk+u/B0w9n2GGeRx04iFAA019xo/qXHaZMJf1iucV7LJ+l/Ct67Ch+
DGjqFinx811tXHwmhn23urUJyn4GzTRluuuvZGl7iDdPEopuyhVNu04F5tH1foPZ
mUzXBcUMJCAcriQQn8GIkNWhonTpfUQx2A9Zpi83xRPgPrKX3WH29cxQ/w/EpOX+
O32D4cpQsyUbQcPoDzBFepSsGvtXmU/OdTksievEdpWDjs30PCJdNx+nj8SIKXXy
nMNPsWjLz5x7TQaBRvGCiQ9HCpCMPxNlwPmG5jQKKmbUuMG8vJaHu36/yPJQWLQU
byUVDHBsGVZRZVriqSW2c55/O/8Xw+zCdShYddaSy05wglUYKLA2j5E36CfAjn7G
N2oEvghunKCQ399owD8cZjx+cthmFetR6CP02aW5cb6HjbdG7pXj8YLeC1occkNV
53ZxWBCOF+IKM6vxYrGG9sjcpBtChhZwFjsYEuoVyYRT7/zxjCO069FWX00lDfB1
yyg9bKL9vV+0DxDfwVcFxaOUPfP7uXGxDnOzQW2+YQpXSzRQkIVc1HtAP7PWIG5a
oygmEoIpFkDDbjT0Izq7d8PNwquIVTrPKjxbouwLFPrlP5jLECl/exS7mv9wWxOH
4YmkC1qZ6vG8WB1mxxof6vDu5giiY0uOLVrG9Vu3dcbFO6dAJgt1erF+OO6OTi8/
Wrj+B2sMG/MhQHOsKOHHTJfouZNOvXCED7cvCaToUObj4Ag9G1Osj2hVtwxhjjkb
hdK0AxoNQLbdcSSWemRL8YQ+shzqc5t9R2/5j33zn2AqJ66PxUlm/4e24OW/B88Y
i3pTBgwYQ6lIT4KX0REqxUTUFcm729gzPE9/h/yjTexk4zaLD+vPiLCsCstaHmVD
PaIwP57JZCvSgT0BSWTC1eufKJF6X/g2RWfKPJYoeFDLbEpjezHQu+Ol/HhoX+JT
I0xbNIUDPLwouKXErqvYJBpJeaHVGuPlCbsTIL1SKRA7bQWMJ00i8rdp5DHfIfUa
lvuSyN3WrvY+YvXW3UIN49qGoxtM8ablCkQA6Tp6dc9QTNh0oEZyGeqKWjQp9q98
8ehqsAdqoXrkM43BjDApVYGFrMHp2KxBQ6nmjJZYUE5yuCn4hF6mS4+4tU4J8/T9
Crf12AADSJyjmNkENdYcpfuhv2CcSuYsb7y7g2fIiV6EMcIQ6Cdaei2S9fyUNZ+D
3T2SH0Nmf+PvjiAd/QsSwzuFnY2VfQq9LUnkrGwV6c+FoRTtuAIKL1iPCL97hPF1
XLOvrlAfNfeNE/GbkbOeHyR6uq/RvKOx7/YFE3jYQ+53GB+7VA76iovh+jrPipRm
RQmkQ7SSPTysiRFLBOkt0+Pcs672AFm7TemLkuoYZc3qKHLXSN5oHZzLuKk0SSL1
9N5NMb32v5UCTWtOTtPjay1SLIz9VDC9A8T7Txpkpxl9OCTIXxoGoiAGJzgMWmCV
X3JkuDXacliOn/4nFSaf2nnGjOfAE0FaGc9NGM43eiT2ZWH15/mbXV+lFAsO4YJd
cddItFhXV6FybAutWcwdulk3swewvVOFsI1/rprZuOEQswptpLsFxA47LDaR5XQy
546XpzJVq18uh6w0SI7aTXZpb8WaAFHDAUpmb/EstUZPMbKUEvLh8BxAww59PffG
0AaTHKku1sXWB12nkkrdwXPCNZkElPuWq/KXxS0NA/ZgOeaF12TNeW3H5r55/FbI
DmtEcry3VSIHeWDUdu9px0SUkUID9SmXttulaXFGbQ8zj2RH9q51NiXVKBqz/OMr
FvyeSx6uTyAqjn8bCckoeXJ5+bOQPTEFnVTq0PzValYN4NqUbGJmCs5QMdVbVqae
jUPxLMo1mT8TuUZoQmzy1AEhLDHifBCYJjib40lyHX/ZyF75JCaDVjHsEZCb+joJ
HGliW57c8RIMRJREhhFgGSMaJeDH0MqZCUygwDEbQ+6aRBOjniPcmsEjCXAdeRV8
gwru6na+wEcSGkvQq1iOceHbwgTXZr9BXFwotrztKHJelwvFM7OQ65giCF6Stf7d
sPFQCnM0T1b5ltbkbfHtCHMulkIkgTzGTxewg8R6vxCD243vnKUG+OY7fkgSLmsI
x4nGerrjyhmdeQeocFc01gcZRkN4Gl3m+zqAD1Ve89ErGFXIB8El/uTwEWIQIwL5
A9C+p0/Eq/16kGZlCSo9zOXD6mf6CmdZp09ezqnuetWIPBIXTTUt0OukpCbi6OaR
CuJObEcPSQ2jpSqOXZwEtp3VSZ4afqtcvIJVHr/saZI/fHgqdcx+iXdOfwfbPmtb
SAOxRW20eRyk14Dl8A8Kbl3yUSrzfYmBW30Itvc2bogkq+b5h8ZMLFMfqYOazmXU
E+yhCS/p6HZNAH0i/D5Bhncq+uMFWNvDKQXPZiZLimB1VCYqHrfFCMNlrNGVBb9c
NCTDAL/zyRT6m/usy5/zk8jtOuCdq9WuIHlMzZJD3ebouzbbJcRm/aMMylsvHeqf
ijeCsrHBPrBAzSTKF8uhYZbGT0+IpDakd/KHELiti8vnu7jO2qA0ErvSVFu9Xw7w
q5hGAXQyLPXKuY1k+ZjJrtLYpB9xdjDhXJE0s0OkVBE3KEwB8YrfLK42qhHh7WGG
B7lANh+LdSImzSyA5T86LCDaF3limPTNGk9gr0rOoJMxdT5GlGpFEQ6SWIQlGIs5
cpAWY9Bkq0Nkf2AbqtYaD9qxMhr0v2Rp3wPqfHO1zFXAu+PQzYs2jNfQAkzVRnkd
73tEldpB4ffFY72oVdWg16042WqBYFLOX84x8UQNK1z9mAj+Pw6f9nmZETlFeWQP
9XGHwTGYI0MTqJs+H3nq1Q+Ht6SwimqarFilnjgr2flfshIjTC91AP9eMC7gMDco
AlR3w6qvyjncn3zc/IsbVS/5ulLTJlE/BVWVdx9j5gcxPSuXpONSq3Mft2GkILbo
uXHGceQjcZ2dBraa+o0WHiWlrTWZsvBfM2S2OWZq7MfhUydoReBxqAF1DsppIKYr
KNyP7NH3L7ZtF+fMFxEYfvpM1pN+6jIailPoJ+pM2E/s22xztWQ6cqrm1ZAcMKCq
xcxhIJjVaSITbXsJOwaxijs1Nzrfcj1EyndoTv1YTi+k4nQdZJsYfAHpet3r5qDZ
ka7ao1f+AhAr6gieFxEgAfsZDxeWs7KyZ0aWXWiKsMYaLPt+1Xp6KMxKbHxhJsmm
lskVwmLMkOBlwt6kGLZW4E4Hu+A8Y8TOwA3Uc1YZ1klyF9a+2k7r9JM9pXqZEFky
ydCBhkiScW7wyNr8SPcsy4AUdevMkoZH+Gdh6Zhwl2/rw1PDsYMDypdI+gUAsFNY
Imbda+ADWg+lOtKEP2rtPDRBOqdiyi0L6+wi73+ihp541pXgEYf05pebbWBzyS87
6FQZMRQLPWjZ4GlR68xZvtNQK155LJiCyXidymLYEYb40qby7gg0xK2IGS2OZ40O
3nXpWqoQYnucIrF2LpQrMtlQLdzDuxXR6E2ftEC//tJK4TRsnogkNtVoRjxJVyH3
NUmKGP9/apoCz84Sn1uljMznFUKGtf9eyHns6H76RPx+rYEmGVSGMTPNk2HdCqrK
59fTPffqB1y+QZ+JO0cZBF9AqRXQphRbhU2YITvE0d6//O4v0QxdcgGpuUTT7gt8
91GHObjaj8y8o+s5Dw9lT9eKdEEAs4c/T1OYXm56PKq9KIeMDV0NRYfoYNXta5HW
x+weXFMcpfhCKd8jOGd70lwIz8UP9+T5AdcuZo9DjN2ogEg9jqJktJSbPF4juO9U
Vy3/j6BMJR0+QUY2jqI9q2/ae/F9Fe6jOzW3iwlm2I1K3yKerYwK8fU4Opn1Xyha
V7wJ3sKWyjCMkXuiUZSWZb/0rUSNeCwn3O4FOYZLIAJVTG46v4CIlSwrEZYV5olw
hItRo503sRxpjS1AD+a9OdV9+INq5sM+nU02wj4yil+Zhmx8O9XPkrxUxvAb7bjQ
CjSVLOvs15SEQEcQ3Kub8LCvJtQHHH+YrJzG5Bd1Dqf1IA8pOgInyWT8vhpgLOWQ
xc7AExFY1GoQhcxUqeBiRneHIln7SzAM3/qROu9MeLu+QYOXqn1KFv3SFolWcf3X
4Ub6P7MXkWez7ZeaLwYUbjhrLgp3el0oWgaNP2KYinQfse/QgFEXNIlApOgaemL9
8UP29t2+hQk6cqXAhLqA/bFUEcO+gt0yOtAKi/JKNpx1o2hhhjjE8vK+NjT+e3xO
bWmIxlWFDDMAcv8yIA6ohKbljOD2YYKhOV4b64H1IBvi5OsannM7ZzY399KHElWT
LmNF3cqVQFfryPBXHZ1S8YLTNYQea+Ke7ONcePTtw/G2Udf6jokUigbTH9IrUqyu
h5TnGsjp2QevqqHITPloZoNU23hIaCujmFg7Hm3EXh3fwEyADwBkdT/wJjPgG0cY
ViDXcOJYyGjY/+7jayUVekZ7msWtcaOBSd8fIxEk8nJYoH4aceCKJ9dnzx3h8nDr
4OMwXOH1FTGNpDmCmvm+WG6SDZ720yjJC4l+r9/K6ExVhbtQsP4ZJ2Sz4qoov7Fe
sDRTZz0MKyOdhcx3Fzajt+X12cJ+V18iR5ZFYvk9cmiNLoOMokpaseYp2VSA0clj
PrfZne5HOtDpRzUvTdxrYGKunw8V9fBFAigGe95gBisyVw6bWI9O5vhQlxSCK3yb
FnZr+BGKAL11KSmJR9EAMm9iNwVDT6fOzDjELhUYZd6Im9BPWjakvosGhusBWzKm
+vzp01pydY09AE1XJ95Sk0ct0Y2sbQz4Mmd1t/9EUXE1Ra618nlhAUmjshaNk/ua
hKZkm88Cr/U1cOgfYQ6NIDb0ov2nasLRBfOw9/rSpaAwi2PLaLBy3zOEwkD+7v+k
36EmpJHFCDamWIJuqTbmVEsTPbmsHFO9VcZDKuCoC2a4j3wiczl+V6rn5fIIw/NI
Dc/Un5+NFKD/j39X2ZM/xqE8ISPm25/9khuYtLEkX7LkgV8skjEyq+l3AzLVjdwC
Hfk/6aUci43Il4LjwZTTbPaKtX37bzXeXcjw4UMQTQbRBFCrADns8NWu4L+pv9Nj
Y1/Fog/wznqgGqr5DnDATaViMOnyhDMMuYNFI6+1Q+RCXc8aBtZsWJP3h9rYM48J
sthE7FnUNYtLhG/ePS6PUgtPVohBijSxqXWpefqPbkGHprmznhLq2eRWkF2GQ0Ae
72coRKoBiYJam43/s4Flf82Ko8AlQo2w3KyrebVFTxaqrl6QdA0nF7z6eRriGyPi
DxeBuMNkoavHYc5rrjeCvAlpjhj86cBnMk5muxqWq1uL+TKfkdgKsRX2UIo29E1V
yT3iSaSsr6NKSpERnz7oYT6+JUtWZPsXtxUgCFj7jm05HeLkq8hPrN3edDoqQikU
jrZpnPmDCHt4QR1G0EojlY/I1vm9HFy9wt/D26DD0Om28It6+p34qflRNMFmJdGe
uPI60pYhAPUaa4RQZyLLAHlTuJdcJc//djDA/3Z1fbdTgsyHdWn3SeO/syNJF6Vr
iC1LeX0Sq8M4HoRG9xQLtVqHKJfV/nZs52aYo2BITwXHxFgDcfEC2vaNxM5Jt9N1
zhBNxIESXy0ACfIVA4mTUcCeoUXSpiByaWkYIVZGK+m8nF3KTou32Fz0rEkMXU7S
FRC5MDpxIsoUtTCC/Kwn0auQkeLmJDZkO4JTCf1OKtwjmt0lUxeGWnKqBfsVlfzn
vD8FdmjQH0bCp9THS+VRFEo4QscEyAPnPydrTAO5gqe2Mv4lCGDyMvKUvHdVBW5p
0A78geaFOKFe8Uer2v4fvxXF2+L5TM67Je0DXDaOJfUCWUJqiJmfY01UKTFDw6Wa
XDSrlZW8sXFWGXYe0P2/Glg0B7P1mkl92k5sj9BqqY4lZtIXChH2Gk8mH4XJaVFn
hIQ2mvv3I4I5Q5n2I2/XOCbzMVww9QhWZckpNWg7LyvsJ/7lU/e7ZfKTbWpSgPFt
IJThFjbx2VvdjazwkzHKEIZvpcuXehzkRFpzzu3JKhfYwjQJYJcUNdd72ZU2rLO6
E0siVXnuF6UrGjVHkznn1vtP9ab6q6C7VtkATsJ4+tnHGVid42wPY9R2QjMC3MnX
Bf2ieBqXlY//pnc4w/bNEsIW19IxG7+mk/A8hC20x4F3vxxNZmC3skqtLmYOnd0u
MPpJgD+fiSYAKrPbHp6szz2XrpfqttYSCmJzES7okLC2lO8zNttAy6Jsm4RmClnv
pDvTJ6bsVo2TJQ/70r84gO1iquV9vtDbg47FIRI9Edb6vU/+aUbthR9dqgYlTwrJ
ECeJF8k6kgnhKkqGKgLAtK6cnqsYNnHRa6yg/SBuIif25WmLpbZzYbpuZnnGP7Tj
CeITHBsu6L4W2JAyPzipG2ZDo/v7qgZXpXpk8jun+pyoSzIMmWjERJM/412NWgEw
KbKyLNEMvFwhQZcbUoaJjXDPEtEr/UhjJXNEm2oep/K0cIFAsqo0yEqrdtl1R36a
hCmDoeAonBLPDwkDTlQmwpW5H+10X2JlhSkiSZDwOnA1ugYVSJ+lk0vejdYSeEmz
pOOWHB1lAD9j3Q7sTHUzfLhptIZzJgqiN+XlcDRYH9oaQcqx+MnvNDWwv2OiMeBF
yImpcMJTbw6QVnN8IxDBjvPJYzRWuBOG45NOp4Wkl5SmGDd9ZiSO+uoTWt0MEafu
ICyOZ33JN+BdTw//HYUE9EMlsjekuxIoeTF5bMMRiKbbhTYiPcC/fCWi+0rNuEI7
mqFoceLuLaWetv97V47VzPocuj9b9PdInnJX7B18HT2HvOtmTV6og+OSEOwsgx+d
7jk8MWU4Khj2olEME0+U3b68LDdfjrNuOdz1OA6l1QkOEL40j4BR7By8/7TVO9gd
3KQcuR6eMxw46wH7MASQ/Gny7rMJO9K5e+2jvcY7tftg9gwuWtARAu5SOJlJ1dPJ
puiy7pJBuZyCCFKzjqO4wR5Nxq3h3LX7k15HQB7Jt4fLZclR/hXBDK7vIgSml9x/
OhBzdQFWXOlVI7lHeC2o1N9ZLcT9Su5CFW4gtGBOJr5+pOVpHE5UcghzVmsm7Mbm
mAjT+qUDv+NEiKY4fuvGiTL+uS/xAiddlwYJD7fS6z9RtGHTKiJvqnb0p8x/IeFX
gqhYlMIL8oDz0Ydlre3OrrFoL7Q1pzV2fZoL6X/m/paz2EElpspHYGSbmUdeoFix
X583oFyDQvjz16eiZAyZ3q7eUHHjALbLwKSKvDVbXNW59W+OOM497sDZYVKP0X5w
LuB1Lz2RlDrm4hzcUqynOUvnjfXDtO+BMtLpKqmItoNbCrQTNCGf8Wrh0x5EdfPK
8Y0rCpNVqZpv3w/rJTT2VOC/eMAB/RUe3e9svmZlZ2yzAU3rv7pqEDxCj+uoa9t8
AIoZKGTJ40ybMae+qnZ2lJMjJLtG67MKSVOOnpri18MP68EKfsxINzFckN90E8yn
16i9SLHGU4DKWtlVAJo7nWPumDp60xCGzP351/jkPOFdiFmX7RjIRI1sJujJY1tE
7GXTOWTDvGccI0lIwfH920KwM2zSMEhCH8iZZmwYIRAZa50cq/FeQYG6niFgBY74
OgCFnEfllXzoBinH099hTPG+PTcU87XQqCL0uQJKtek8qf7fyR4Annz4YjJcSWGt
1wCC0ZU4Ny7Qf9jYdiPLLkM3ym/MDoPC96qBii9fcTLc3jB6FNWgWMyCD4brYvC0
7+1s8hKTkZCzy4KcFXEqO0o6+IRtH+TKnw9O/B2sRM4a6j1oBbPzPXZgxiphzqq/
ImM5L8Ev2W7PZR6pkYQd4/Mi96VRA4LB2keVbxn7Sjk4kaVgLvKVvuKEYO/bua/x
CWoawqWor1pYAY23pkMSUO2Quz4mLAa30Yg4QFXesu1s5/eWx3xoHhQphAcqvBNR
eg3qesduc7DUG0unFp9GOK4VegOKcbjYELs4gpyoOmiVUta0yMCxDTOG/dqrkPeO
sTEUk37F4tWEaK9FZGrvhMUfZiUGGA4DnauPV3f6YkhintzqcVzl0XGwbL0G6eNq
jn6rfT8JH/fzmmbeW+aoGfABzivmoZVcjAl0xPOCHM7JnPPgoRccMjuCf1WxyUeA
yols6Ku7xGvit1ZlSrl3iZdE4DEJyCU1ssqaIry5UtGEco0ecAGzUyBV5tXp3Ed9
OGRjIK0UUOdK9vuF4c0T7NlFVrRV+q2Mj8PNNrWN5aJmxi4GRDti2tnPexduA+Is
s3UW8jw/IpvzJB6sVCVq79tO2ht0FH833blcjaJ2r8tFwNBX5U17CvLe5if2Ss1z
+SA95kh19GTLvY8K67U7VaWVoM1f1Be9Gx5xVq+h2hbFkdHvuGOCdUGs4Ur/TqeB
t0TroyiMidvE1Ha5A5jHKayoK/XvlQPm8ERWRchMmrna4pmpT1e/WIxaAnhrdR1j
0B94eWcRnS8gRVIJgFdEUTV0DPD/4W4X5eU++2LZhdhPiRUOBqGD+DagkP8fdW2G
CriX1yorL5yhf9WVYmVDyEW7hAn1ZWlT2aQJJDREk7ulTXunE1d39zejj2ibfF5z
cuadlMz7gYKPcV1rQEh4XxyW9rKl8bom0qiD7tlq/BW7o2s9sxzEwVvcNlKH2FeM
NaXDpxRWOEyPjKDN4Sc3e9wTFPbxqKzlIoYqHF6hLM4Wvwu4Qg+GYfdOimr5aT0t
MPa+zc0dMb8sfyRW+Qyk8CDh8VfckcfYmLwHRuRFyPZKO6iNfuOqCHNspScbeLSE
Q0uY4wXt4cKOjCUhj3wIsrWNQfl0w+yUbYuDfeaHCoN48MkwgRmBBCxhLQlouPpn
QsiMTYB6NsjnJJoU7/4tgbmQr7xHN2NL6dzpiRYJ8Wa5n5OQ31/shBPuqtt+ZNa/
awJS6Twfzxlb6mypkN9StAku1fzHyhQ4ORU9Ns/djcnFUVjVkjh97hgUj4yeqNCo
7LRXczGhiIBZ652rnnIhQFaqLJUQof9xe+OTyMiUWl5a6f/sXnI9lMByEhcZNtu8
Le8XJcjY1n9WiGkjWdUu5PZi+oOsWpZgflX+xcofmYiDhAm6xTNKZ/9dtdEm1Vfc
QclmC9qu3ua/ptipUWyVPXX28etBqdfFWEB/xeew2vY6kNeMtLPKyqKGq4jwfZK7
ILj4p37FjtGh//rCZ0elSvhF6bG6zyil665niqnQMDMgpGfzzWh2XiuAPEOD+cM9
VsJT9O5GobxQdLWKMdxgpYk+n3VT3l5eASUmr4Tdv4BdPwNVVdK1wSOjulmj4e7b
YwAF5rFFkBSlVgCjSbUIUhoVW0IDr3SLeJefvGtnpoxXs0tve/v9QNTY4ea7sC+L
W1a8SDbAVQ/VPzD2mOqEaLHeHRx85+zUbO2inlPsqhQaerqp21zGB52T7br7GC0F
OBuHNnXRR/bAS28ipdsi68PvNTTkrgWveGGInEJtdZrnOum5aoKmIee6COjBQJah
hF4gsXHuPh30F5VYmb2NyqOIQasQIWTvnhtBM0VEG+oF118CnVWhryYYFQXXlzYm
IkC12sNW4R9v5puZ6ajZZs69WY7pH0q6NFLJ9DAYI6T96DnCw7V1dtkGvlModKt0
oZOrXRFrHEVdUabs49vkBty6pZ+2uxM3ldcvTDksJruY1edbFGetzj0+QjZPgSZk
Bgj6pjk0qxcGFRpBKuRtLHuIqpFyuvDPBAV1Uf9H2XzbbSgPVLeOKsRYF84+AhzE
YoUq2UTbjvtQIRV8VEICYV20DJUF1MgFBhg+rb3X4cGhwcWbonEmxCOjxztrFWSj
+qegl1YVbvk8jMFUxI/JSke4FT2C6PExVBzDBVqFZftkJn7xDoDyKeLKaH0F7I7I
/PsAhTeTp43wphgtgXjakyHnPO3Q3Rlqywj8kzpLRh4fchpTjQ5QqrLPP0+bjZPx
lmiMtVX0rz81jbBe1t78jZyZlEgnZSGt5M8OUaVNaPciYFhkn9JB22SKFZJOmvUU
aoW4nw704kKJsYKNs6dxUIW+dvegoYF3rJ5R4iDbzCzsRxxmN5F9LU6g2qbW7FWq
SSYehG10nljo5mP3/YWRH7PqnOlPj/U+YQMIwmpZp6YMOy2RmJ8vKU4fE0mV57zQ
GC6QzSTZcwQc8kIwi1l38RtMvlqRjGz85ZqLtOeMAuEXtLkadwDjABtuMyBkzvSw
3omYbYL6dxijV8FBFrWSYWjHmxIw+OvsjMpCyNJv/UB8s5L119qIehKTzNQh2Rou
W44jdaLVrp6GsekqjvvzcVVOFHW2hSSgPW52Vc7kRIhZfhZuZQxKuMN+3oqeyYeY
Ttmb4LwBqKFhw0Jm9q4a/zn5DXCVqubVJGwUrp10FHdC3D4lroPBeyCAnsEPPjM+
SMYC563pQ1AUqNdsfQS1bem1BnrwshfQNx0zEu+RSAeg6w/TzHTVVeiomNcWieoQ
G7BD5H93rz8oegpqcip5mD3lytF4eI1aKmS2Ak27qLnt/skAS4PqOS90X4dB/0JI
6zB3tnuCRt4ZbVDet5I3JnPOy8GiGH09c6GuY6FmT4eKOB2LIWUB7cA5bSGOQopR
c/zzNv057ZQpZaeQ8JJT65ooPcCaDgNhpYs9Ca0VDzMzy0Hc3A56+XiKZHZBYfTk
GjraBsXpYSPdWvOf67r47IvveES+GH7gFuQJV1TQulk/C51Xp382NdvqKYs/1M85
fIVM5cuE4ODGnq1sNdifHBPW4NrVZDWsgrk8I5Ld7zJc9BNeVSCrE9/ICXNcA3H+
lPooYr1/VSnHtIUnyCFA3NG0GWfVQhHvtuWOdYheh7wmJvAg18vvh1u79h8QWgaP
sERyifnZMYVgMMoGUH4gdQ/APlQlFGzw9hNi8FubJI/uAiOoJuLpMvtS7ueC4VVD
VziG40b05HzuJXPsLDCuCW9rfULyLFQDUR0i8VBsVsBBakdJtMYLogzpN5QukQ6s
xeNhm5lt18lCadk8PItyrEsX65YWzBklCmDlFT3pvEsRX1x+CedPXTG0iExEp6bI
m2rCt7A5GnFK7FlocD0q1jssn0Q7mLjHzOHH8aggoTnxjdz6Ss1Vz/+zUqAm082d
8o4VzqJOp97lR+VAXlfGqyyCYAc0+tpHR9IC5ZnBd0g4fwIjiC6+nTI8Qeh5XKtk
eRnEeY7KpsMA2Kl6S6AM3k4uBecsPgW3A9NHQFUZEkB5ead2LAjPh6vyCUqiOwM5
CoOKmv64i/G9yk4eu1kSaIjqEi0DmZICFQWYVEmuv0F7CI1yzDzNrhgQfTYfC3PC
LurAWDMAOZTwPZFcHlRlbxDTiFH3dKQ0VsWBdCTfqv5u/91gAxieSUJ9/6gP8Pza
BzDyyGWk98Mrfpx5kFDyWU7B+BumpddI2HBJ4X9SVDscIr28LvQPdhESKSfAVmbi
tT1t4YFWf+aVCv/n4g0uDXF9SPbwXSff3XNZ9xhJ81hU0WhXFaMNOAPZo12Fc7zY
lCebQ2w/6iwXkUZrqwCY3hl4MkueNrvDFJhMWS6BvpSEJk8TKdkvGa7KI7WaMMtD
su7P9TFBWnOFvqOz5IHuVMiegEd6m3x1IaCwlaLEhXFUzpx02Mj9qFjvnwrZ2pbG
iu4lR7lCEdz7OEVO5XHBxvT/I3NiwysonJSGIhvvdtdKPnZxUe7pvr0WtRk/Kyi2
I4XqWNG9A2ee34jqz7nUbMFcwfITAZIWE7jal53phXmmGkKDNVG5CJDCIg6cUAHD
qIrogjB1U6IbHt0SCk/lGOhkF7NFzwIqX3lIRGtoxFv9LRk0AP7Qtzc3XIWeQgvl
pMoEoY9Z0Wk5CRKnAkIjYr6O4ZF2FYd9knFThzl/8Ucaz74lEePH1LJn26yy5vL4
BCf4dMsHRbefoNBd6Ddaie+pdSe6wFuOxM7WnE3+8hCi4qsjYxxD2eZVPDSTht5T
jeatSZ4ITKBQcednNM5vofAOc62ZtO9cVDvbFBkPUvRQxAvb5xcf0j3OvfP5+pZF
nUczu7gtpCvXh3MiY0BXpZDty9eLlcQNFDGa0T5FYATxdR73oMfBuY4QJa84OKrt
svWH1npuQGAn3draghdlkjB11DQPDE4wkqFXeg47jIRnoXaQjpkc69Wy+cLmAWiD
WCgX4/p58i2JPHwH/rUotV/JFJTcP3QISfFHMNpLmqaqSJ0Q6V94hD1ky2vhlrAQ
kgXHN/agCtGMP3fjXDI4lw7kU2EpSg5fIYrEM8I3HOUNbmBBVmfikXfSUfmD6rCc
zfHgUNWnd2DJuXzSYRejtd3ctrbQ8hU+GqMApeW73GEZ/W4TTe1VlaS6jiIZOiz5
ylZGg2IkpRJ1uqj1kmx0h/QTjU6Q7viVAvfyUdNm7W+L9MYuzZv9Kbbki7UezlYo
0MBvkzHlbt3ZJRx6VKHmkvDhX/LkKFlm02K1zNL/jvVR8zHPSX9sfVV5U1rdfUFm
ndSDFsnWQRMT6Q+sSr1mpJCArWsLJMpfvAAL5AZuUYBFovly/oGIQqWMTT18KNmC
nXjMknrje+O3Ciaatdn5xiKo6Po1m2rzg7i8/m4Y3KW4DvF7cJPWd6iJsDqHHYkZ
C8M3E5hgjX0rizVwjijlq1lJDUzudVSYPIEfLbumXoZ8keD1ideT9HOVDU6PgGi4
kPyh67pS0dXE/gONVgY9Zp9nR/DMyKmx8nLpq4nNPQkBiPguwKBAd++OzaX2PFK/
3H09NMHCcjmo8y54odoVJTd6+NX0o4WkSvRaKk2eRUbpoR0I7DgeJoNQM855oKqX
Z6Z4Yg5roVFVpeB/ekKPHRA6quZ0XDyx+Zz31GhN1UHN7qbB2TT/hAacGaC9r3Ge
seGrgphpa0qEB7tn010YsFUcyQ6CebXmJr52nkluLWtdHwU+ZurgHkkffwyVjXYY
JCw1pqyl/HgaRxxssXUVCCeYjciz5F9DMaIiRImv8knaEfk/lP+KOJvA/Ta28Fwu
li4uH3vq5uMSyYQ66L9HPTB4LlzYDKVfif4di7z3tjt8u1WRgpY9y+kbFT/GUOgP
wUUM5HZY58qT2ru3+EODgQcDiN/429zcj/9yNXe64fyAFVJW/RI4Uz7dq7yOrKJF
hM9GYW5PTqR/Np5DMigkozo0Q0HOlA7bnMcRtSqMg1/VgjOigBwxzB/yxDw4YhHY
dTbtz/0Zc+45EZ/DJvHFeeeXkCCycu03LQbcMLxr/D/kNf/DppI/+XnJnCmSEBJy
KPccafzfsb/lkHnkyf8WSZuz8RNuk2xBBkINsUoAojI8lwLTAFiOGGyzQjLd6kUG
wyLLrDPI/SqQNUNJX5FAtBz1tzPvvisuSs/3RxE4IRJ1melEgPBxysuUrlAMeLAW
SMoWUoQVbcc4aoCANiryB6eeGg89NFAvyfErP49LIqe/TQQN+uzfOhcy8lVbnxYf
9AnLSzbZ+tfmUUEtVbKRuCjAU3XTHg6B+DCnDykdHSUTuo0U2xJ51WrDckxo3sw1
QzcY3Bj56UcJLnuGiFAwzNddsy1skgjbOd5qYa5SWv3ybdnwOkTQlFGtrGySB3Wh
KpvrusgxsT1c3GmsI09mPr1e4pjWITg+2bOWkeGequ5K8v/asL3h/iXKFhmhyFfR
VdWxR12CO7uWiLDjbgcUS6J292rnWnP6IFAzL0+jBMRV4Q25lWUbXdI/IVUBgzlY
qfQgQqg/lt2R9cDH9BKneyF38uKpQoUdqECqOQNrgQ6eddPDikbwKTDfLWt2eMnM
G+yVmsRD+e8QNy2Qx9ldwRWnjdyrrZzs5+gd9joDwRlLRk+NM6caj5FYKuDOJf0S
cpDWbV6eq8nmezKD410f7N5ybD2dHYqYQF2mnxS2d+wa57UPrMv5tLltJH5ORbCe
2npS1yWY8XPv/VEg8TJV+pXkE57D4dIX3vilXnX3Ik0nEX7vjizRmjh8opilSajg
ezafujsO6J2NbvyZYRyuiD8OQL6Onp8hcfMsysRKmWo4pan2ehJI/Uy9ri2KVDM0
gaWu30AaAavXM8+JP2RfYk9W8/aS84H8qDZqjs8+5r0izXRchKsiKqn7wgsXu6j1
Yy4XD85tyG4uNTMxfymn4ZvAlV+lRvns6R0zTcoQT9Uib02uMcBZvTLX8urxk0jf
BvYkx+EOA6RfgI8/2ZUwSBR1Lh9hqRD+rLx5ap1KM1mvZBoP848w7CXhYYsEiA6X
QmsF/plhYshDaiyfUvLtIF6/Z/Cw7SG+GVV053jzXPR0AAd9VQwYuxOyqhyK6I4y
z2iTMgsYWcQGZwCptCP4SedyANXRwEcGh6aIWKq7mdRfgQFkCD5u4dBlPbv6/Dv0
hQ6lIdx2kCWI0Bhegig27cVRHZkASSf61pVTs+sgKIzb5mR76By6UTSYBEApl2VW
cS0mdy9+MS0voPu9uFak+8EfvflfqMCt6umOZp6DA/8Pm6bK9v5V4Wzze+EkcoSC
triyq020B/Y9/NwPBEhMOd7MBn1WLv2IE0QeJxRZFiRy1RVXJ/C8JqNpyo1zeTFW
zGuWwF9vOPPXAtx5vF+gJjAXp8yDTshX5eH8OB60cz7bZduWy+u8swFtpvOZdJN6
Dg0OYw+7IPgfzp+gh5WNOnMwi3yAcJcsKbDc2+aNOcvuzrPv++J4WuWmPiA+RKzN
HKgi9JM+Y5efTBZqo6w0Dcj1zlJor8uvWodJlZQ5UIXpdyxvvfGdZtg3PCtr+qre
2W98s2j1lmTvfZFFjADKC730MgeTlg10DvtRWF2Y4MBvjaf6XgfSC6D6ClLmvJMh
BEj5h5f0YYOts3LdV+IKFG2CQOA/rD0cwxRy7GfUvU7iJgTdaJjeqPd4Z/QDB8/X
bG8lQG3uqlB/j+nAsngATuxX+m1ZqC4puTRqm9c/gB++omVsLxfUA+Ofi5HLzWEr
X450HI3kiRzXBYdlquemGrK10Zid64VfprovdCOpaqmNFfX0Jasld6SPGLLJa4nN
bjJZqhdgW49wU+nJJOKuxHnL5hqoE0o1gRsHbg7NOYVMtr88wjSNAYj357A+Vsjs
Wk2w3Q2zWO+962IiLEY/uk5WiHyTuof8M/wF3Aiq5Tb3Eb5koGnlMtgsqAzHw20e
5UGHfnwrZ0ok5shmyrs5KQqYml6J0ck3PInnLVBOuAxIxc16s0kAuhsNDCgUjgt6
T5gNyfNKqCXmu6bX1SqM1KDM8XkzlfOFxiD5KXxSxMh6ogsyEs9RVhGKZ63F4qHg
OlDwz0h2qg2jBRTgvnCotoLUfIEd2mhsseM39PfccFPXjIzgj/YrJFT7lmI9jlBV
1nmWCvf3JUi09RvKcc4rub9KV/4Tsecq1tD3/nU68PmchUGFK2By9K9UWlN8jILM
xZ1xeWH/PhdL4yYpBlcniqGnwVTxG8tYPt+MGzw5AyNgwWUFIle1fZsTI/KxM6xi
ocKCfagou7ve41fb75G1HngJrxtJJP8LSYP6h6iaTV7+q/klGlRS5W0kxED9ibj2
om3ck4g+MZrtMUj2dg43YoUmY1jyMJE/wSfHn6/1QuLuJhRu4Xjy38PdhEI016wt
n/jj1QepN4LFmnFc3XHDU5z0f124mkftp23QpesUZiM5c2TKtJoNL4qZKIX42KYZ
pnOx57+aqRY2APZBlu2oceO2/T3XmHfwviWzujrec//OhC55wNI0kNnmg4Ole8S0
oreMQgw/CbbUh4MTnNGTco32yGLmu4/pzkaByH7XmlY+alZQq8KFjvKXLxpE1FrU
+NQbouAb16NLD9iwioojTeUC8o5L8LYKTEmmETi409XAAEOhAvIONjj2KGsY9urO
40vfkTcYzfEWPHiCVqC9DLbAtSjTLTrQv5WDFXoy8XmPpvz7RCgRzMjiHdqxpwJB
t/6OP6agRi/3kcKXaIhJ/rI6931oR1Zp0vutDVwqDRjccgk8Hw4Q/eEE/oX8a1Sm
M0zU16UTCRhj6lxoZ8BoVnQuPFicHVo4Pl/rcREkRYjcONhMPJwg4NxKImqaM43e
lcpFbMLvvsj6vIFHGbr2KpjimPvpUOQtoGfoY2GXCiO4vjwj2ocRg0Ca7mN9EQle
bRCVMhSGzbHIjHPRaYFApv3HWKjzXX94K867pEIbkblZ5MhL235iZq5op1B5E1VW
sGTq9N96lD4h0GXpLxR2qkF/ejeIO8xQ7+ItRfqZGwxAtXOnWu+FMCnF97kIzM6b
awxf+1pLAsC4q8Q/IkjamNbfXXK+fomvNTR6LpeDCBcgIYQuXEFxh+P7WCJeyJYy
G/vAd+ubNKipQ3DAA/dxmOFqxz2c439xOfS9zrS+J+aktjwOtAMJjzaNJHf23QC4
pdxeeugXf65kh4KRPJoyZ+rzcqO+uaBz5PwftjKItOSoX3diB/y+dXt/cJgkC12p
qlj95W2DjD3Z7zqD2f3XwdCKqUTgz0LImblPezpe8fORW9tQkHpX0c0PrZ3uMBVv
gbRXSHUbCKvdzls9t5YOa9JVgZw3ZZojSGtvSQ90ge1wckvXfjNUTQnUWbkk6yad
h2Ny9cSp50jYXQoam0rppHjshTzYgyKLhbFwqE/XxwYUpijIUgRn6t0iyg+HDs8a
PBDo2izvuivILswqBWFdCZHD1EKbm9FPjB7QpTJKLYPCl6WhrsA2uhNHlAvjJ7Z4
l/iWAjG3XlkvVYgEoFRxZMV3DAOVLb0GzvU6SQtg8jGWiq5nNhEVSt1od6YgV0VR
ZpaSdjWWBo2yVUDy5sSg8pLMV6BGQZsAkRvBpCZNbQXK2xmM4fJcJFZJbIFLGz+Z
9fbPid+3Z6YLr4zBT2KwtJEMUB3Sr+Q9yZ3ZsDFl2WDXC0O1TuSK1OPvCuW2myKZ
VMLOlgkblsmepQiyCUMVclMPA3FUqXpbQ1xPwdkzuQspSK3KIQFMSM+v5SkS8/5g
nVVOUSaRVtb9vkLlcyXxiXPF4KE1f4cx/6lQZDkndTz8gkrb2CPV/sz4XP8Gf0zW
pWH2W+OTBhMWSBsOQl1ZFWgSYOz161NdEfAaW9/rImTwcBbXa5wIfBcmVmnBqS5U
5V9iUqgaiJLn6jg/eSIA9ANTyF4T/OO1QScupj37Ic4//pPH08GhrkVR8zJ0MFNp
jwH4Nbv1ix1GqNLNdsMlUfYmp8HmWcOkG5c/vUc7dN3CK7Y6W8zMwOuUiBfdWzfZ
MiMRmF/wAFxSRdb9563EjWM9N7QN7l8wkh7jKYx2UoRs+/huRCx4HZhJs/ULfRP1
hZ/xujk4KMdLJOb6CgxWjgq9cDRb9CST1l8OHt0Aq1Z9e14C432KDTIAmmvScrLE
QOuBfDxbE4seoOwc0oJQSiqcEThW2dD8wqbgPwi+IlUm2gpU00qiwerZ37lud8UJ
CU60F6G7IWuDoCIrgzgY8dqPoT8jxQrqWD5vUI3vqkCtCHQ9lD24ZIITXke/GP8o
j7Z8YU4Bt4eRvzilWFx1m6guhAfrNuSzT1MgWdGKIEm2pT/MkoLeHoxk9jIqOIDV
VU9BYQaIJWw19wJxsi8xM8CPxzPrX6NAkKSsBzK1mz7uLEfPLh0aTGo/vsAaCzel
/LLMIkWBecCyYVhspPU1CBIjCZeSokl7aWF7CfcXnBnDVIhWKN2ry+hRzdhxxKtj
dg0XjQYJQJ/y6a/NzExi1EMsHbQzuudI7gmoA6vYET4clk6vEsLiiKCryVKuvSrw
c68JIwtu1/1+TmMtxHHNNWcV7UTsQ63s1VpSdFEcuaNp1sbIF+9hkUjyNlNGMWb9
o0ml3FD2znBMlY/1fR/IJyp+41HkzfwF8BXhyPoxzouBBjegk3myq27OMQwQBndc
eRDTfRDREXldh8dd5dtk1OeDnyKozMDYqswe1uu3ym91+3oI9hAPiP1IL3M3dux1
JnEovvIcIb+a5Tpz2xc0GZECxIh8+ii6NyjB6dmSG2PfIlw0Yh6bKEZ9xe/LJihE
UQGBGy+zA2ET045kTFqJTVI9JsE3IbiMsF7EH3V9VEYSKHrbCWco590xkEwvBr+Y
9UHAc1fGYtkStfo8osx3yW+BN1sK3DIL2IAAxPvE6nD+E1uur7hUng1le/KN8G+n
sQHZI94XPTUjOsxaPAz80mKSPFnUNo1srYmy0831vyEVVhO9p1Vc/X1Ri6VZGJmi
bRniZLCn4fa9MaX5psoZFvafoCPta84JEHsF1+JGktktOIarNE6r3vE2ZIEGO7cg
YHm8T1hvyp/AFYhhi+S/PoMa+C0Fmq/axH7Avzvv6Zf79euWs92nDF0jzMa5YHpU
vh4TBm3MfsZVc+fKAFvHPBX65DE1o7hH3jaTed8SPyDLcVKeLhv+I/r/ZUNdEvya
81/1k+XvhyugTjtqoGoIDT2i69CwxD9TMKkg8Bbeugce5uAQ2OU/KRhq/UdPYfTD
4S4RoAgAnUMjG0+20kuFk5lQqd0sSFSCp0CzX5nQKRQpHU5lKbX6VVXVlEhqw2MF
It8LRBY7gZaSm7tCDvNLbQcoZ3rWYXfeedr8s6uFOgmxP6tde79e7oaeuIEOMZtf
Vzd6mYxj3eC3ZpKSmvqUR6qnHc8uHmMDgREs6ZwD7dg5zW8lOCV+I41SuwnTbI89
bgyJZDj+QJ5q1HD/RJ0etBADD1qkgJcjNCE5beyThOvfPrsXTPPszf7j78EJEAW8
kybml8LSFaNRLty/7OXtCVQAHndaohq4dIwAOHFjhGPF8CamnLt+pu0JY9f7fYO/
D5dgE44xw1zXCJBG5NU43tKCH42TJpr7fTIxBe5vD91kSAAMIfy1QjVMTRvVBKPn
22sFEkEZvQgz2pbMepYwJCG9ir/sMWbk3tEDs1ulrXB6tOgd/g+cj6pJuY2sEHvE
9LwJvy9Doi2q7MYz6S9X9STae23nS1gqsl5Byc9jdGTcWW7HevZS8YFSz/zWx+w8
ZyvdgYmxoPPuH5MC6Q1JkT1epK29he6GRTO30Zb8ru5ngDTYSzU+ZYnBEpt5hZVM
SCo++jWQx1OgFuzZNlPSUklwfkQ3uk8xFFRQed5G6S6GOAR7a6AmEejlF5YoSR2d
dbsFR8eO+P0gC95Udmv3AfUD87Ub2o5T0EPsYRareuKc695Emy20qdcGiTsIBLo1
XZygKc/sxlfpwkd+AIu0qWu4qDkUsvQ9tA4M4fzPndzYk01VyWfLfUBlXJdF1WIW
AkfhIO31/PcrAtKkHYmmsX+XJh46XIzMYLbQtWtvnWLojdV0C91b5IwBy6mkEqj6
uUtJ8py7e2+F/GAKj8f1kdCNNgAzBtGnm290gOznB1krnxA7kHMfwwAgc1As+C8j
D0VFaWhP6SbhwDdep78TQs4TSXsyTeA0vF5r2OiMZ3nXi2n2Ojv32VcfOI684Gn9
cBAL02q/1TiKN4lwmmhnZUaV6l1ssalHA1pc2K7MAdCPELa8Z4ba5lH0V7lAVjE1
OGmuunvd30OILoD3ZpWUdf7d6rInFNoSOb7a8VkYotPrRxhkxsxKRv1LsPvZUH6j
SSU3xxjxDCdfudOLpEQwTSWh3fnMZi8nZP6uhQAlWzwe6FUa7RYUSDjs9SVxSlnS
xiSAtaAP75UnYvV0+8a8YaL+k9IeKGi/IU4AjHLHRoH7+sxYvBp6DOU/PRaOvRji
iUWG0qDr8VAhjt7syrcMjqHQ/uNrm0++4w5e/Uvpt6InkH9Q36z5FHM4U3rvUDoF
Aec2PS//S8XcJ4d1TpbqizBarGcgFkU/D0vb3tr/NGUrIvWR36J4j18r24IlBN2Q
djWjMTfqwvtTcAK/lI3OhTXf9NKjvakRnnppIKKR2Yki/FNSRxzjimj2yZ8IC9YE
qt7yyTcXRrxyhIzvXpoFcQr5SLf+OCdZ5Rl17PoxW6IA6tUkvHRiUMUn1bpwX0jB
z4K9md2vUEzJxFbYtlh5bypgbwiGuO5SZsTT3GehaLReET/Kg1cpbns7IAfoNQX3
FLvjDFuBFhu0Ah5kwLv3SntD6gLGbVffWe1O4rdhE8PYcJAoEuFq+cwCIOcPLoUz
oR75Kk1Gz0+kzI+j9s83CPI/11d8BaGe/2YgCwp0Xm/tVQpZM04LB6Xre8f+X2u2
e8D5T+nmm6/BfnNQsEss7rUgFfJaCkTYy2/AJmJ2uVl2lmU60XJirdt7inw9QwOM
R8KtQxjYaEx6dy8T3bYXupqcrWHU0NollIX2HwmhRJxLUfbIdoib6LkkYsDKRMM1
DT/LIjoBLPPSXmkbrhhcYY98mHf1k2uokW55IsML47J4qEvcKQUYKvCzHDfOOynN
hbVhS5yQPNnjLuBpUeL9gRDRRQoOcGQS/QraKsw+np/Y0d3x8eenIxgK2ddTc55m
RI1vsmkn5Nj2BX3Ji4jAUX7Nw2ipD2hzpky+WPBRAos8DtE1g/hEi4TiURsoNgQ+
NwMs8Yu2ZLspfMrMjQZCl88hbxGJfcHATeg+Do6EWZ5LRlAIy3LM93jjavz26ifT
CNRsB2Nt+3+qbyuTcIkbIgSY4gcWBGOUDGnRDxODsf1/d7FPYBVydkvNkv+3KN8q
Z4LyxZT2pESwEgieT1B9tFVebnssO3QgxMa0jafxqAJuiP4z3kobvtT0LfxHOsyD
I1Y8RyS1bftCFwVJeMYmautddAeyOvKkKdbBeW9lUEQqOkzrPAqF63OoNr6Xtixz
49qvdMoa8RzZQtGxJ2Wz48hMKqHCgHivu21cZqwr1SaikSIgx0q22e19XRiaNsup
f2nQF7qb8tkoXninPwsMW3THmnHWQApcDOZ8zczqm+LMK4NZIvyA/nLVs6bUTUtK
l6JJpKI1QlqzTDCdmPbxTXWXV4CpQcgqDRq7qu/kYdOvqEjb27nl9ovzPD8J0KDg
QeYBkmYimNOP00v1Fv2RSVaFENk8tabG3HaQFNv/DAK3lGTA2Z0IuxRP5vmA1mti
VB4qoLQPSVXDt/SxI5vAgkSqSp6/o6DklWpKcm6FlbfvRxmvavv3U6t9nxtBr9Wo
w+5beUV4UJesJQ5Gu9L/clsAjoqiFOOX6/45HcFGtpsBt4dRr7o4Gny8rk1QmwvB
zut0CG++5mz5E0GerL8y3yUpu/k841jVcWp1jJqKHkFwPEHR0eeCiII4XB7uj4pw
7nfwB1Hkrc95pGtWvg9w6uGtDcPdAMZHp8sCe2Bw5i5kwdXi36elX5uh0nAGhBsp
FuNRBb4+qYN/mqqERCPmtOt93dLDMcXj4C4cGfc0BHR1wdeGkD1Uyw+WgCFeQHyK
RcWdAxD3qEBEbJ1MMP5UqS8UEDEQQh87Q5r6ld/WflSDZscKiLb6Q43UVr2mQ/6l
T9CXAivfcYOC7hMttK4HwGxCZWs6beUo6vB4w7+AJU5rghe9wNBrK58dHtAqXQWT
vW94kBCzpMAQkKx0pzo/flJ9ccuRvvbHBZGIqNEkP/NutHUahDmBvgvVJ5O91YCF
PjfKR5QcHSmRCEcnBG17AA6NVGji6UYt71K/7uQk23mpQKc3kGI2j2CYoJ2yhBKH
jbMncI+akKsefOc4okPiHJMAp0A8P0XHXddvWO2Bl1wSALxv9sXjNBklse/sqcyy
8P0z/WMWnc2TB5lOr01OEtnMSqgHaM2iP/gMUh17IuvmKKb6P9eQKg9mrG9i0prl
em0gx5o+SOygUXgBRxr0zWQaqwq98brfDkSJLePLlsF5MsFbywyU498OnMoBpsrb
JCBmqL9dQQeKlHOSjhIT5er565IXqaAY6ArXLVwBq4eU0CRfVjF+ajt+ubvNgqC7
3UcOPmNlCnjYbiRIG62HUhLOLbE99vJqdNSRZU3cnu+lVZeOfpwXcPlWslEojZvD
GZGXd9gm9ccd9qAenAKwwwHfeGNW6mCK7+wz0fFKGyr6PMiL19wxB8aT0K+yDBdp
3fY/eUB1U8AHw7lYYXHaObYlKFi1RO5bQlLy2P+G/slDpzkcpMlajQQJKkXz8MOO
4dgHo2G4tus96+jes7beS+8ywl88igPwgAQbcdVnzgzzzzcOuYTnH0C1moMFu7HM
0pm1ZuOWbtluGBMqsL3NMnO1EbEHRyAc5BFDd2kUjHY0z5aE6mgSJDGTX34iEhpA
1DyBMgD5bnpXrptIcDT4avH8tWYYW1U5l3iAIQbXUvAHK6RCD58/vJxF6lkBtiGZ
9ZY2GkuUUG4LrY28nGs1/2JHS97JmARie3uhqu84kPD+MsN2f1zLkZpSL9+g08/a
z0W0b55ZlEef8407y4zc+B7fwIrGtwbl8CbHZ2yUa0jMxEXk+pGUrCclx3q8Lu0j
rYgpEfUDeBHMBUMk1p0ImUnTSYAfzcqZEOiJ889giMJRJmbQ7g4WodJe/kHB5miy
F0a9bGlt9Xk5iej5gdOoOiCZhCGuvGwO751gZRt1AV3UHMrR3wCOkdqL/Qh7BAJ1
Eq1jorhQ1trXh2W/o4d2541KTyi3t68C60YqMV8cC3fF8aZnXpT9lb3lc8VhEAb7
rYhE/ran++iLh+WwsC1GSl5ez21KKPVmc6pepKfe142W2XJvNqtySLcDzTtkUNRJ
7EWy6LpdSYoTUxkfZo7pcoh3PGoFcljECiCt2Ttm0UQn/dRpYo/yLkVcqBgRnbJt
FXZGMMlBtwKQpSdPPLNLVMF9snhGodlfcld0iKTKBEw4B+XyjXyiGZaZq659dkFX
4TQadd6rHQj8R6jhSftgx4AnA2H/DPvXYt8UtUo9ewmUul8L5kqR4mPAg4oBmqAQ
3j1u0HyNwdf+NZTDzuMllara3N8/LrjsZzzuhpdVRz49rp1WErkRLCgOotgEYkRY
7F9yzuhpsDw3naUr734SipaZYnOVoO9mlCVdjtkMZaWGRDtYFNMB+IDxnmpDJbXr
408dr3zp/x5t/FyEnjjgXFRZ8UMjQgOmzWiPExnrzAGa3JK+AGgXfwmhGjd59Lqj
cO6g9CPR7AGLn/T3+qlgnjH3JcAxHRiKhea1cY0fGEkz0ov96blZDc1zzp3b+d56
wjbjE4QSShVMYbHmEAW4wKrE7UgS7SWVMUSiqCWLc8iDTiWm7Tn+hdNoydiFCuR9
TlD/5TK060lYT/EUxzo+mOw+NVakBRRdpQ4C39nxUs0g5PLWgZLx5Zf7pKNd2n/W
P4jlS1FZrkqd1zbELQ27iGYHqVdvrmhQQhuwas5MMs2Y1lmiaMf11bjYLgoxDoGw
DYUEy7LXBehiexgb13p22LcHz0r9kI/+c9fL+l+hFyrZwbqB2lXec5Xl2kQVl9yT
zLbs8qZtmoU1ni4CcOZT5+yipDsSl0IJuii9y3Xpt8BVe3asf9CERTibjYc84ytY
wA93kPKiNfLy7R05hZOIRNmw2u8uSh+slyagh1qAMflj+NxEWE9JctDBCQCl9dty
oBy3Lez9cwPpGwJQdBjVJvTMWtFPzG0LW9Yf64fWsdO8ut+EfG72QOBzqrOfvZLw
+NB9OBWik/eNOI0/Kf6X3l5eYj065tQNG+lJWMaeT4LC3kHTJ32i4QdOl4xwLbMd
54EWDYme0dPN5U4Ugmjbe8A4lwBbk6IZRdN2SgGqZpZyzWbp72nkVgrlxRHeEup5
anVqO3R3L+SrxayIgkH8QEwE+KRUNJ6nhLXCuMBoWVW7GEXYcCictQzrzXwokEj1
QsvJEgXqj9xEZWl4t3rXu2cHrbaqBAwHSmmnpuhEAyWcnYtzDQZqLhN09d89gujG
Hx6uRX75BKkwRpVJxsr6JQiJH5Arxjcq7SRLL6RBUA83qmA1k8api+/b4EPiu9xa
Z/0tGtLddDKKNJM1VDswF56f40kgIRZRF2e2x2/qRtAfX75lTe4WBHX06uQaYCQD
bOIsINi/Wh1jqebD4gRBTNzYyabp1XpBCrumrg+aDNwC/V681UyJDEdt44h/FYs1
LsEwAqfcOuNGuPLhK3WveOF+WUWpb2vwZEJ2d9eDA7Y+PlkgpsVGsQl06iBZPoDW
FrVXxIPa31/EjnrBcMW+S85g2VB71eloYdPaSyTHCHYNVtYZrfci4q9o9fqyM69a
3aJAcbPmrLbTqZ/Q7dihE6fQxn3hqOmke5LGi1sz0tHsioTks7PFRdwcY0O+3Str
6F9EfXO0bcCpkujJvP69l9WjEAgZ/YUFsPwxZStuRtwi2VE8WibCceqoZEh/Fjin
l8euoW+pGi+ixMpMBxLMO7B1ES7IUabYt/nhbrYtT1pCzPs8WCACRmDtd2Eqa/+1
1USe9+KPMLT7Bya6075azt0EUeYvO2i12nfnir3n2WRzRhQaz6rrnc6Kj/MhlBnD
I6sjTuNQtHddZVwh0Y33R6lZjGONMUZJYBft4uKalgzV/pqi2xyUweES4z+h1Qgv
n7qlESNox+GHSWuoMpHDz/NWvy0aywxLRgMmNVIRF+OA4rMGZ7b/8AgvHnf+WKSt
z3Iy6Y0I4WtCH6bRm8nDGTBavpQ08shdUr/NMn5gJz94VUUtx7C5hv6XEbLN29Ed
vcFsXlTmD546+F/tHDd2Jz/p08CU45m+z1JLy89HuN2UiNLr7IUFCnF2Cia9GQqp
XH20l6J2bg7mdMCfVwd9E8AR2H6YzVMD3tSRd1nH9NiQZaZYET5+EPQeR7ZjQKBI
7Dgd1zjvZg/sgBcL82aIXp2aeXEyteyOhrJpZ6znCKtS8KZ7qA3kKlQCdQXbdcTG
tTvPxjH4MDf04EbzpUyULnftRB3zaF5/3i1xt5f9TzbF5j5DpyaH1pxiaRmnHon2
qfNBAGbW4xEf1TXq18SSIC74jbh+IssMgIxalfklklg8Q3d66ImNMdTURUEcDTYu
u25e2+MmX1WyL+GigP4VM2v0Z7gx2Xx0WZPN9Uc1u605m5egAWEVw0a6fLLLH1Bn
JhkjRzv57SNBZRWzquu78eVwxmrVtv8Ks2o19ynWpqjBnqtErBAQ3b4a8JVvBl50
MU1bm+hDG44GwBEUylbK45/JI/WLATsZCXLGLvnk0dn6A/hVaDk8B+07DCBLsgMV
uKq3ktvovZzdSg4cXWBiKEnqYDme78oDLWxEwz+5SDi+dnJ1+UrymkMB4u75mePE
N+YKdvx96aExIDU/zIp+yx16pM9LKtFv6HlVh9VaOKI4AwkMS1BjwY7D4tv0aqEe
Qls7qS8C+UeClzeZkerIDvKoGY0WQMa72idkh0/NX9xKpQUrjK8ZGor9eEIRkPLk
dbM/r0s6OTHwYpl+wFLI/RqDdQWNE+s6ONioCdGcvJk+jAKXwB/6/5MBshzJhmxQ
owG/yPUGrKL65n6oHV47UJfVLNkgqHVNbmyMeKTP1ddHqfO7FD2iLcYx/66CDUi6
sxMrcuNwibBiX/1U8ba+BXbH9bCkP5VqxewKyOf7tXU2s3LYG/VAeNJ6us5c4HLY
DcNKfRP+gjUP8niudqmt9ArY1UWahrLwMOjKvK55ofaZcjWaaYwUImwqXDubm/uN
DDXm0Urz2WSfbAOWXLpz2WJW1HWC6l5wtwBCQvCDJE3QOR1VsbBiHCMKVE0JJ/g4
kTmZj8MuxpKeaB140hFPqZJfqBUwO2CsDWNIbQY3dGF+YTh0lIR9HT/uGl+1S+yN
ijYHKQKQ7XyEPRRsZ3jZ/8NurM/RJVdTMQmOhs/wEHzkzxk3rWjE6jXaNm/ciDVc
yiNgXQHLTA5H9DkrxoSBXzZJwOfmfDG2Spx9tFzU8pbMad7hv6wOJIPIrasF64Ol
3cXnXb+yn/Xov36OK8xqSMYSDDjl3dJ6jD9blhi2U3mjptzz6PTv1MIyzNGjIfRM
+y/Zl59zb6KCMzCti7+majVfEzKDWOxvtm5dqFJL9VPO8r6/MNaA3Cny8sPW6lAy
W51UFeVQ8uqbP7vZua58rFAtpkNFEJrvSD4qcwK7Xo3uFXu9WqSw/QG0gv8vuxe9
MVydwyd7GU1I9uq+KVAAw+d+5v8MvELNuykXzjjc8DW0tkJxgtBFQhs7FSfz4y6y
cUO07mQwPqoTixH7K48CMh9qJ9nAABPSUfI+iF1ExWVKQej53B+gaVHcGIkOmuQH
FZD0JgIIqBM7Srr9rtT+teikjI57iA5Rp4tVf+BzSLbH4ATZxENil2h2At0lYiRT
LN4FF+OIEQvQb835ZjkhJew4AFFFJz000VTBRrjd85WOoqvv3gRW+/9tY6jOTBln
u6eYKHMZjL4pVpp0a7ohc5c6mCWF1Cy3bJTdIE8FKLL7FsQ9uE7oqL4STW0cLehD
wgEIxMoIwtvwQ942h17N5nXuN+cMS+M6wKuPwep3CrkkmoBVkw2awC1edKj1i+9O
mTQzzBCZdxG8mNnxzmz9R50fOeH7gro8Mjo7ke48JgMQRQNO55xxrdqanFe9A6SE
7An34xRvLFS754fqgcX1ahkg5F3PYvDy2a/1GGwPv3HkxG5jMYvZXVp+XIDS1eVO
jnK63/p5Hl1w8ab/XQN4dHOg5C4fPaPFF22Qe/5MdRXSNwjAJMoH9BKC5djy/3ly
7vV94W75xE6AaZXUGa0/KPPGSwG1zMgPJoecvc/w5CI8s6gv5vUJSCswzoOTnMXa
FCDwG0SL8et14q3jINfYMQjAzPWSYDkAjLkHWgfT+OB5DyZi2yKR7effux2S/G6a
DOwjGKkorkKVrNjBOXiAFzoBV4YIDQtjE6b6CCC+xXp776MiEfkPGRH3+EEqSe88
AX4i1QkuhVQbz3lFT7UiY4EXQtWl338zfbIe3I/CfN4LwxaorNOhYtBiA9LFzSyi
4wZVWizw6JPEs+sEFuimXyb3ymlK1xkn509uxRnVIO1xQ4EOIkjhx6iqCAh7chS7
3QzeDnkj/Iarx+FW9UIZWOqkEYytZBH5di/+5Xb4s2UDLJ0NoWc3UiqBVc9vkz2U
v5c04OMELYzfy3JG+JQrQU9j67tprfnJ1dGdBpVI0s5fOG4ZR7eDFj/cQ+GDfakD
NosuCATSq9IqER1fp1y1CbY7kRC3Or2Nxh5MlfGWMacFWvg8tX2OIOzUnh6OnEmW
WRCsnAFzqCLBpB1Ew1D6IRU5Nes5vTKSi7MmqQQ3SYwq8lFPQtyH59sbjZVgBXA7
7SZecqQeGRdinEqFZgjwvN0WXClntkKeHII2ydMj2FLHEiJ/n014gMrRvjL9mcx1
YkMbnDrBdJXrMKwrKFUSZ3ZvtHxItO2fnOemy1htk+3B/5FhHN1veJhYh4HgSPYH
pb9V1TREoHOwrSZYYq121n8RX5aMywofxSIGxNvM0VzaWLyE/WUjbnmNjAVhCSae
zs6LWXNeWt3C+uRUgoqKY6jfjrRIuJfgM6Itk8IoLQvbGIAeK943fDHc7oCFqIT9
+eSljY9eVyThUVEoCMliO7d44H7W/tWWlbg4eg24BWw/hDXg/cRhgZEZhRohqgDK
WVzmw1ggG7OiCB9HzXXXj9TAMuEMF1nYytdPMJp61WuHiqyB/Rn2jERFuJEUutN4
tTqr+I+Cy3/W3f8qZx2kGfLqNicTkgJVUH/9AQMWWwkEDd48GPDgR6R1vRlSQc/9
IRucqaKQ7VI3GVm79sVdNj+eQjlzKUhIwLpfultUZ4EUyIGKcftkMCK6cjtlF3mR
m0ebXF3ob5GI5e4+Aueyjx+elFUe3oUzNooTbdJY3CgSmr3WdF5tZGoqKY3eaV5D
lIvBSBosepHeo9wuDsvokqKOcyHzBJDjoU/52JuAhQlaV9RsdCZwKbK8P4io6r5S
Utef1kgkp7dBiGhCMHrpebkGdTirws6JYQi0kgyBgwCFBVVkT4biM/Ky8R0KuF5L
TvV3Wi2MJGkPtb8X3/7QsQtU9q65CfKG27LpW5XmVJ7jrZGTb5ylknrJE1bXSOgo
T5jFP5eeu6+Nqq98k70EV1qA3zC6MGwuV20+PhlwJ960huWIpkz0wbAb5xEKWXH9
r+3a1qNLob0jwbUFkX5Rgo1RwZ1uETvbJOCaJDoSYUKVTUmOv8quuHClGS/nCp8P
cwgalWu4kMmPrXXoZfbaWhGIOiKwwsAtP6WGMKBZ9yUvbJyja3U+k9BrOkOMG4jQ
ETi0dvwKNi5Pw573BDHdQxoANZY0Nm20x99UIDEUORYJs4CoRtFQGjTIS0zFqXS8
paQSPuvKtVnSizi+Iwqwz2V3E9S053FHQAEca1jDTrtYg7TMP8RIeoCdjegAg9JV
TJxPbjaEhWA1/Vmd6Ak5sSB9Ejhy/MJAvpKvngt5TwA8/jwS0QSIaSr4HDbjkxg/
1gFKmdwsm2MaOLe6HS/IR7ufuaRSQe0tRFxPiVyCOmBZxwLb75sbZ7uGtI9/Tqlp
fvPXgSb3006iRGOj4f6WZlDzZ1HhMY0M83nSjC5EE3NDtIJgoGM8J2Qr3l5qIphf
uTa6hHp90dSFgwofA8fKA/GusXeaoMlp13SETjvkebltkYczak0kCN+ANLwINx0Z
V0pnpKpAvJ1Y55Mj9+n8u29d0RQjUr7h9LqsShiLsZcTXhc9h7BPhn+fdsytMEfC
m+OI4Nl7CtCxlmAXeHtpsHQfo5u9WGMWQVDjQzybZdmJc2sFYWBwuuGCAxWHuw/h
5o/PTya2of03m+6mlPBipz6uMKNv6I91ajvMFd1R7AVEYcwEdfigQu+KZRFBMqjJ
GxWUTWcJmOgMN/QIfycSYU4Okilt0ap6EDWBKpPgHMlrCRjPApCut+JCsSAp0pY3
FjY3OCkPcjj9vt2Tb273Ttyn9OVTinP9055hS7p/sJhqo7vy4YpqQ7+MGNkwtZyo
r+ShgZMuVzahKRuGFGy3zo7derdb9pgohyjTF0VkbpDURm0AP4flQCjbnujOjo+I
G8DhGmS9B08L1nssAHBplvI9AeiQfmZvBK54fyf90wIa1dWApwTRDpykIDXwXZsB
Nvp7IjVp/G95IwtDvkzmAs8x+OY1urOUXu+f5YzbK8c6mKonDkczjaM5oLwpLGX1
xfqztnAL1JhUKZDB16aDIIATViewcA13v0K76SFYeSmfwhMct+VQjFv6bOya1GkM
CNZ3HXwrKpUofJrEELHcmeKWonROOf/5naloxdqUTt2BQJ2PaiglMUOEo6pglsqZ
07Q06QXr5MQ2bYr7AU9vrX9rf3BlTaaeOiBhFw34eomM0lobSZFXfQTmM6zpVQKG
ocdoPJnevfFah6Wj1bUg904/yZT0FH1Afup+Wp/8JQsZ+KP0a5jeAw3gHI0YdwQQ
N4ChhMGGvDBG5rVTr3MlgeLvKf5mV+mCE2TrzwEX0oT90s+sgfOnpKRDMHKwhXzZ
9zDqJHSFiTm/s72+mK1DbXdFwzFnBDPuJ7bx8f85fCms/xD6+saFlV0DLGh4+xjM
hwAeP6A2Bhd7lfQ/DwKzsZOZzxCHxHjUD1wuj6/TtXxpKsoxw/phlMamh68fj1Jf
hA3DMnB9UbKvkKOcN4de+Et+3RsBC1KY2+zwnZMA6QBLw9ZcNdZ6V/mpNRneOfly
iYGbD9EdBZTNou122Ooqkdx0wlXRSVBlC60JabiMEIP9MXmW8yuVjndHVB9FZ1Hm
x48dAP3OYqXvEiVWiGq+XbwKfTBc9hZkp0l+k5cEhhqA11r/cstAPqgSOUM7NJjr
GaQ2USZMYR4S7/3fdPs8DCwuvdOBBdkIt0Mvau1ie8JrT5qA98yFribnJuY+09Uo
v8ASqzxrKQl5gWy22hERGPdEtespFUSeisHkOuOXWOrGPBmGcVZitpedxKKSkIzk
CIM7AyqsxkLotXSbZMCG7pyvau0QP81x0eapHbu92kEqUxNcQoj/WKerDZdkx5CD
IVcOKJWFMvLDq0pd5ehZ8CsSo0P49lVF3/DLMvTciIUAiktwejHMwNFd+3lQ9IxA
EPHFLbO3DvhTq0w4FSZj27Q4AoQ0dnYgZqbpiGlpZZfLm1VehYkWGkK8ESmZJnrt
FhGRfVObgZx3tV/AW3IBOdtm4kbzZ7HIEj3F7r5kosQqyXwrgc+tq2HmuO+XRLE2
Q6U42HkJSbbFWh83VKfYuThHdgPKzvQyiKehopfY99S/ZToKMH15bpV6N9uuQVlI
nTtstrufqdEP14IXJ6EZL57NVJ80W5+Sl70+5KikZws8FJRZXOOJnMQdEn29bKnf
8DQSUHaLH3+kRFgxV4h04a/0BxYy+14i4ojNAObsqcnGUh5JL3JxEGFWCzY1wqUU
1TZn3kfTLcZXI4ENX8iC+FYNWS4y/9kzVMyXV+nHtGorP7VLEWypDpffN5KLwXLN
krUIHpVYrsOAes+xic6/h4UUiZEqh8lzDdFunlXgc2PhKZlgFMdV3Wpdo+7lCs1I
vHmxCooJTTF42CXI/73io+2Hvo3djLgYV2Fksu6q9xp53pcyCp8vvfKeDg3KD/SC
eHA8nVQ7Mj+r61Fg4ztXFagZRzZnFMWghL9JziLRT1J+KYf7rWfwHdn7HIYRuE4H
OVa6Bs9t68i6UlZPaOnog/kXa35RJn6dkpYhj8LOoQ/M4Ln79MjsXb4E+Gm0O/pw
IyaW2gyqbs4TVatmpNwQ073O6+nxYKeHMEU2X5qqTOopnOVd3ldsG6l5JIv7g/3z
zXv82MeRAJpPahw2p6ifk3WC1uQ+yJ9YIrmtJ8l9CODc+3zqUWCCNBipdYtFAnV6
gHd1zN0ixE2EmlMJa4GhpLMOYYDUVfCx5iNrRdbW8jgPvFXnk4Zb6Je0JSdXp6hj
1Y0U0hj+1rr7tJQEJhA75enK48On5Kf2sb0gvnn//qCilpyL7jGBtCQs0mFJU0Rp
ddtruUBLlfZ2oNP3F8SdoV8QeMX9ZyzGkRO1AHkkFcgnFCA5s4X/uE2aqNu71yIy
/pLLK4hjEtwwMt9W5U9u+jtSAolNzLmRO1gcjKBxc8Yn7QezDQa+qOn4q9EYdlGQ
ny/jQo1FLd7fqjTzWXTYsncLbduK8Njf+wG3acvsRqmPr75DL84sO3WpPqYtD23N
pQi//v91pCiQML70FC74OqfW1dUtnbNeUYDe4DW00/OC/X/0xQeZokjuGA7ui0LU
Q9uoZ1LK9ODlR4HgMhKWubUlT3WkrdunQ7xmZaNsu1O1p6WBDrEHUsRXsO790epJ
rBuDQnMKLdqNxjWO2ktK2UQd9he6/j9deCMkFRIm6fPqP97Gahmfgpqy0IywaeTE
7sh5Bda8EwiQ1wnbQvXW581N97S0BmaRWDhsUvQaBsx4TlfCgo82xVWDm2B2jPuX
uN5KS+xRihlhcjXf+oQMeCVc4phinV9EsRhodJfF3fBayhTp1LpuTF4Mu+7o42He
uHLEfx2d2r9/UuCsnxvj8/JR7WRm2xgmoQP7g4SbVVP7bTVBSpEZNgjE2M+3l6Nr
OdbUCV0qzvUM9WQi/RCYPWaWmj+W1/+cMm8iz0OnLkxLZ76GnmutZ1iRk1opeKTW
giDMGNRqjA7c321ZwhI+J3rtU0pK/Be35YsgZbMRxw4J21HbzuDQj0jJag9FsWiz
AZIT6Wne85eFsuQgtUVJZg+p4A5XIfinGZWEWD8sqeIwNLRBt1EpAmW5jeEV3hDM
6wVmbOp6PVP0dFmJcJZfbRX+ELfbrDc8d6h1Xdmv4AH92VDhyWIvAqV3r8bRm97Y
2lks5qLZNZrlMZ7gMwRcexT/7zmJLGzQWlQCR5urdeYpYEdp9O15cAbWZCaA3G0B
QlrivtHHrwNNzhFVcSBugMSWTnEk7GwCB3ON2TF86RGx5W0PZyECcn6X6NdtZ3e+
Tdp9BdGvej0a2I0a4T+QKmB/Z9kZcJ1v9+2yknTyQcw7nJS9h5GHnfI4TWFtqJR1
pwlXR/YX9KxLL5T32MRnxZbMOsDm+Mtwa3JR9n6i0bhl/y/Burt41lvov7i4Ho2Z
ijY+puhtnQGsUAnVOxuetYPhs38tNgr8e0ThSPQJcfm2upXlwhTnxgSlltlshS5z
74fk3+UXMRJIO5YMpOrFSBUy3MBvmEH8I01myo6x91+uBSUj4sFBwsy6M8C6iKaF
Tq4a6A4756rZqFMbDccVeSJiG7Rxi4KrBFulSqAO3E4UZHsK5y1S50tjunCMSH10
RJtzlgtoQgh0C2ltccK2rMwVLMvUv6jHiQ5MYp4IZugK68dfreu1S2y+DBTQYI/A
/h7Yu9X+cGITKzSvR/emeVrGpRilDNGFUIzlPa/pErqhQUMvYdb9WoP7J0nKpNh7
lDtKMOHvCZas8w7jO29m6bT8Vsc5SJ3PYqprHlnYnpZ3XcMcdRMki2Le7ObhIBD1
3o/ux2TJWSMV6FCC5z00RIIh5rFzSPWjyU9u7njnrNtvn6LI5roSHBSrExoZSxzy
p7E0kpw2SqT7ucGyZSYczlYE2dII5EBDn1EgLA5qkTcjx+vGN/jLMPoONsQTfRNs
NAgsiXfcGP/h6WjRd51ZH4SoN0l2DntEMTb4fEl3L2QByCHYfB8czaHMGQbQ0ug7
NKRPghjwakqBYPBD/xbASg/yPQVLj4RsswHifD2DyNmS6j/pptp6HWgqREvezq6/
LidSxh9obf0m7uWkBqnfkDSqLSjxdtIchsa/h69OI0T5ZdUgXIf06Z1KZ2saEbIk
MroQr/KLG2HhRrLjwS0+tzCTzKDXDVV8NAo1NsuXZexa8X91YQBFkIS9JfpbCfow
w5SWNXOwt68BmBYQlItR795sYiE/W8ErRLoHslW9q9VVENxUVblteThNuLEwOvP4
CVcah5PpkvYm9brFThnUPqOEpHlv1DvN53CRhEZyyMI+DIXZM3jUtpZXxZLnxkl9
ONDwO6YplWnahcUArpxiluYpzG20oYjWp20aj+ljAVS666J7CCMSkU+mFJ4uPXjU
31yHt2wHpkO+qbyvl3BouEuJ6SYlBJDdy22cJXXsOZaPG5zTKpeMWVDuu0Fc3v3g
/2vAVWdcqizxKO6WenSxbHWYC5WJvAusGk35lpdYVjAOhsRBno8Ej2kSb5FrnSTR
krj14Z1jqIJgprSe4TzVyJwboy6jw8n+lp5xX2khSbnhiOAxVP1IBX7CRdjQVXN1
+HZLwrHcwRDGuII1VwqmqUq4LYAEVOB7+r3C39aKkKhk1b/B1z+4SF+fjBEvG7AK
M/kWBBCPjlvj8CeoJMaiFzfjSLH+pb0DjKkNOfvRu+Be1TGTYLvL/LzuNCZ/GMdp
+6Si43eepVbjZe2ffOHLtOpFdxKdyhmNZtzl5lhe+hAZsnhJnqA85SKtfDJXBUyU
MKaWSE5ZErXMmgoyOqit5PfEFqVEbV0PDPOmUgSWlo8S/C87IJ+Y3Ou70zoe5jOE
OrolxQ6Jrnu203T7FiEETA/0BTIjyb/epiV+Ze3X9EyVvSXsTPIXUb2kDoZs8K70
UdVOb3IVZMDeViR/J1g2ooMAqnVRqATA/DHVpdisG0NBiHPd81lL/yEUhuuaquhn
8xceSF1kAtM6v1HUJ/7pGm5fnFRxUXgQY4nY+oMAJ7VoQP9WlA+0l67qOZR6zFak
kcwRnAjGYfNkmXPJpyoj5uAsJwA54e3FIwl9wSGn+QIy9ZH2tnsMEC9BWeuGoL/Y
UN0ti5/oSusoYTvpJZ8dW7JdTsO2EeU/qVE71m7vT9evKVU8bl0tj2W1nskWAVfT
5W1B48PyXNyt0WOqlnwUQyAKgH501VZDd4jGa9KsBpo1tA9CzTl+RukNUUvKW4a0
N22Ep4NLrIk/mTjxrVwqCCzVxKfZGHL2zYXw3vOO5YQ3r8PPU7Ssit2raGLY72/d
JPIRRKv5DtpeZ+RqrMB5zWxSdEJlcJYyXJn00qhRINQtePeHN7S7s2pF1rm3S4+5
P44M7nCivRAYCOb6CxWw/2jB1VCo7hSTx1PaEdxGXTKVCexqwsgugv52hypEK9WB
hdclwoOULpcn/9Ui5zUDB9G5oHvkW9/wJ1FD60YXCcscg2l0HGCj1rV7Mn/xg1de
RxUTK5dYdvBUe5sBeiMYGMVg1+tU3q6lE2FQvUBTe2aFrnGleNejJBEJbOQdPyxT
d1tqndG19F5G8cc5OuYiEZNibmKMVkkf1hr+hGWUMO+5zQXKW00LaJHZwVffU+fx
GZaVIZ2ul9DleRiQRIGURTARuVGQg6F7j1Dq7O2yy/oY9+gsm7dBolLTm7/ABizs
SE48sxl8upFyLw0e56UmzffwrkySK4/LH5DUEzTi2Iq4Im4GejuXGdhxzLJ92zx6
EuSUa/EK3A3khOtr5IzPi500jyYvnHojDMv9zZYnjYIgQz3HHsAQmukDSUl81tag
f4OFRD1rAh4M+Couz0Nv08cakVYTXdO9oDZ0MoA0wL/s6Z9JJguZxqflW/XcF24J
8V/ZICfEs2b5m2XEE9pgGLTboLHwTvhI6DNGm0CjdbXrWqSVPmhBXnXNG9seceR4
IJkGEFVOL3ipfZy3QFwSziTnkPJpPLOM+NfxRTpU634M8Eq0O9vjSoCDpPQDon0J
3wq1vkNNiXkeiyEFD9hqaS7eVFBsg7ykIGmDKCw4vVwUzXyZu77j5qltFedC8Rm4
ZNHl0ySnT4dA5oAQeJejHPVX8oYWjpOmCBBy11/TdHaMyqzQTuAPPV5nQCRoU13P
NlaNt42MQTJzSwDaKVIorBouaxUIFKRZay3JrH/o1MhVOvQ33qcvBR8tEi1G2bdf
1exI6iqGWKjal6+QAECVo33CuwYd4rtuMEEAp2BQ8lSH2JMhIuqWTbtnCupd2BK4
DCeM+Wc99f40yTXFzK7ICKdlMssIa8Lh9g+fDoq6Gx3DhfJefZ4ZRtAci2iTBNbm
GvkFjEgmfxvgf2JK5nbH1E65OBOJurR8Iffj4Ipi4+RP0rYEO2augXDlIrx4GSWB
cYIpmjkgU6BInja6T8LVXB6SHrqDL9SN7RM0Jez83O2tXXQiI/MY/3opVbrnpoQ9
9cwSUysbkbLoC9WIEsPZJ99toqBfGNPZX/4S026GYvcs4RhrGzf6WqJ50aErKZYe
BpQwVXkGGvWTO+ihTFr+Gl6gnqfM8tX3sYRsly8uv/ZIMLEkpEDQzDRMa1Yh62Za
lIlFBXmSctsHDF2s9tYTcdhnCaViGTGOxlN+o9UcNz/6D+CMFiOmFEtfMEw8FMwU
uhbnApgNm/AKSDPHpNLYb/kkd520sjOQcKelzJ7cKKwsWI+iCBJWLWlxMvAdKwXh
q9Mo8uaas9Cz+0JiX+R7g+k3vl/+8AcmgHPsWx028JjgJve9s5GZWt/erFEJqym1
92WIUC6L6acDRugdXt2F1ej1acwdtt2CA5x31Xu4KL491WWH0FGCXdgbn9M2G4+k
IkJ0DigvJ3ErRxiqnuGb4CzBTQYXqA3eBF3lHHXL4kv3RNKH2S/rDLATL1XSanZG
1uddZsa+7UCT6rfJhcJ4AlxzV9+GGoI91jOqVqLY5kijcbj/rKI4ifxxgIOZp9Sr
+U9SQAPAMcpbj0lNx5XnWUeUQjngF3+ucFw6y59rYMUoGoD0gKFDGCFxQkk3mO3q
nI3Ina39icDKnhS/86yLAF/Vkc6xOSxXxX+pRHSQu+esl8hbkEgW9NrHt+/zkSCu
F0GTm8hsCvEuw6mF6htuvqdHIECoNiJJz3jWcqkbrgzPRb8tHpnHne95U2Z635Nn
EW603i6iV6foXXFPtZfILmyniJAw/JWqYWzJ72F7ovEAvYpociQi9QcTVFRsu6JL
N862ZKinSJeg6c5TxbtzKeyKeen5JiyLKJx40CdIYVV9rt9fvkpwj05OUlsUyrWe
DF0GiHeXxlDuQaCWdv0jHdno3Vj3HVCunoioPFVanA3Xrx1mIUG1pmzRS5uAhqHA
uk3m0wSEgctOk10Hnbs85b/zmqQApN+5fYrX36N+0diGJX6FKvi70boSgG8CbUdf
QkxgWpUUCuNqDR3CKz+nY2Quw7VKTJUKYosRRyZfdtwMnj8yN3JeVKPnvqidi1tI
fW2M4tTPqR8egE82OOQmilNHgGx0vETtXQF4HlCf9fW2lcY3a+YRkegfQIi/2DJa
HqFn0dgg1Ktnox5ikmvM0w3O9U3qJM48Z3Ry+AU4PHDBcJWaYj2apyIEzPkahz/K
3+AptR8HWwV/95ptW+ZTihj5iTP2EHcHBmSCrT1biolokp6qAgSd8y1oYfpDSWzm
H1sTFbaH8/xF39VTX91IjOZIFE7b+j+jlZGNhEwEPikxrmuAy9Dm9rqoCNRg8a9T
62TCQY3De3xDexXutUk8JIfjlLM/pKRDS4Y0VF0avmiG2gvgCAbv044TGl+dfCDb
9S4rYyJ0/9GakRZPUTSwhB+BcLAGZjPl3clNUiaPwyVKt1xDmqEBDzHhjpcDfhDn
jBJ4Kd2L7AJKGM04xoMlSUcDGTmPnGAluXwgyDDn+5dfv967XMi5QIosKYJ0s8dG
Nc+tNL1ikcnfeMOitnO6+0PQy9BfTNCpgZJ4EWJdwCRiQrLAeB7d9w5GV99ia0JU
f8It/GSlrEDEuwRzlPZjWXcZRXLWsgwkYZs2K0mFoUttuAFDZ5LBD7njcWeyWvSY
A/zYYFwHQx8zhN36ItFTPsPPaB2JQAe/l4WHGJoXkSu38KgRQRmjsS1Nued0dWaQ
/H20hmteBnqanN2+NaFt76jOCRPSr8ecjkqL+Hy7MEC+MSWcz6SI0kzn0q0MRV2/
eL/Qpd17JpYNNyx1R1yrvV8d5zbZHtlmuqE/8/WTqel6Vn3BJiBE5ef0z6aUKTfz
dwmkqX81IYXqPMSynnkoC/rgjjz4sQReFUfCty0UfnleD/stNb52wumZcod8RU0S
ear3zMYpRoOiMTFXFsVDf7/PyUhymJfX9nR3/GNO1PxZJ3uuApH1sbBN7RMavQIm
d9vzehnrtBJPHSl0OT/10ZCCmZ1HFAUAGuiLkMiU93zQiShT+w4k/EPVaHePUV6s
uFfUoUqqX4GTfIRBLiPuLQa2VsXM3d1BVkH5dMcy007THQc+s1asZI1u2yHdPUcb
wqlaN38ioW5BFwpARw2wGw0yYtbNlBtRvfAZJTyjHAZcUuX9+XJFIwLD2R8ECwFx
er7BTOJh2e4kQ06FMIly+R7yC3Vcq7DcUNrag1MFUZVZR77LucOmt4xTHJWzFRTc
Co09thYPfgxjWNwzxooa6SuPN5utiSe1fEukeRmKcYxx6nqAi1xOkO4S77IydZTh
COqQvvAk3+A/MQ/CuioB9TnGvt1+WOUhyh3YzescodH9hsiDZH9FNEsJYk6VrmBh
Mp0fm5MUapVExtjC+owEUrHuh+3bdsnsimKA9hhy89bBspS5kIe4tWVRa2Qlb3L0
BfGPAz/MjNMLQEUyLDqckc8EZ81SnZ50/OMCjYHv0t1A+HULFM8/TRog+tm+Ee2D
m4fxgcvvBeo+Wtw0L1U6WFf5VpzWEaLHJ9hHi1B7RgVvW8OPzq0IXA45R2fsbAcO
wWMal3Lzn8GKseQTmBkIaVg4hZEiDK9KJD0oKFuv907V2pj4f9G55l2DjrTE1eBu
HQYJPgwxsr27MC2N1PrBA/pY21VzzpEVjPLMlqN/+BI8opsfk0Q4zUaIJWfXdxi7
qqT2Vi3xtXhdRp1K8Ac6nOFveK9MW+jF11tDjOqWdtK4ulX+ynEiSRwx5MJYNJjM
wIfKg4llTZ9yb/EqicW0PJ7CIA0/dNFH3LrLjwUlj5Gd8J/43n0AmxuA+vSCltFa
KvwmI8bkfnoyxyU59CYxVElAP5+1ZiDIxQo8T2/tYYO00mon+z30X4UakQmGzGUQ
SS/r5Tfo4ng7kogXpZbZK1RdqfZNuJnhRwr0jzFxPrL6oflchjl34IGqWzaf5Qg0
c/koVk+ROU+BfEWmLSpt4tRYlpLas1Y7LvA7LMIFRkF7pQpTKovB6NBD3fSNaKEV
vVuYRyu53QJBxIwpL4AR10xNM01TFNP9PPG06mEjWAHUzNbUPSdupkraHcYpzYOr
kbM10G19/RJKfr5xP4ig61PAFeKLVeIFGY1njmdxTHaC2fA6m1yCY22gK1ximARR
8Ar+NtTJRVeww+PqEUcRXwBAZhH4xhCO6LMtdKaCbfRBnDyctIyNiB6bYL7kGkX0
7BR/E72r886rPaaHRvQmddln6pvqmbyVvi2vvfKyjNB6pM7/yXQU89VRUl2hwq4P
cqnm0UtxUAVjcdLWauJJpeUaQGIqG6MjBv//D77pDRsqULQApuNz3mtxExNEOmrr
3vRAHOgXzKzUuacQ/mWBbujp33OBbiQH1W1j8E7VEmdWSo7XaQUvCs9oF6AH2XSB
Ef01Q0W15NhkGMQI+a/VEm4nnG/Ae6pGHuFSzeLVz+TwvW4bXqS9mmOA42QW7ud/
d5i2/SCch9PZYBtEZOQf3xz4aR7aWdMcN3hEn7JX4uDGWLcftIng0FxoPTJLKbS/
7sfRyv5J1mw8uXhriYcpx1Ms+Smr5GghXpWHhl6bPK2w3GHmKP3OHrhxDnEic4zp
W1xuLbe8odbB0ETx+/X6PLAlEzowOXOrvcHL29SbpqFRCPv8/qkFpvlMwOD417Cd
m9EkXiex2JPKz0RbxmlWSXdQMYSHSw8aP56/wGwwi44SPvJc3Qg/153g8Deyb9x5
e7tMMeeuPdfBnofQYrkauDvkAW5w9pnTB5KbXgk1yzIUGPGW9E60cNEm+tFPrZu0
ktjrk6QO2n473yPBY2URjC0XLCdxDZYr15hKV0GChe6mRiPvata5HfSjO947SNxE
zA9QKm0PMqlGVlhrMzUQoOmyesOpOEsxOkpU77iQrgIPGnOnKHUeZoN1OIKyS1d9
Z+4q+sKB5X9rnOze/H7Q4ZmZIgosalBoGIFr8staeP5Owtlzh0UAipEjZppklAvr
53u/ImHirFM/HZ5F1FbTjuxXfHgvxbTIlV3WVpr4bsNVJiRmTuv60DUGfUhC2KrD
w5LRi+IGQki2nJk9ACmpjIU3FnzI4KIHRW2axq4SFnfACMsu4bX9cgYqIr26nE1S
W6uXyeR0SiHrobEKvfMLJtHzsu8afaVyYVFM5WB2fOudrBha9zBq//z/TY5wZAwI
Rt8OGXD/K/ys04NY81OegFjrzlVEQR3LrVHjs6d6O9F/Sytam0YDtgJQR7swpNcv
W+e5qJoryIpVj1gyt7L4PGulUxRPuCjYs2fmviSdZSLxKpm9uoBH9RJP5S6amgmJ
zpr5jxPFnamzs2EyjtTLgUYLBFyOPyVFcpqrZDFujpbUcGNj+JglXVBafd9vykxP
NZuXLDGtZbKt/tMMM2WRNPT0HxSY4bIamocpwYC1JozuOKsL5zn4t6quvOAF7KgW
rJCcwRVB3I9Gcz7VHSTzgFuBqpWSdd2PpMtqgsm4kxrWUUziP4FxmBI/W5d4Im6Y
JD/QadHLbI9YZ7khrJMClYRN8z+rS3enMuHFO7+aqAR+rrcsxAqoJE4SZtZqSvad
hX6bgSH0cckMB6uCuMe+JOZ7T7vSJvqzKtuUB3vMhRyJBsRsLwQBIfoeuynyS97A
GNhbvdwSqIyw8Fj5KNbG+q8CMq30DSb0GXfSfIfz3xHQPM6K8oWV/GFlXCfN4wqk
gDy3+/DX7BMVVHIVQMvdv1N8EzbNKyq3lM/P6bLrrW4K8Bz6LQ9PiS9HOTf0PLxI
MEZ/J/h9VghW+Vsn3PtpgeKfaZ1Kz/9/ufSK0Jew2ihf99jua7mT3WP88VMrC3+p
gMy2KPyGxK6kTzNCx1gHNQW1VWwr/6WAZlSSIC+y9KeH0thZ+90xiNdrNerSHb+L
LvvjRrpbce5xJnbh5fPwd2qMw4OQzzey5fQHQDsjHJwX+BtatAvtD357xFVeoRvD
v9SxGDNG7UNV1yLksqDhe60yy501wOxuJNs/5ssoLzuRQeiiWcSgU08q2SXM39bN
q721Sa3EGiP5xLLaDg0uzSgnyY1mJzeZv2tm+8onw5B+CJuZtiZ/jeLKGap8pDsj
fM0ueJiEY8PhGZ01N0rRKi3tn1n4m1HI6pGzEYN+LIfliYxuTAmaoJqPLic+dj/3
hW7vshBaoLID4e5VmVPopLJOannWfuAOP5XU2f/ruiS5H57f9bTg4VnfTbmdpcSc
FO1tIm3rTjUyXY9gy/YwU6tEXDnEkcLHyEFRpEkWfXEEr7/rpRgZmJ8NaHujgirc
unecsTG7M0uAcpMulGqRoMDccq5/RlM9aR+X1D7CPpqSu5x5sMxt7GECdZUsxWEz
+avwpYR/1HV4FxzvnQF7wYMJ1Vg9YNW8++xkoANWUBhXjsbH7nBXwnYerUt8j/Jr
wUnEzGaSM0lx2Jymbt775JYHlLqgGPbYeWsROM6ZwudXo6YKDsvJFfXM5NUiPGHn
3u65xoEfSFNqfyPjHCPCrLpTg+6fiwVxJGtt/OPqb+iaxJmaJXS1LKRNXGG01/2+
cymCy/kZ+dVSQEgolkvSiEyFVN8DDlEMGSSs5L+N4qTNPcyiwotepUsGXlEmzJtG
pDyQ4md24wZ/XJEH7heEgpfG38hIajQLs3lKIRB6GpPEZpKVundQLokSWju67kC+
eV3g6e1kGDi3gdt5Xx56Bm5FHe1IL5pBOSmi8bzosMcOKL+a4wwjprn95JVE6nly
/2NQd05I8/sAZiFpqd4Xy2+rv6oSOOXlWYChL6KtTA6ASOcvtaB2s8rMx3bX6CX+
ek0aOeNobyeNM9OZATl+22U71FHWFS+KVgzwux0xDz1hccVlSy0+UlyP5NBjG6sT
VBPVvHiPRDnnto3ZkTDufKXp2tkGki6aRqqzCP4qYIxZ8IQyYN9PUaEWk4gyv/Eg
8eBCZd+JCRdGypYXgunS2L1sv/iTDwhtEL6/oKsZlauOm8bXyb7b2CLqhCtYcmLj
FjuEf8bYc4TTHebj/i484jte8trAGQ56FQ9eLZskq8a2eb3uc/lMja0oGtGP32sX
sSY6rCElGngOvEKQVEmvSbI55V1Ozn3RtZuo4HY/Nt95j6AcyQB7tzrxIqVBvQG3
9L8nwZXIbMyUlcQdiAIhjYcRRjZdyF2+k4SDD4dwfjBWhUufXLr1/RUnqKqvBHLc
EApiNJKkyTRh8C0zY/73aNNokDbayX+BQQnsXtqC93T2PTwS5FiZ3g0cexK3tTl9
ihMfBExv5d+S46cxefYqrebjdbxHGVeva8LRtNbKZko02MIGyg0TwLlGKf+Mx9G+
2IUTXY395EPpal0+T2tOvdwEKakQQcUcutA7MYPfYBnIQlmJy+iSABzCwQYRTsL8
9WTXmgZvFL3n4/OxkVQOKIL7grVdDbEvONtKXTC03nzCoXwCZfx3YteQZpS4somS
6Gzw8eRHV25q9epby4QXZEVKaFbjT40js0wnHOz36ncu/AaGCK2YygY3QUDldH7m
uPauqa9WXYVfLciBKbj2gddeuvFqPfKXQyb12G8CoBW+7RbqAo5p8SywnCxTiyZA
2yVKrT0iP/d4B0s8/Rp9R62XuDYSDJ2SmmEjG/KtROs325CfutkchfYymbWZUWt3
llb3alXsLIWwbB39lyVCJb4byoiEtKqaWhGJYqIdXAvk1/mFapl+hYSjvvkrULvR
0nh8hes7UxSZMVNFOFynCw/24StEDCTIVTzdr5RIL09IFwFle/UODdrVKYe54YQC
5mXTE7DW2iTdOd+M2hOfjrCVacytzyOcIWdgj0vJbTtTkuHJ0tk2/h29nTV3jc4C
joRKy+JbfQYNQQRgB9dhiZyTRHWhsqP6Hmk5VZzqnA9hL7R5NDPXBt1IlRfczAoG
NfWg0sAq5pICdWcm2Jnv0fi7YB5egyup8ChFKsGkrAhPk1R+0pLiQXbkGwX6xG5v
F/1ldlZgm9krvLeu3CA3Mp/Pcg4u8/9GHW6iuvpbdomhLGSW/7yXIaqJCtESES4u
7B9mYzQmxysirZc59ItiFdUK6ZyTf/FE/KEqt7kIRRU30U9FLKswmU6lbq1wmjfO
gS+UarJb45tc9vmpQHWKXE4gCJ7Ba52e5DcxAeNBvKLdvLikt2xtlr2+h3sDv5t1
l5uiw/+OB3FJ+hmD/B1CPkJdriXfwYobPzkeiFWNJfWiD4ioc9Ay/XEiwqJJZD2X
TkQ9EVuekR4423IATrXkWiw93X24tVaTKhQXm7FHvSnNMjW8Fx8b3ram656Jv7Ue
bOcYNd5qZT3bkQ8JCYPK/Gn6/uYSn9frYs4aC2pmCqWDeZVk5oRXOhSRrQEgMOPV
Qtc5vyRnX4X5rijE/ydlxX+/6fKeTl+VmPRFxQi72EAZndHws4b1Z4q6agwzlJKz
BQttRkbaI+VfGcQMQHpK4oot8e/p7y3Q1EMAXQLfW9Zb87ztGhwxlaDPErKnXDNY
KPvmXs6UZyXmnQpSgvsqUtm9eCWF8amPrDT28FT3YadaE48mLeK6T7F4KXKIkdNg
uJT6C4lKx7WLqPmBgkKh13wBA59lwogpEvC2w3Gcmu0uIiiFIQzwn5VVkzRQ/6AO
h+GqT4aKs2sB6oCzS3k2n7yLsV5XuJNan3U5c8jrpyORBN5u5lp6xmeXbl06YiZy
k+LVi+Tqhk6xurRo8buMGSK2lr6PCh7PcPxXVb8Oc67OSRa7yvTamEw9NYT/USg9
HyAFtXR+qFI0crOU7xR589kOVTuFzMz9xtI9dUd70QBlqteM6z/42gmKY71BZchY
VDVXeyOTOEdqGmfmhEY9pghCQB00wk9uiqyUYwSE4P/v9Q3kZ/IP/NrP6wS7dGvu
+N2vR9JvZW/N+Fu2WV+jxt5vET/EjmFQLX1IBj1jXy6H0zJ76tbqV9enrPky0WJn
7mbJd9xaGOfT66LRPsAyJBf6PEN5zm9krK0qdTVhPmR3zhEzbowOJ1BOZt4jx4en
8BFwvRf+F9X/d/hkj5yrQhwk5P7jWckXmfL/oL/UPCRLQ2YyFvbEdMVVaQ73Ez2S
svOo7RXsXM6dEJA6GA/b2WOaDRje5SHPaBdIbstdR+S7rICsKH+61s5X4/ea4f7U
giBbqeJbV1kRK2NCD+taC+oH8LPAE18SNHe109uRF2w1IN7GuqPIYf5pJ4F+fC+G
NVNQZjPhGGaTPxePvj5UjIVj/DXqNJ0QmdlvE5jRwiQ8I7eG2+SYyUlqwBmnb7fC
LHyLqVBG3kxEo3uCi7D7RiaU3GxukRFaek1Pdtse8CfEhzBz+ajGDKo7kCgn0wvY
m4iphIh7FVBk3QL2Dn0kxWu0j8bdDoUBW3NORkBFeV+C57jDR1wf2VHb89M+ZF58
ifnhJlSDXKtjfKZyde/UeelC/Xnu0hTsBYQiqt9tiA2+kOFYARZD/jRvwhh/bKZg
NyojqO+0FgjFnlOKd6Mga+nw6jYn8rbfaGj4kV7s2nPkxFwjr1JX2o5QvJWFpieI
9C3CSvb7q7K4WyCOqL8TPBm6gMJPK9JqBVCfB6IYfMAPfKSVEqNm2CEqzR4NObi5
ZWKCNrhLTZyCLRwQeRUkrY+Lex7tw9LwcPJhgjpNfNFPGzeOPdh68X5hsYjMLoGa
XaL87cMweDTYmvz+1lWJn5Xy4WrBDi37IPYEI+W3ohWZYFHznIgnrdgHOXPR4ePx
iFMrNyJ+tjphxGKwZ6ksD0g5G262rAIYtaIM4/ZE+hfwGewtTlEqM0HtpSwk+eyB
klYdH+Fn+1CIv7VBLG6c3ztWJPVkpn1NiBTVrGAvYnD1z6ttXYqmTVJBkcofowgw
+iaSOG6EFD6LKxxbRR9xJPBwmohP1S3JcDW480gPiGn843vmYcsci+B5cqlW+J1v
vGDK24Qsw0bfsqu3VzYpFmyv8cVQjqumjql6NWzuEqlK5hakFRTg0WAwUzQoIliN
mEl0Sn5iAKM3JoxnRs3Hgc4KqGa8A70nsgldHxdCz11ltwJaS+3db06jjo3udLKS
C+fW2PptKpG8i5QvamDIzcN7cdJGaLc+boHGWP4yOA7saf8m5SgsUwBCL2HN2qNp
40pDV8W355j23Xy+iaX7Qupe6wSwBj6bbvhwJQjjJxxLNqNC28V1H/pVOq0w4q7Y
eppWahZK3AvwqnVmFehBEMaPG8GlDj8eYEagzOcFy6B5zPvfP2RwweLDjL7bKc2T
6lnPRr+hFyyKDushqZWP7L3SqQnm0bsnCtDgHTqElxbaz1m6xAcHNZ8zJTfy36ei
AlsB1d81K4nTfTKIGEL5JD/jvMxvdXvx2hovJ5lLG9fz91Oyg/+k0Tx7ajjPtbHM
s9A81DnhOS++J9sq9axg1tfIRIQpk+XUBbXiJc1NaNw93CudAR1VSe6bcbfoLj7i
EEAJQSZTKjmBJCroYdkbewzIAkot0Mk4rtURR6/MpXOgYklSCQOF2R1d5mxvrlVh
P9PXMVPQljNt6w0HqbsOuqYcZcLV3F5ip3E4Bwo0t26EXvCYrz+Pbu63z90FWzt0
YhWfcnjzRoTALldRNNG55SGLG7oOB5kRpJIrCrVPQ6zLcx/70YtLO8rEdE1sQgsl
jGSCINDY9UzAOO8N6IHbh8hsZdRwiHi7XiuOV25FRKDAUeQ4nbwsh2BCx8cFZSia
2lMKps7bx66fmkjmhszhCNfpv+m9+F/Ts8cwDdTPy0JmV6a2MVUkl4cWS0uLY2CX
YrHITPoB1wHSm2UG1q7sSQ9uzFZn3V7XscpiWrlznjZ2tzSAxjd9r7wIqmlZmVee
C2UQdwNBTLyxcjStkwN3437qqITKvgFnQ7M81IbsSCi3xaf7Ww3sHV83fMFO1sf2
H18iedliiwpqXRNlkOVa16Bc2wY/nnQmYhgVY8/RR5cxUG5Jj8c8ntGjYgkZd9T5
QD+Vjnd0TxpFFii3I4abs9H5n3Y8ZFRDUlmpnKVXRWyJkYbPZ8zey442exUr5dgx
CLMxeuXg43srNf04M/mUbunNNFO2JrZSxi1M+ahjHYC5Bo/XxWCIXL1QR7KBSPIA
x3eOsUJw34crMPg+AxJhvg3LJXVRsEWogdqHEln7c1QIXsjzZBfai3cVXc0UPHmN
iA+TkW5R5MgoGGY3DlVemuChLwWmB7bjYRtURpZoUHOj5I4yfmoVGk3113tec5Iv
6Ruj88R8dyN55n+1UGg4kCOqpXEslB6kxsimCIEM4YmPbyHYdbWOAvy9XDbb1Wy9
2LEs+uE55JbVcrCyrYwwPx0BtZ4yCpgTSPu0UrQ8As4R0AmwoCBYmBRlMyNrhAZu
hX86MRJNlmj60gYEkUPMzGETUBr90bpKCF0DjIxLL1jFO5E0tpZ8Icv2LTj0Tvxf
y5l6turZyjC5+m499K6Sluwtdb6jIbSGCZVZphAmkIe52pVdGDcHPeItmF/6gslN
n67YVKtv0vQL7vrIW38A2+YdoQe0/Yx8so/EIMNfJnr2bfq170+s+DwgAjXbKSqE
91FVwn+h52p+lNQvhDmcgdNVAUSMO0os6xCIv9NblevLKVDwAblV/Nyxk3pxD0B6
kTKDKZJcpqDAWO97rXozGwCBJB3gcMgRPbGuDKH3Y2jn8JShS9eHX6OHuLsVQUBu
lhIPzon/YW3hnSZTJYCZIDaDs9lSRnq2j62/KRzJ7M4iCoGMqiscvp8CJI6xrlse
AeyeNEeJ2uRLPP+CMUKno+L8COWuaVNr0fjt+0lArkYc/a6nd1FrhUe0amLdf6Ce
CYzc3P0FcZBtkIvKN4SwMMEb7C+7hNr49ZZF4QyWOdpTk/gAcoyKneotKd0FXlZZ
e5RE8bx6UP/dDhr+lS1WPcrgozeK01B3PpQYtA8NcDfsKzvDRx0eZyuTUDDRhurp
xhTsT88Vwjt2KPzWSc1QgUkKEz7WmM68WRZixcMdSkGjtZxjIuG8uJ9KXw+ERvoR
drVaw+Vi2gnoKO7M6bOgmKGUaDFydyyyF54X8c9MxfQ6Jjdj+cOW0CIXCWUzkz7b
oXdus4Earh78sVQS6prAw/megzDZoAqKVZs0Me7V/Pb8rt7fx7RyKVGrmSM3Fpbs
mqlhnIxrwX+Xm6zNOta6K9mIV6HLXwsIrbf6b1ydFxCpY8cU0WYKPpogeFj/UUIc
pbckRTf72hagoIEVpRwJsR068KFjnreHEMLHu6DbC0YVAt7dFOcwUMz7X3+th0Qk
XpDXyePwYRbgYaTpg6JPCwZ+hd+Q4H7Xcsxx0TNHdxe4L801zEqX2NCyFBoPwuO+
yg+6EZRTO5AtJw/zTQ4eEkbownOKwqyTw90YdZTZ7RNoF5LBT6BbP6XvYCZNqMB0
i1pmYYIgQq21abRjGWTLlKnfgnz5z+MvbKW8GYs3pe3h3tcFO9FDcncGtf0/duXJ
WBI8BRiU/7bMmzFnyiMrMf62O9X6S2YWbPm4+Ux1XJ0Z115W5DwYhhL35KlHLX3r
6FO96jveNeads4EHR14Q5hdNhv9Mm6tZ6wXWDhvLh7QYXk0lz5fwS3v9Mm692Gup
zRiAiYncDDDGEO8yMRnBJh+maqcDw2F5rFw4SOgLZEhUo26Vu1wneVDsP1wE64JZ
2c9J9RRoHCjj5ZN9dwG38WheC1Z4KFo+JPZyaBZzeShlnCmwpRr9/6ooLyuqlVfx
mFO2nL0dQmqI+jBNE0GqxZ3E5KWditoCAW7td/tSFcxBaYRE/EFghkWm7MiESoOv
7Ks0bDwDF93FfwUq+hWmDwgRVXBtn6JkSiV5oG/InniGyR/SVZf5rW8QElODVRxV
XAI/eZ6X+PdraX0IQltkhoV8aT7CFbNXzmSg6LhkZthXABZ+fBsG7uDQuLIJIQUG
8cBiYJPjFhK3ioAhHA/UPSkrsOgtf1cYFun2B0qVnMVkTEPPzmmBCFKNfrk0Qt4N
950v1ZPOlipSofxL6ZfKARomgrBWZNizdijD3F4eFXjAT6cBPt75prTsPpchkjpq
6Yiu+9GB/0OIMHfQETiClKfVX1ll3q41PyJp9oafVxN6vB5gqnKGyHIWLTyZjr3a
u4kwnkNC+3o3vTW++DaWkS+85TMmVXAisRl0Aio2sK/vIJL2Zq9fp1wuKz3J+fAx
Nh9Se8CTr4so0QicK4U694QDa1S90pdqe9VH/Qa/JBjdx5w5n5p+M/9/c2KjEm8o
kdzUDlws4X9sLMfUDhDVsGHLc1rVVB5ZDiqmUYbGMQVFLlcsoy3yX4vqpXdFupiV
BX5mzLkiOpSnyNzZLNIjtETztQwSa6sCA06vyKvvVAejJNCmaeBnSigfnwFfYc+Z
v8sCUvbLJA6c/9rR9LE4FOoU6Pwu5ZxQ7OLPDThg5gWwfeOAOXVNNZIUmwHDevjt
OUqXxPNdb0Sj1GzL4QBcIGXbtm0BC9LB7ByaO6Xc/WOCgyWD4u4O2pZwcLvj9IKv
jS78dl6NdrE5+RaESR7NaAw/Efucf+V6CGixhLpM2ewmx4a0W0gYrl7+RPg8JH/b
utgZ4WyVjM80OsKVWuiBcB5zmHU/fOYMSPoC3hl4LcbSlqcVWgb5CG43apgU7LZO
0S1NVDYoRee3qtmRrej2IRnfvpP62pJGD5NRmUDjsgsdJv+WU/gGRBvXr8rrTgH+
zQRV1ORcENRQuBUGm2szBYr8kL5FPgCPw7FAKA2NalllXpre/k34iZHGsap5E4dT
dXEhP3YTFjsYo+5PjmKjC9I5C9jkzUT9OW99U1jSLaZ3V5LrvbhcPF1iAIXAsBMo
806DreiuJN+xSoSTgHIW3sURBNuypUS9KAuoXA67fGftUbXvry+WbJ6ZiqTqGSkP
pURkQNsOMZVZ7/8WBFQ5eDClSAdkRAH5+j+5i5GTGvzznWfOmTi+Stpo71LsNAxw
hndFTRrbRONDpMTS0OpiAa7VZqfcv16jphH4Du+8Of5A7w2Lfim6QUEcUheX4ddr
YXZcI6PjkKJrRFgEh1i58Ggh5K1DbcTxWn4AimV9K2eZYNMB9g1+FGREUTYicVRh
qzQ8O7KZuHrLS9g7MiCiBjDzMXk5f1DQODLUopVo3gou2gDBP5vL54dERIAlp+l3
dEY4z/8JRjagFkjDcKlZ7OWQoC2XrSvYeaiqpVdW9LilQyLgTnjoMJjejzlftdBf
OlujSrE3AHp6xD/JdzBZ8HPYYtGaSIub+VoCFcwvOPRvRKs55Tm4MZltzzQ4YPxa
92SZRTGGFSzFVes/e+kElFW9ypA7rmldKnsAPYfBZsRQW8uVH6K4fzDXEIx3pu2A
7yIs8pKwgmcc/8rvxCUcGmr5H35hSL84VbW5kdJJP22f9vhrPK0EuWVJznavzOBj
S9E0F8Y36U42/cb9vvzohCSxrTdrAvdWdRbalLTPIVt0cPnVVUlv7dTzg+4ZiWci
Alh0ZnLk5uU9tx2Cn89t3tD4rKM0OBMSMab56eHaUw5/rB30vJpJnSB6vvsDimgm
H9yX+Eqyao0xW0//htbT9JIRZ4Ik4J071vTJCQ8ZxyL2XYECK3JU31eAPlAx5TvA
yXt+u8sRQQySv3BsXyIkaqlK+kivBBni7fBPioyDuKSvxuDH/YD2f6xIou2/v9RU
usO+7y7Rdh+s+m7FeUzlYJahQua1uBlbOpoAHAVjjdlo6F8X0FaP9oynJTZgMUVx
Ru3kmXkpd3dqal2KdNTQu5WKz/f83jStQ5gw+hTLSAVijLCtKTo31YDCjQUHq45a
8USgx2K8CyZ765WRlgRIR70AdIquBgHyNp06r1/wZfDm0RAiCqdCeLvdUjpXhfEW
tOc9j7IrqvFq4MhbYLubLmVB7UNxTMFapKI46xaP+2FMz+W+SnYIQNLMGLQP/qlJ
zD8hVrJ8U574Jl+ZhJsJLdLITJ2ouspmivfXRx6IJjJye9MYojItt4omLUQgtFu9
pKwU/irUcSAuIu+WDtaTWf3UmW7BnAg+8CbPv9uY4l7tDqnHZkbxDWXmGvWIaXtd
93gJ1los2+yItIw+qQp41obA7Egh0+yH+JRAgc9QCQMthZjBbFsvKa2xd2yvI4Vu
W3fztdurn4zcF8J8Ub59QjQ9HLWqOiJbqP64rJ7JvR7v6DS2cvIFFLWylY17QpDs
hdap1iWWQyPofLkoJ07PWnP8CzqgAmPvcCgTjQ5I8/IdChnVaZmCtXrtUQBoKxaP
+INqiN0WfSK+fgPQGBeaxqOQWxjndjt1fiy/O7SJF9jWyYG68EToHNRKMiKLkQLk
EF9x71asrC4Ig/3ak2lLanA362E8rbMy1Y0+CgPPljsr1OvfcfyYsFkZaDdJcs+8
Gzknx9bPwTV/Ea63+NrdwEgHsPE4TcTgL4Th58Jy2+PkLmhVtzNf2O08TSOtf2do
2Xb7i0H67Yn8v5g8y1nboksVsMLwqCOe8s1dyOWdYhei+53/S7LZVRV/9EeB84Ru
VuR8HC2eXLQ3s25NHyaUVkOqqVyUCTizDpSnZqs5xc1Oad3CqFYuJYfQwkxO1fgj
mZpBNpMCEQW1VyJEybFUdBSXBU8Rs3VgH5h2wM2KDXDw5JIfVVEsVxSJbdWTBw8O
LDgNHTfkq7qotXpwmkwmqWpqJdfMlX52p0yyr0SQLl6Y6bvJesfmUceNSYK4DRrY
WrEIQn8Qu76Lyfmn3bGnqZSfLtWSETH/YyaBz8qxOl/87F8fZWOAaNe1f9geYtbe
wgHSZHsjCB78eDDwTEICHyIMHDbqK8IkejW8pe3jf+YWKQ9XSHTSodN8kxgsObvI
XFJ6GPnixtIqV1+DLAAimoXeAbj5YfvTW1bF7DgFZ0LQL4x/VfRBZS9mPQ2wIbcE
y96giKyofaARP7p2VXA7wzyH6X+5pb6CCVTEbaVXuleKNAOgT0fSVZ2UrtBq8dAp
HcuVFuTVlm6p10wsSABbnMJqlQ9jLp74CKccRgwhrXIfMQ5bmNb8j4oKWzJsZSzl
yMIWJokNwavrNSGTQChHRDwaG/mXPNhkTW25k7aD7i3Up2QGEDge2aoZae+M47Hz
rpN1pZCXbRu3ayqDhjnZVbjcO504CT5IuOL7iEIbxg5FpZwsiynjY3hcSTspaK60
g3jCQRJoGf24epCBQG+aD7CFFc7P7VxfmpePm82uk53mo8CLNQ5EPJgtpMCgk2o6
nNaO2ANennFgeYJdFTVkqttTgGxYjy8vz9c5hk0sXTq98AUHRRo+tAiGC39yuV+D
S6VvtJWvBi2naDcyfb+MCdTnw29pwRAO4fVv39KKH83yhQdxlSOg1657B0TOrmc6
IaRVxIV+o5DHahcLkxWuAfWJnDg+IUkONZ18cfTtXSNpDy900Zdo3hnI4A1JKxKq
F0tLb+GTMFSU20r+ld5ov3luH9gbekrODoGYxXknSIjcJC/ETnsmBoL1DjYy8ahn
v1KOFfcEdCm8FiwzeCOCLjzsGRGccr3LIUavGTmlN1efbO8wv/bKAylBVgmpwyoE
oP5fSHOI8wrT6EAXEm3y9U4DdaUz/n3ef4JsLNIt0oQxiIAW5sK4MehR9BrFqOyl
xYlZSclxud/Ak1SzMBS41Bxz35+E2V0njQlXM9T3YtjYexjhDX+qW1pc2+s7lNkx
YdkLHWa0b7aRoYpShPaUzca3tC9BB0KtqwjwICqOBPke3xGB+YxDuPwQmrH+Jr0j
7cfj1d8I5rbumncxFEHGKnMeGr3l3721/J+7nvzOdM7xwNSy/JUdr2sopZUh/WEV
/dSeJ0aS1c27oZRDl0btRv2yLB9oa+BFMkGK6BwckGd8uU7nHwY2uKvyxH4Ibwtw
nmzNjlYsvRotydaIdF/pVX37cjtmJrtlePP6esSeYEiEv24uVp0VTJeiibGI7FMR
1EROkn/m+VjtLiyIfRKnJiviuPX8uTIlATyTiZrQBFxQxCiw0EtzYsfOICT+MjrM
bwY2+KGMtIobEqgWiVb8k3/GFyKP38xdGazX9BizKEIii7iBbMJ0Dr02nQcxcc/0
wvBE9my3DOIWFOY8ZCvFgnvADIjAHepn5/5od1D8lhwMnlciY447or0/wWZTWBo1
8zaFaJxKvjGjqfHKN8zlWqx+SHZkVXQIyY8Fxblfc4fxm4/y+IGuNmY/vqYwvrqi
C0OyxZ8OowL5W8qGlSAaVDUgVZMqhZcX7SolQ1yJCzWala10scSnio6VDoYvM5oJ
k4ApkuAOOZRwl2EiFaHawp739yfEJx4lFSSHC0sQJ5l11uENDk3EMjNkC6tBiYw2
MXqeZidO8Ycdw2v4k6ZQB7KkTBFL7GjwXjyWAzrRvV2nLdLLETyN9bPneaCglUE/
fP22B07vCrd8tgPm3Ps0tdtls9EO1aeTfNTv1vRvGcU7hzr0lx9X3DIazh1RtM+N
qxwUZoSnlxkWBuTXlIploNpDdrssM5Y1Ezcpj1Kt4w6kbF8SrCJI7JssbH3BdK6R
QL02Vft+ezavPdbg4+bmhax2TE1HpvBtPewLifVZv1DWJAbdRuauhig7++VBS5ft
N3fKI355fv5v4BB3NTT0F6DH0U8f/AndkXruAAXfVhWgNfzixp2c9efIitok9fRv
hGLLMnOebKG+Dmk2KSt/gI/sQhgXwfzhTMnYzePIPKjMKJICvIsV0eiG3Gqo8eMf
e95y96UpYkcwieynWP29VhKcHR1cFrtj3DxSabTN4A9oGPQiaoJ1p0TNQUm6FQbu
ZfJin7scXSbRoePcBHOWIQSDVYMS9ouvmNBfhVDeYoIpZpmNydh0a7wDP4YBmg7u
JRpDRc7BooyD0EqVaZKhc3SnaO+oPSkha6LEZ4ktZm1KbPcZ9GRUAvbXC2ByLkam
j7wKWOWGVzoqAeFk2JY0fHLTMhtpfXKO96nJF84Kn+ND4NytVb44IrDWEqJvaKy6
/CnqUAKH7127heXU0hKkNCwZPMUilPG7jKmlGxEnunsgacpHVjzz1AthhB2pmEnU
WyewV6hCK/yJtSCHz3NvkisJ0JOiBdkBVL3OwwW8ritNQ1ozHpfA0vYNmSQKGlkk
BGt1f96FxZEyPb2k6or2Vdlp7YUVXvtvb2nrxcG1zLqKvleg/6ofJuu+ERssG+VW
oDDAhpMAfznyMjWg79QmWPrIHJRcbEerOZ8zjTqk+47ygGXJwmAYfQs3FQsBM/Ln
AA+Ppf2KurLomQRWHP8seMAlCvH2asj+jUPWk1Rn51KSw5vOnTsLwvcN86QJa3d5
L2OUBtkwCuowDmYQK/wn105C+YKo9e4c4U+8egpXC5ra8HVwg0/zDOedyRvzXk98
pM9u0czFivYO7wHYlI+4H1i+hkL9setw+/J6pf3vwvkAoEPjBGMqU1lJYkf9KPDZ
pw/I4ztTtPtna2y47oNWOfvxGpKI/FOxkAJhYkHb4R9GNnFa1y38dX2oSaEtW8F0
NaXihhIgqOT7Ut1ELcnUcsatjxTB959SgO+Ne/FF+RoUJTAQtsDPNOp1cdjGfDry
yGYqkly7vOsicthRqlL1DU+x7Qy/mCzNJsJ2RYSxXr0uAIBSSogbr3FCX/2cmWnq
UQnQygqNC5GTwo1iYEK63xSObqPJX4Ze7eZpkj2VFhcfbO3zOcaZoCm6o0CfCMae
hmzJUAAdD9PuEw8OBkFS0cEiBmkzynuvZYI4MQtymqhDNAK+l+49EfcAcnxWJ87D
LhONizrY2dg2I8vyLi0GX+XMb8cNFhoCDyXTfc9zmx/Oy48y5OkavdxQXeHanWQt
r3xWYborp3KPg4KsOOVsLtrXRfHiMdNRUzyc9vDuJ9WObjfAsXSwvhyG19titcl7
s/LFYwaePysBIS9kxOdoNSV00GO6ZvTKZi0bZN7v1a/yYe82dsSbfXSJPyWw/pEs
wXNELuS5NbKBqJ8rI6af0qcwiTBA5ie8ybzpTQ3Zf2UEhevd+oqiKspMs8omZmxT
9RVnOqhkd5jnzYYcSod4ENlIJsspOg/H1CbDtqOuyQX8F/WOTa6DzLhEepG5rFIS
zxOkZieg5ThIOK0+eUva4gZRlqJBaLt05fkKsDnBVayQB86SJ+UCUggCkHswqrDS
TVPQUypmr30v6ndrlQ4aRwNh+fa7+Xu9un0nKOL1UQcui/UtqW8I7WIdUtkCi15B
K6ke+K8dlTTTO7/fjin3UFcOc6+rYLg1ROwrQWuhoCBZKUyDe/5dXBJKIPUQQBie
7wTg9ghFzIfuM2QBWqAHFSUlQQwPe6MP3Sfmn6Hr2NhQ/+Cp1Un15A0TlV+6vKDf
7goyHwkkboFRDefJ5udMrwnktYi8j7RAWOOx6Ue2vdvxOJ7eWXXx5XmAgiQoShkK
0cD+9aGprDcdRP+V0TLIgw68g4WbRWbIuBAkuYAIoC/0dsd5d7uCspSrl6LXiI1Y
ivDVF08Pk5AdgFMuTlY0Kc5R6FVM96BH+L60WMFzW66hLLvRw9GEoav9bVcpkP+q
sYize3cEYqNNZrEC+q35ryFeuejPu+URIHurYygMZsqLxFJaw512yXtMbt0reKbS
jj/+1f9V0055XN+hR9zSSEfzkfw3Ai1ybDK4q2Kk2jvutMX1x/I4d7ugrDJ61HjN
YSbKbmcC8wHpptq8IaEAtllujF2uZAWtTm4fkkcHkXtboZ3f9+nrLDaIDy6/2sko
jTLpyffFjIOwEfkzUFftrEN/W2wlAl9Lmc0/9lBHJgRbRXWVw++KA3rlPRq0d2bF
JuWrgW/uYDsoGWiBcqoW3AkiuLFKnZS01VeQ+4GmHAlJ2+ZvTEQhv+/0T0T1IxCs
aEkh5368ygpB/Gv9wo/e4pMDxuQlgUEYVV2nuEVTYj/U3xJHCxzvtsNf9oX5+Rix
7X2VLGc+6+aqWOo0dHKqtair7XdOqRBvuMB7xDCrd5VXKWQrrKbK0BwHvaA+R7QH
cDkOewsUB72LsprW8dL/5PbyyeuDJpaE/0Xx8FjBjEhI958nHgbh6ooUssn452H6
Zy6t+0XFp92gWROc637rzcpmRJ8YBqLMnAG1plNVXh0ugl1szBqLnOygURlnWr+e
21lrPiB9QzJzCjVVX+fBBvKCeEOuiecPkK0dDc4eDkCKcJRXkYPJqsjqBki9eEoJ
ph368Q5ngi4QHEUXWYX3eGmbF6rd+rFMLQZNKxhRxXaeSqLe7EwsEpY/GTd5qbtS
ERy6omjhJtKbBXqjxFUJtZXIQ42R6+/zQd13X7yk3Nm0CJqnl3gheoWya/zvPOV5
AFtWBYSfURUpTL31d5tY/doU+ApWKNe6AnLef98kJcL2uSTdEQ1iDVENo6hsGX6k
/YIDODCDdyX9CoDLEEbvNTcewTnJhs/4Z6OZxMLsV5djsX/h+pGoj4RG0zXEK5vH
9fOQrQFqOY995cB3kJUC9ep/DrNaIdXpCmMXaTSsm8C4rtWfo+huVKGMzGmQ6j1k
EoWcczCOOzvr4NJJZV0RQWGdPZ2iHSLtB3sYM0RTpUfGcvcpuX3Ele1kNcais63i
fozcfVrhSlcmsoirM0WZqjJFrXUyCc8oNybpjVBwx4ZMB3HRjPhkawdjMKv6pbO1
izgq5ezwjpLcscILuS2F1eLCwGtBamRN8ODRx856kLmKpywsjpa3SO30hNqSlogN
R92a84+igB7qn8MhIj3wvdwHybeLSatqxE2xI3uCO+rMoRET9TUkPQ0ytTs5psA6
qxmY6uWNdGXMx8PiPQtyBc4Rksn5TGdIU5w6iB5PJtVgOmSk96+2IFYGERyPuy6B
CLQws82pfy2/YcS44XqjM8zZUKIlOoP46wOBahSSl7+SiMcdCy93c7UylXNR7qQr
QNdixhBd6p/TtHZKUWUolPOwTnKnV/LCA1ovJqH1rozafVl86+gcYtYCu7IUMDGH
8vwfYmu1lE8Tu/tjX2j6tG1bh7ZyB/MRXdDmY+DjtNuUKkdE4B9a4fLXFx4GGW8W
d+hXZrlfiB2zk+zqS/nk8j8AygJPO8+5btfCWi8xOwHz51SzvbFmypCHAo8LlEPf
UQ4oz1Da7jV8zEy4PZZ0Q92yctas7o30WeEeWtgHtjj3nSjRxpWGMpd+Cygn99AP
gBl58c38eOrAgIjO9xDvwdSERtcLjyplu+lz6W2FfcKf7izISL5R5l2rwRS4yI7f
twOjEaMo4+sBfoDQYDJ1iZVoHrIKlXwYBzYl9KUTypb+PRYZmnPAZoijcNGW9P5h
ecJYr2S3OqR4vzglI09BtvCsM5NvYUhhEM/+KnoaDHiaWqBiGqLcYOaizjr1KSOj
La+4jKEQ9skAcvJSX/Wl2MFz2BbQTpAKO70n142kzT30LGPWHFvSbXGOrzEaFqyU
PSRclpwPvuwdwKkGiC9jOd59t0iRiyXj89RcA7KvHjkAP5SEMfmDTLbbnGpNEPsy
oNFbIZiYk11LEFhQEcnl6bhJfCWRstLYDapHYJGu3mhVPNCL1tYpjms/d05S8hC3
AaDlHgt0of1C2zXQ7jjVLXjFTIT/yY9abNDUFnZXJBvY7yUl3IDmuSzftmHRMHyc
RfdXL+/AGkQnTgl972eZUZ9A25NCyxDQCnEitHAVn6mKhPD9R7P+vSRtL0HfsdxV
k5OOIlmZ9i1K4ce8KwJIrEunvLucb+sIsW4QqctWcQ/ajRnsEA5GhSjtgFFe8oH1
mRC9e0fVTm5GheUqjFvd8R1Dj0Brr2/SuhMIG7xkaL8Yl6AqK8oOrUeFitOa3Nbp
ROL9zvIGzzBtcEGP6DQ87P39CnBZl14Y4yiVnFqW9qrRmXIh0vPujNt/om4JxLZJ
6/BY6o1HMb6QexQ00a+W2uA0qmQPau0URQrMUUQC9/6BH47BJBEmHrUgNCdBr0Tj
tnXuU/10GH0zGxMwOzn/EkoF1IpCCJ1qvFEyUoiFUUB0pJsNjMu6WqgWg+tCroRN
ir0DpN1jCNi8gD/latpOwIiLq5t5cG63LrVMAPopQOicH/HG0xVFSZcS501fglaE
rTfWdZoRdFQqmi+f0ZYItHZYAqzDr3aDYffkAIzAJWi7PyO+DP3FpNXqKWAXMhQE
PvI20obu47YuRRIWOJiCVonwpcdq8dMd9AlZoA1a/NV2KO16uFDg+WUc7jWuBbSh
rBciTkMB2gORel6MZ6vPhm8gVDWf9JwFppSsGl7BanzFB1m9QwEkZ2PkPPzjgTsU
V5KKFk5F2jIxmbVin36UdS6yIYuQKet2UxCtTzQ8TFdmq5Gwu35/HFlqpcGHoWnF
Yn5XGFEzhApztsrk88nrIN0TXunr41AUsUN9BuA6cZ6M/46joznxNNeJlnSm97Cv
pFZAobI4XiHooWgdDCf/saKUsJstAqMDxv++UgLpSAJ6s9zjfox/EvbXNshtwomG
twexDScSrGcpxUKTVKXvlv2Ybn9r/gjTCaZP6AtljtmeKIQbPSSgUY8hbspjAUo/
43rWXMOixwlXQId9tKkN8svZiA7sZyCWbZKzQ2FMkMYn3XixarSE/ru4CW8AiWk6
aZrTHi+qdPUuvzGugXhhu5VsSezESlsx/dTtOQd+g0Nu1sy8ItVF6WyUliptGjR3
JhHETh5X98GrJM+u+kH6wIymzW+E4Ghb+bah+22pYoa2Y5CpesR1wG5AUKId64Vr
hZ1bRWGggz8aJu7Gat7fRUrbjuFY+hfJ1UMldmntTNS5sKjHebNKJUAExXHocnem
o2lz5Ki9ldl8JaWJQAHwBbvVMB3gs/AxkQuVMccEavdImnr57SWhJJyzplThdPDZ
LZA4RaU81qImXCqCqNYLRAHCDMq9t0cAlOglMfVvDG5aT8EVcW5jInEL73IOXaaG
xNaojLtP6kPW7w7xSycJ+u4ov0JIzrBQ3owGfXoIesXY141MYtsOVRZD34pLhI5T
4kwvB8PpQI8KiCfguh6VehQxX6Za2E/VRTtImfcpKV31GI6SDdlkWSTgX0r0GVZr
APk0ZYV/GhVdXf8zTrdHBJ7e0w+pxHcdV7C8QxRjamY2gflM7KNfWb0s0hzb8hId
MW2ZZgd74jg6rmNzo03y/ow1DvAdvvNZhLqI/QYAjowaPPp2gZrtJ8h9qtUWPS0C
CEcs4MLk+D1xWH140mdf2iA+TYk4v+M+jlss1kPEwnXefyEw0c6W8e1TLGgFgz4w
RCtCw7S4y5y4GhJnO4Yai5YPdtQLakKIQlFO/v7sJ9iA9op/n2X3iG1YQD7IFnZc
M5Miu9vcd/sHI0Rn6dlGquZFz/KQ1t9F4jleaRFM53JZa70owDrFhQntkrJKpI6J
Xkg8YIVRWBXQNA7WvpBgWAJMdX5FJKKeN4Fs9O7Y7SzI7K+YY9SIjwfH151StVUp
PWamJ/byioXLQ9lUtgMXKup741VOFonBP+udOCtyQ86AGrt5QN41LYfU8B9XPlvq
YmvFBlioXqb8zKXdc/yKvUwocCTNe5HGKWYnmpyuIX27wFRi3bpDVg2Bor/AJPha
+lJek9gLuTuCco5NvDVeMSjMYQPfArRQfhVm2GHRgwSnMK6nHhqRpKD9nKs/dZdM
sov/fnk/Uhu3V8/tpTXgFiq36du4ENsjtPaIF3waqVYGPQfyhvv1BQYMLpmxNT/1
qhLVChayvKalvTHhZthBucmLReUAjlOuZ9zpIdzcfRJXEVwsV/oQP/1xvkv9ZXcC
4i6UqUp0Mtse+oN/AXHSrBbueX4AIOKFVC8qhvZP6L8vLAKHSUTwn2iadvoFZphm
tFI8oQsTQRZ3pR487rYDRQlzL+Cj9Lt+Mh7EYHE4G0wr/zo2nVGDm5PbOdi9/f5s
g8FS4SKyWEil8+ppamFosJ/MuWmWNjEhHGMwQkgRpGwk0AnYq9O1G7auBaP9Dvyd
G3VahHZeZx9bCzQGv2WOE2MpgPM23Pf0Eoc206zOUFp1bZ+2epsZO4xqa6HVM0qt
ZMhZLoewI+W60Hcf0+gIxuG6edlNxDxii2tW8jY8CI+tbEtKB3SkHuFppmTK11/Z
2GKkZoXDGkj97hfcfq1fBRhwd8oiQvMCzew1gJnr2Ls+8E6lmk2tSO6CIpnDlYHJ
sljyQnd/xOfEWQa4fMr4FW2P3ogg24JxLQXzGxcVc2bc78aWf3zoVkbGiqX7jel3
tn+5WfSirqZzUFqhKuVgllJd6gOcmCDnLQyGpOgipZkCWXSxT3rx+4lEZuUQIEm1
1hncRq87eh7qusJ7NSqEQDY2xK8/UI5lq7qC67kEHf/5ljbaOyCcUPQ3eaoFvMLV
+ejErpSqTc81LnhgmaNOdSXmnXZP7Gj7b8lWM5678n1B6nz5R+PVyVcRP0JKBJVK
8g9Vwqzjf/nlOqMVYBaYz2BquCQZKsXvhsJO21Jw+TbIOrMTkICmnWd6ODUsSs9O
9i2RoMWOrqiA5qG2eBrX9W6jn6RBmxqbuFGEYz+m8baiT10bvMH3uQrNmW+svVNP
05xQcEHOAoi7f7bwQmvyv/9BOw25E6qRUkOVuHUVJ53MkYrzgHiKa5k1Mf7prDq/
F4JNm0x//Tw2smY+JwHXfuYwAYIVOfeDKGnQ0xTVOZ7OVkeyIadpRk7zbU8RF+HW
ZCQgADc3MAFnhbovkR8tqLBk1EjOxS8qnjkXV+oNbJs5EblLbC5/99GH1flZXUjB
HBVEYlM4ZY7qkm7QPq47HmlASryFcoc75nHF1dFcs06DffRC+IULx6dMkhk8iAut
XzZ8oTnic4LcV8998DfzHjgDf9mQ2vEuwlhS1EOiHxVtv3i9X5Jr7cIJbNMR9OOM
aioDTvA+gWCUC3885/i8WDdSsDDHyKIq0Z/L1aMduMcoihVidEK/E4EANiQ/9JJl
mvVjlGqXLUaD3wU1m6bfXqMhftkJMNKgAAbi1rXPMAEbG8qeb6O9Kj8+mWR6ec8e
JlIsDzSzxdrPMRbnf5wFldcqHUQ6P0vDAVi+fj7g9KXppOw7LdZl9Gm65BH27kHB
8QiGqq54k593m5aAlVzCQDXDDRGpFu0ZaYWUsDLTG4KTvfP9UK+8Pgx7yejfoSs8
b4quyxRpCBXbvn0Lhv/LQ0uAVTvzpcipOu2JB2LgWfwqBnkDjT5MyUBANEbUbtQj
/jiSeEnpLv1m1UU444db8jbKX5aTrZXneY0Zeado7jyif+sjs2cAIurD1d5aMAYC
JnOyv9gaNHK2nCeekc1R/4LEEEYEz+IYfcM0blxrO55tNSb9M9AJsNhAozGycBDH
ne8vMY9U6+3z6Lg4vQSZUe/a6EHcNm56pbAvvovZ40DbmqB4WyGMXoHzRYwsr6oC
iybclKGWxvC2e2D656V2QAXKi5zycg7LNbi9M9ueArZaY4lgzyUFjnj0C/fA9O2D
qtdsinhvsWWNVv+kloUy2vecidl+LW0QYQVJNgB8YFIooWiK7w9SwG22NnkxsF4e
purvEHHc8uXnh8MaHq1Yg5YeBkPsIOWUdkkY9Qf7QQMDeWOfsBxyyhXagj4PiYxd
ThFYS0EdpeXNAcWVJBUN7fzEvzb9iG9QRRuzwLzmU80YqBxN6Oy4MfMsmolq0Jdn
Enuxf6bhafTZbyJWvBf1b8XdHGok8gHPqVtRpE8sbSfttbRNpUt3CyQ47gZ7UKy1
6jcwE2mOErZJdi6EuYIF8y+4dlQwr4ZrZg8UcABn8bVU2+TkPLVKVvAE4SSmoVFd
ql2lvSL7t+BvidWNszGT+EeTsYrrxfssLCSHCS9rsQVEYkCcIJW+mRtqcp8ff7ez
/y7sGUAjcGHIaZ8PdboSkKjrYxz2VbvnmV5b/vwAdkvo0Hv/2zxSAbXDveEDDm/B
o4HBkxAjRsXnZb0Z3PvFFMOWraazS2X3roz43ijyYd/+/SFiieiknL7RAqDugNbJ
6Z1D/VUYHAtzidpbemnmqmHGuHHFBC09Y3IF9C72F4Ru/ZMW56/tyMm3bpOQfhax
BDOd5PFO1EuHYf9PBZEgoyrldjIqFWfw1Md6lSyZ2HEq4Z3DSV2A3XO3OpGCc6Zq
+XNUxFF5TwSqLN3OdT3iQKoYGWPXlA6sMiis9+QUIKFvebpwkllUuoCbhq7xRkbm
ynGnsJ7grm62mVb38VxoF40Fa91qLavlA+jPHa1YbirMMgt0QAvGgVBzZIQL0bzG
CyEtnC7FE0tjE/Uo7jRGylWp4gHrKgc+rTJvUju+NE1/2AKPlqTEvWGEJafjzbZw
2N/26YDVliaM2Uf6EcVf5fxM+3dsL+ilLm3V3+jjUssOQYwQe+y0fhJKyHrYa+vt
uJNW+cDRDn3owSbQ3CHy41p945ht6k3fjkUzc75Gup1jQmd1wnuHs4xU/aeGBQ+K
WLGJQv64vVbzk5CiQtv4Nreg4wT2NeQlrSFzoMMOjFT3+nlJpVemlJkGmNh4sZoO
E5WbaqaYLGtC9Ug0Suwd3KG49WkU/iQNp3KPaZxjSuFNNevzyjLDrJ43dpvd8CYU
jLNdjhJgO/5D9oerVvyfVT++ipTEWm3TU6v9BHSs+XEWpfCuUIJSU7IOUWTX4AWw
emLqhDwkIGXs1e21YPnh/YOSelaQo7xZrSDgPO8NcAoXQ6t7h8tny2CxSMDrrHNu
3Dm3tZwTIJk3R2OWmcaFB6NZY2IxbgcN4Vv177NmByvp9a4nmm7Wm6JbmxT3iev+
gSWsIHdwKc7VBjJZnCoy0DxbtX1sdnq+4VNbDBj6rm5srRHeY4hGiRcybJSAZpA/
KUG+bRM4NdHCPLe065xCMy7Cg0HW/5zk1gr6hVFfddOYJslzp1q17IprWtw5sg+G
PazEkhRgV2XxqZSptmtadsJCQzIO6ji04UaRl7aTPSurQLG331CizE/rgN+4oaYF
YMiMYaBwaubI79hMMnIuBBC7KmzG6vuWnbf65JR1zhP+KQGdto88OFiBiJFgovvs
RUEU5I0uFl1cpXok/ZRxS/uyShSu9ka7jJwk/wZtnU4ZLvWNk21r/24/SUf5Bawr
qXtkOnx7wh6YiynPawfxKCUWVz/rKqXYwSA7LEEJ6TJ9pPfglT3j2s0VSyo9lkus
gqlxOi5yNNIv58s6mbax+jZsyDJ878f1xqnkVpZf2P/jSCPqItha2L1k1IIERNWp
BOtE5z2B6TnVQTc9K3sDt97Kjjt6qFiSxZC88qO0VDLu5HRlRhXTT5siFtRtXa8M
AplvO7DiAcSGAe36EyHy1V+z5Amzbjk7kicekADkxVQHTns9gKn+z6AILNTJoHsP
m6I3KoJN3evFduPeVKNwlcK8NMoTJEKynKOf2LGAwrqd50IbChH7rtm1HVMLOqUm
vaTmjDA7GoqjCX4APLmKqKVjzxuojU5J/3XLFE7uYjJxJXoxNcIAJpNzqxGsbOEJ
dUsMlWNGwaQhF7fwpZqknbh3avK4VHnPVWPxx0xzEGmCgufqvKglJ6rs2Z5E/dnb
Zyd/WijjUlq9ufqHgM3Pa0LWgIdrhKTJ5OYYmnNF9v24kOB4vYIgS2Wts8AvBo2i
y0D41lTbeyf/qvcSWcV3hizOO5hBDSr4ZoC8df660ixqITFRcYPqAEbZ9irSPNS2
KkRaGn4F0UNynDPA/WV9sGhgXvrmOoYbBSy5HFFHzegg67JlvXuRvZxC0KBbWBkC
nNFL4AHVE/MM4V6IIOnmwBxA+ci9noAn241ZrvFop20859oX/F52ZN3UG/Jq+Fp1
FqxLTRqVDMVimZJkTQsIWES5bxC4/Bc2cFrrFz7Gn1VV2atQuOxw+9zZ3temfi5Z
EQx1YZgUc83UnzMuBrIXKtdYbaIRpnTuFhQ5c3UEQ3TATDw7dnfC4bOE3YVd4BGe
nTbkKvpc/EWWYh7mlH/1AWfnZEIFXCGP0nMp/Y3iPs4A85gWR4xnlcT+myYWJh72
4at1F++XHpnpXc4865WA2gnDhYhceRcA9RgBX1i4nLh/WSzl42wKgRD6asFsEcuy
vjxrhXbIIqQnA006DrojBGVCSU75N43buB/UiSRr7BpEFjAhKeaq+odfxP1n01Vq
DL2WERufcQETvkI/IlP8SqKL/O/fv8M250eiq+72hOVr5YKFNLOT5MxwEZeMy/qz
JGiPSrWdkKVqVPP6+tN8lLpx9OMLPUEEURn2rEfs4l/ddgTwChp2o5VFBH1a8iGQ
6s4RbzGC/XzHumpZNvhbp5/tCgDJMsEIxOOeBL2ZtPQtOniBRWz8CBkDrnB513Ko
7+5EtxFamFct4rm58lRDeGvwFJ3FXzaEL5mB72HyP9PFpLtprBYu/cjDWQnmq8aU
dTCPiQoMiwIwQzNkTAnaEKg1VIGETpZhp96/W88qfYXfFwfKgC9gJQN/azdGVdW+
W/YoLzyRZ5BUeZ5lc1gi+3hTWNzfR/WnZW0qvhU9iHNTKWZJU2SHJJ9iFkXC/zyr
ZNL5jbgivoRcgNQZi4KqdHTNHMU/dg1w9gwK4h+IxZBYMoUOllZKE4hGC8PksRRc
00cLHWrpzrFaSFBEITLFdLhecfC1PcGidPjHpHWvoCAyYps0p1zk0R2Xmj/gM6Ib
D7VOBMEtTei/7kZuq2MIXiho7D6aSgtbPK2owSp1yuvRrGLrfsSVj+NT2pcekh/E
lK+nOYXiCo/MbF0RTYG1i69V3N7qw+LoMIt1618WdWrOAlWzD/GEt9tbhaFGNHIS
1C9RkMh6R7weS1ykJnfWou76MDKPRG9JGElDs10KRsVy4uATBnTJl3PQD+14IXF4
2JDKgkPURavdbCh68Z75e7MYWpYfAnOJ7JljD/wdvtKl+jsH6FMqJejwbN/BHe73
IXBBysdBXrbM/YP23j5Wu/1d/kBG6rxvSJns0dMpUYSDP5Z9PQvk57IG/rfbmK0I
cASJtswedjQLixx5gSNaJhl/ayLS3ObZAlcw1wwTox3OByjqNni2rJ8OhgOcU6kq
FUD9ROA4eLqUpGJAS6A/+MT9NmviWWm/xMZmRJwJrs88rW1dK3NYTvebII1ybHov
w4rpOSiPNNNHyhC7MwMr+mD50aX1s9zN7A2gjM7ZRGzZ0wQNKUPzh5QrxU+5MRF/
HuHxwzo+LHoMDW5lcRw34ab6T5TzSmaMz/+Vt1e9/+zVIas4i/g/FzNBSdqm8zJa
wHet+IHmTTWwr0Byo5bVJ0r3kfAU4q1bexQFWJk1+pOGi0svMEyY9czDxBOGXiLn
U6VlbUJNx6Ch7OjPBmoY2jQt8pBg3TFa7Rs0+bDjlkKG3wryeWWqhMiPv3MMKXfy
XoykJsNpFJ6loWwdtjz2S3qhdPwPLCVZP0ALzVvRQuEo690sXkk2nykcheCsNFdy
G9ITi03DO5uadddpBuBh9WHltRG/D75wm5/HpXsJEgTdfw69ea1jNTUpzWcwNsYi
SrzDfeEWVH+PpEuftCWqrxmPCo0fzAm0deJlorTMJn2fGPlZqFFVK4YUn8rfAQLP
eRTCxZSiVPQJzO/qLgxUTV3lhoDINGs01EoQR99ldABvq8N7OGeDjZH78LuP1RVS
AeZ1SeSQ0rtwAIXUs4tKEc9nUjE9rA6SXYA57Y6X8YHRuCDR+weFLg7Zxwr/BRlu
OCKOuwJkI+Yi73Hz5GZlOzNwm0IXbqDpag4LZ0ioh2n0Z6un3eEo+ZeSuASQOw5W
4CsJMQN7M3mCc+xdGaBKGEpHgCrvwySav5r+NqJK4epJOS8wU1dsjsl0MnsOFz4Y
6GRqbdjnk2O1wWF6zx4viAGleSXSWQ3j0jnmOHkhAXUDkw0LRNEekUFuQ2jxnpnr
NJG6wwTjPVJ01h6XVwiZ398+PsJ4vEFjpUHHYYOMsDNwTG/Z5Z1jTdDutvlOeRzo
PiJ0a4GO/tZyiSKwpWyD+Tw+CviGc6UL49Wzz+ziOPNhCP/seWPJaxTkMh0ptLEO
tKDIj1KpCDHYauMkQYpX678adSMZU4Kl3E8hZCxmRvmKEiYVjgd1Kb+v3ehMBCd1
XDwFFhmhhsJN95oy+WZJ4UElxw9oFUkyiaObnYxjkuiR16iJduh0900v3ED7tYzv
NXhGFwsh+b6PV+0TPYRatWqPURTL5aF+cSh/PH14dCe40XwII129GkWsvhIF7fJ8
2cSIK0rZOpJL8qZne2Y9nD3sR2QMmTygALQMWOqlhIap/i1rnXwrfx2kmWc37DL3
NEF9qiIAQSZJuz8YVs/IMh4WFvWMH31ETFgGLWNixhmtBMfEbeEwYo+5jobcRW31
SjIq2f+TVCeB/vpzo0QJrnAvI/4/A50ry9A+WTfGyFUCXNNHAwG8oH7xJu27uhsB
VNoUir/3c4waAAjXi7VY+RkR5+G5n+kHKNQzlInYn7+cTvUhB4r3xe+mvwDE3p4Q
Fmn2uFD5gx+JNgqI23oLaXHlAJKiPctlS2HCP7WYy0YtcNIEI/a2vHFaRhUuVGcg
Dkq+1630ly3mCL0mJAxz5pbQYT9l7XqKSf7uRDawGeDg42wF6i3MNPncQ5ETGzbs
2MemfH8cyZ39yqshi3KUQX0p6uIhuU1q1I9pH+8Xwsdeo9ysNAEJ9vl8718etUnj
+QpZ4DSyBJS+0Q7Se+e9VdgrcyM8zTN7VWi+ItMzAMArO561Q7hTnn4nrfMvB7pa
xSE6aMkSMU7QKjwL5Az+QLTZcnuNEhCXUJdoM0s+Sp+Lx1OxOO3tXBdsU0uSuOt4
2+rtn5+f8FgYc8/VMqotDYkPgN8Rn3xBNLkivs6GdVNwcoy+hwZaZzRIIgD122FV
4jygmmFqEq12dLbYbDc+JXLU9fbKdjPbwm7oMmDuVGtq5FdcwNuqcH6D+oxg+QhE
s5OgxnuRtspemZMWddDze8QObPeA5VffgRji1zBstSDm3dpoqLnC1iXmR4EaCRra
KNtFmU3u+e/gZlEfTV7IHVymF97ivNqFbJV2+PT2TN13p8aQTEHGGDQ2T92jNxxx
f3NH5Cd55BZcUvRT0WS3QQ5YpkuSA3mR6JWdGn8U9j5l2Zv+0tkJz/o37Lucd0eS
i7tkReoDhq0wzLqN+s3NT14tI9HpWkQ/1+M5GgxQ+QEdtUJ6B/oyIXlR9+Qj3ct9
lIk2WcPLJn6rAXJHIsJcPlzXKXotA25S70RgScDV3EPmML/VLIXdGo1Sou/FjW2y
7hXllb+I89++CAxahzhOy/AXtsiJSdcwaWPcDsV1lzJCwj7LjkFIETF9sh9Fyoni
+faAZJGVOBG1KPgvEXPdILfg7Fdah/muE9T3r7mbSfaxDpX2Ozo3zsUw8qucpBzo
3JEajRJI90iUtk/XutII79A4jA3u/gd84GOkDovjfSuSzgMcQg3n58HJMv9z/4oq
cuBVUWY3wmgv5Qps9fUDgfodXP8iac0nR4QVBo/dSXOD0gme07L0hu+UuDihmAQK
dIUssY+nks3l8t8TEKu35STZqqdhM301oU/FWzow/cy9X47c/smoY4jyQXGp00ww
wwPcky3OqYQ4fy3PsUQIx7RCCcatJE+Lf9pP+M/Ogs+mnWs4n/JptlteC2JEaMaL
kf1OGD7F5ZicdWMScemjC6/EsXjSHF3bEVrxLAbSZdfnNe3KO7JqEHEgQf3mNvtu
QAPKnTExYnYmUqQz9Etf4zjI4oNfRMYXRhNtP2SV/JHVzIo/LBURkl1hWTenlUPN
8X1n5AX/QVJ6RIDGZ6UoFoBN38sr9N0hmPIRNPy96eoeNIncghgBb1W9bO2p17HK
6NcyIc/EzDivBmBw5XFjoylYfTsuH35rkJz8bNwW35i67Ba5v4XpVGV8ysbpzmWN
PklJJxQyFQr2KVUdLxobcq/MT9WxZ+Cv55ULWebMj6ta7HWmxWBDJ2qKfedQ6FM5
M+uKoszA3eXvKKBXHM5oQdHyV3wSNl+KchwbHSBGCrvKJJoqq/MXZE1ZA4ga+HF/
yFXbLRxvE0EtmjSEzhezbYLsc0zRLL2cG4hgG54emIpZiI1hTZy5SHlMTMhQslUO
RNVl/ftkEZCfZBqI797doGfLnD0LCBdbq4513M/ZiXvOleBdyM4cVDC4/k6RmDFu
XBwWR1c8XORmM+ENxbJgg7ECJzbUMo8vqhbP5jVpkXvrOANfg1zN3yloZuLVDW4e
0kCIVNs7oAEd0m/ucGPNZhGNgdCcCz/As4qMLhF6BCSXH+L/1MgVXt6Wk7QWyp6C
Kmpw7iApeSJYbk0/qmtaSrO3ewhXDe9ZtfU59IMj1/iqtclLTPuJdEmFRN/20Qmb
qxZFck6FtiMrhE7tDqwEM0QHdawSNjdyGyfMTZVOivEnKaxogMX0hwAcXFAlvRVd
Cy7MWGHfEINzSzw50GOoYw2UPDUCKqvvVvO+SRm229/RyIfBcmSI/rHaQgbFlKdD
VzMlsI/MkiPRDxrEMyquG9VFk6vFOYbMmT70PWLvALAS9FQh9+hsc975E86lSho7
TkI7nQD9ACxo1+s7rn0ghdGYFCKDDhmBYikdXg+gGOxu4ZjEsUmAqvll3pg10jIW
wyWt33Fpq/l1KYDvPM5xEA66GGGh/ju8GE5Stmrp2wtu02l2XhIofQMQo+/VCvtA
WtGzoX5xYH7Gl9yMZ2D4ygzr25Ona9pH9AkImKJp4WXmISFyJgghcV5nUr95W2Lk
gNz0gyX3sP4wsiMQ5EqwIDQPy2R/tqfoHfUlkP97zqWvT0wqwQ6HxY+sLzubFeJm
6gJiNg7WeJorNh7FSjy3HAKPlxts0Mh4IfDzhOeiCcQ1OcdDO9/+lbkG8k9ppHWR
JHCxYnkzXKJNLTjgEYqBMoJpLTsNjtKDs/RJ4Ej90m/soY+S/EVPSwIsA1S5bxr5
26NOdzD5GvSqbaerqrIlYEQjTdFAfYuP6XONuAPMACzlb7pBkKL5ofRbefdWjRPS
bUdhTAigJ5FuCkjbwFnrhvvOhkTa+Psua1+Bt8G3FJJ/JlL8GZ58w3vhSzBGRDT4
+lTC2nomvs524kJ3ldf8eolq5AVHucMtgIxMvZNo/OuB+2s1qo3HQfCfPIxWu8K4
EfpmxxFhBhmvyeDQcNd/kiVH0BRWpbhkFc2+c7wOsgcuB7csKGzUjVF9IZo+LVdN
MLXRTfeeImWO9DLiloREWTb+wQ6p+Oq62ADW3K3V12U6KuM8LmomQ1/KHM06JhnM
AEbyHzEt6DOgK+BSZMoOcPBg+X9oJrFilhE4Pfj6j/jTIK90gjPg41DsiyS0o59g
kevOE34YiDSWuPpCAwWTM5TEcEqMD2+R5/U85Sv7c9Qv2BDSIVZ8CqUYKmUmPU9w
mmdad7ZLP01QkJKmBgewIl5mUFPgF7rzye8nJJwglX25jlerMymSI9BYB42vQQGy
8KcjgDyp9CPJTqgfoMMLJ8sJA8QTztUz+cnH3FhGqV/mgj8QNwjlBXrpIuWBS2vt
1sEilPcv54ePop3s34CJgX3tP3wkRZ5W1IbQ2ZTPWsm9/wNjkL2+ANgAAVvYFHzH
ATcBl3bkgrqmeb+3Vxa9tYzHM9YrRw1bGghl94YY0e+70hj0uJ/ao1ylBkf+JN7x
Ibv7tiSyqhyFdjyUjCEH+jk15jPNMmvGLY7C6sSlNNYDnRV6mns3nvXQQrwR89DM
mKSWM1rRj5q1M/S5fJHSmgfXEbk7qJF0BwSDe/EyoZQrw+ANZ3VlHTkwzFLoFibQ
97wTOfng9WxzmHU9exNgem2HzwpAXP+STfGqm2EfFfBiXLDLsW2m/RNJmWN3ZbsF
QfDCGqjGhLqsw2pdsIoh6iBH41VPxFe82TvnO2pofTat5bQREbjk8mPbIAsK8wZT
+4IxR/LUXqcH8MJsps+ZeSdwtjaGeMRHd8c2ALupiMB8Sf4RvJ9PqTzxEGl5Y9gA
2cNfZ2haqq/FRRu4aqc4+H1KpnbilWhkOVrHgJpKMiJSg/Vd2YOgp5qckePNTceQ
6PNx/NMsfiGUd0VND7d4Z4gd1i9D/ZNmgBMIf7V2DUloHvZ/enRoqC5ZhwAyX14L
g3PKX7xBnwMlpZ0ty2rKLa3vVQFI0mv4Di0Yy403kaX/duPwry4LOuV2Eodsj5IR
0L3ECOsBA5y3UKGTXa86OVSoDvtEB2jrsDO7kGKwvv2ufYxytvR6N26bR+jfNYD/
Nl3Q2SYBD1hF0MT8MKkPWCtaQREKUj336jANff62HYphr6bXywMaMJXuVEQVloQA
Xz4IfizO8UK+/LapJ41K+cpfLYWo6norQb2eeglfA0ucrec/0Qmn/gvRf6CC2m/9
Dt6kI1MIC9GdvT5YvyVlRl32Be+XeFAd0oQAmUlyG8WZTCA2n1hBo4DeMf7OjVsQ
1/L5yvmi6MzfKKSAAcWBfGbMChLshiI0oyPTPvn+mmE08USQD3SiyOsFGxkyjEvQ
26/+bgGrHJjySMGnlNWR+UP7CKb/yjHjaEzWR4o1i83nm6a3UqvS58mXV+zJqNpR
gCQAuRGw4l2Ats0w4YEKJYAj2V2v5GiJIKVNrfpV+/QvAC7x2fjdRM9uHTWHn7BR
Tzm9M3PaUpnSQaMrSKJXhMlhxOAbU5js4hmmkjNorYlo3hStovSWB/yA+mjK3Zkk
5bAxRn6nsQ8z1FFj5UgY/WiwGYwqo+iPd//oVrKTOKacdHshUrUEXVNIuG/Zgs/O
C2mi+Oz9aJcgDGU1RWvskK3pJQqfvztWXZ8jV+LyNA++tIw+4TxLpg4bRVE7Mchb
CnKo/m2rm3x32mv+YboraE940nv99RfABNwpIGIBu2tSB3fXsseRSQw7hto/+gXv
dDUaLOr5qJl2Sh38EO56WoYclF9f4CDiHqqOkz6RkTPIqBawqJea0aCcoDKOR7M2
yrqF003N2ZHpAnzPyzdZzWEWxvJQTtm6NhlHNHZRp4qqnpBUzr3ZTeTzZwrx8Z/b
fHc3aWaV3QPIoiI7nRKmUb8831tFeWFYKQsbQKV8eCHh+0zXpCS7V64R5iV5kPwL
xleOE/2CxEeN2grGN7YIw9hpEewdS0uB3FCwnw62BbLStPCJ1aGJzGvABcd7xQIa
7co7/YGLScFbH3fWIa7DxslhHh/IgoKUrrvp/Ez+oH0dxoFrYb8pOe8C7c6bmh0M
0pWKeHIwGcJweAqKkTblTrnm9AKbyI/AM6MSMq7hwuPCPgqyh+lQNojgbtpJvLU4
bhxg8RO4N0vE7BsMkumS5qdJhwVf8tZItjUZa8CafSU91cnVTwp40AdP99Jnzmgg
RZJauS+IHxkPfD3rbLHFG1MTqftsACCLz+z5aBndX3NGEaWpAPwj0l3F5QthDytO
7V049NH3Yz8Zt08QbVFhNk0mgSLf6ey2jim/2ppOE362jS1L9W3zRjhSqFB5tTh8
pZNCVg0//gFghXRrnnWGh0LYy8lS04eGYkrNyK/jvuw6lxyejxYXgV++dx83jhFl
yz1UZanMStJFwNympYKld9I/VoA6IJY1+RywovTNVtfICp3uYIBTxGZdQFgRoslH
w0arywVj9s5l2berBdtnYvv+I5g7WPnCGno80pW/PR7J1HAgqOXgBO3BB/5Fho5g
CbSW1FYSwazkU8A/4oWOMwBArsprcmPu4ZDRwgmFY5JAWqEDbWDOuCsm4MtxgBOw
1NPbmpEs+CbF8NgQEA+e3qM2CJc3opXjJPJNw5FulRrD6odsXT8VI6L9OTHw7+kX
F3I2DUccpWXl8wEetPVOMpi4R7+LAmWlTYSCWEhGwUdq4L7juRZdQxjWyBULDCs6
Wk9s4RwGdyJ2g+rOYXt/LFIT1f31GPrCct/02nBPtwlJh1hFvxoLhoxb3OdT6OSk
6Aw6lm1SU/KfsfVgAeYiErmoBVVk2kGBbD4ZfHybPDY1ZI0kvfxgaYtB55xiZ60I
lvlKkpMQ08q6Mw/eULZtgYlWsM02gK+DqN6aeKfUeuAUDAlkyOsvMKMsGbYnrxQO
Cpbd91K/0zWOA5yjoa1fdmUuyhefS4sZM6ITPXpocspqe/kX+pVBfZbydNlxs2U4
1eD5uL1RNosFnPnL/RM7cJTLgkXmuk7RrRAG3zgd6n+MP9WAJqUFnVrWT3V0lvN4
CBv6QkDhMlOQqJb5nmKRutj6UH2zVePRkONGzBJ2DRJMWwgTATVQn45nBVLyCuyN
AJJuoerB8YpPxn3xtyh1h4pnWTQO0bVQ6/Nk21wAiirTe9R3HtxiqQlsyd28lbi4
At91EPPpnEp3lOIF/jUxipKCD9iQzXwjJ+DHG/6Y44XrkJKn6G5oVSEbe0+qf+tm
Zic/8hCrIj14nkhnSGvFllDzSdZZPabaNuYv24ekYsYroqqYGgcDe8hHrBbj3Olt
GvvR9kmrEG3DDDVmdboLoyQEXGcl0Jp1JUb2Tta29etgussSXbviarpqWI4ro7dN
e3d8IJebvhmTN+qt2doLW4qBIyM+yFXu3I+bEKokJrrdS2/GbB6JrqWBYixj7Fit
2KRhHbSfLQejgW+c9KW9b34Y0oerC3WphPly6b3lP+IBJ7afWya/bZtJSVmaxP3o
KYbNtEDbp9D1GKhfUCq4ZG+WmcEHVFubIWPHJmnG+KGHLXo6HIMr9rcSPUo6SbmM
zzWID30IaNbiK4NsUFhorMJ7fkze0PmgNu/kaYGpXh8e6QYoVOb1+QhlazfBdWtt
o9LFqmDOLGu5JrfsjLJSb+ZXJl6/BZxi2SxXapG63VygZaMfNAbTn8G+zq1fuu1x
Djkqgm39rZ3d2lkP1Canc6Pc5vXua8yuVRkFl1Ni1ROoA2S4LPyPXhbw3m4t2z7N
87Hijba8vlTcq1CPESaqRhcSyb+b0MJ1UMmG4qXTcGD1A7+X22lrSxkk5JyFJRlh
dZgkyelPDF0TH0w0CP2yMt0byY60QT0XJNOpzUhgm3ygZuwj3vVv/mTSGiZPQ6yS
LZeXOik7dfhpMopPBng0PAyiGaNXqknznZ7aPC0PjFUOPidCuatF+T8vR9388N57
W9Y0L2pSu67rtAyJZAbWP6mr6iy+cZHtij/a6Onhqrjl49ohJwg8fgYsh4eUFqER
ODScBJsCGbG6LmC7HeH6kgy0/T+3tibrBq/WVBy5DkOir0gcyTdxECnQ1Msqum+a
Z2mPYWJrPaD01Z0A2JDNhxA8aQSZTnxEBEmE52u1WJ/C2voQv9HDn2wzrGVO1H8i
3rEAGd+nIuCWvhYoMceIRprr82anexKCYoQkFFhMHMGAZg2iPQfGhH/B2nVshYaM
y6ggZfvNMS6N/x5av8Ivh2RwAD7O53Pm1+sN0a3j3y2ad9H3OypXrLfJnvrYRCHa
QKvGhJH3fpgfqxri75FoTBLT12BJ2QAB5ldtUataTLxZW0T5XAMn19rWcWr7wK1q
iA5/9bWOMNCy4GPeBKfHQ/nZkGRmU8rWxbRp9lveuLd/PXRV84RXNe9hjJLRSyIi
lZ1xfv1WeLYg3xNZ1z+xyG6p2256lg5sDZwcQKuuYz407QT1r4TqpG78CpZN7OkS
D7EB7qFhrgUrHe/zFiFY8d5rW8YoPgWo0z2YghvNbuHq1wfvsQc2SNB1XPzelAWy
pJIBSTDreeWsODgoLqeljgZapsATGigf+Z2r8i/yOyC3EqJ/WkDGYNgkfB3wUg0X
kzGgiorg8QzvPYjCnMDFIfAI40PlXW59KoqDIowbAzSQT05gDr9dcYmn9Lnnx1LU
P6FiNiCbGG9tmUsOBuKnZr8Hjf/eL9WN0SLU29N3HbiTEofgwfkXA3aSTR51rv20
cfks6Oky8nGs7NnIJ2oLMlX8sv/tRkdNBLc3Uv/NLrzOjBqoNL7CvkdpxIU/S8nD
wErM6BXSTJgHo9OmpwzgnDkFhEQpb0Lv0hu9Y+u7FELB5o92+Juz1577IQ5mFusy
drXKvlVqEiELEG6ZufaimEqH4k5q+bQodYkl+i2l6HSMDji5h4HwCJFdBtbL8Cm7
sawmcmkzS7QE1JoZ3fuYH9EXsJaS8v1oaPopyXCmvXOXUx1kKvG3vV9OtFS7i+Ow
fuVPYZ/uuos6QF5/r/zAXRXcxPOmGRo/+bh+6q6VbgaRgoX/A3fAuct2MnO5I+fe
D1YfnnaxpJazbZT7kPOmaL1I5WOkQpqnyHz/FnH0ZBpVqSuSlgOSL//8whIJgrfZ
8ExraB+pKPn3UZ8L4nI0osiwfXw1sVlOlwjZ812GKBCjmBDQAM/wn34zdkykgL6s
X/qpxsWHBa3AjOs1yo7S8UidNF6b8Upq+1bYb9flo9RdLqvy+lICJ+gfiMGPMo5Y
o5VNqnyHCuq/uJvttk0AkY4o3AELvm0fEpPDhRTmRsN04u6PdD8MdJdguRRtKIxH
LikdH3+/rSgnpE52/gtLErwiemDYv+a6CzqyJ/ICIGIW/Q6Hv6WN5tbqZopPeZy0
ECx68GD+5IWc0FKJSoHPuUHrb0jLjH5SRJzvcMY4f3bEqDDrX7QPejw7uZ4k8mn3
2MSWQSj3Di2Z82RREchmj7PTLVUKaK5Pim4jTTokmyx13IFq4TylJyYn4x5NjCyD
HyzZpFDK2Nliq1N7nRa/ER2R9xDkHZ+r/5jApciO51w/pXOVRayLQxC1Y8DJf1fv
HjoHz75m/aqB2Mp2xXnqwvGOKUlizDGPmb7G6gWZ+hAcNoiebkrRork3R982DkD5
v2XHllxGBYaXI6n0PR9sUa87kHbiGlVuhPa1EQiiAMN1fMCfb+a/aM6GjZ76heNu
j/mibHLyGG3+jVenbmB9qffCJBoPd+0Zgn/eq3HqUNslqUyvBcjqgqY9LdbihsGY
Ye5q5XeTfQcXASK1V4aaSof4QKCyxBU4HEOdNiD2mPjnuK50KN6l3eANTDqaiII6
d310GucP0Nq4D3t2ruoG2WZpQIDqqNMM8DYI4Fk1RlKp/kyWazntSlKIx8KZ6/Kt
zYBBCsmvGOZ+pSKv2jAv2lvg6cTfkmfYwPHxkEaoaWD+WoLawLod0tKWxetK8YCR
ltwwKH38rZxhRif/R0SLdeYq0GDTogQ6YKgiVv5BSH1N9GRMPzxDm4XsS5Z0+pge
2MZE79Z+x/EJ40SlSGYZ5DWLcCQx6CR0ikt7srzMtP4oAparGP3u6cH9V+ZKazOY
zcaI4yDGoJQriSPNQCIsb7/m0TaHKwb71+l3SPGzCFURJjo63om5yexewRuqQb2L
MCHMZY6fCtqTu6Kmyg12MggpKL1Cq60rNBi/fKjao9bgKquNE76esSdTPje1u6ot
arxXghWU3cG0+Xx5VmF4J+ByLMseL/MjSJOgXDQ76C5dJrqTMkVcxNR+taNc8Nej
+kqbhwUm9aG1H2Fhfv3YybCSR1yhK90Qqs00B5mqpo3982OmZJgopdaz9ELQXSix
Vzoyn3yZ4VqkZNyEYriDtbfyagTn9HVZXbnmUrGRQa7lFSWjMlaLQ8PlpwFxxwSl
46+TprAR6aD5NX71nDKQiwODaxKyQ3+e5IguvilKvG3x4gmWBbdHohL1+r6ZIHVk
XkdWeNg97Inm7DzCIE7+QWjFwul7yrGkhNAPY9Q9VHtvo1mN//xgL49Ig02I+aMC
IqM8JmbMdcDfxV+C8YDtMh0hXJboJIMG5BuP/DH+w4P6sdyy/MSAcOfMbwnWr+zl
qE0GL+szQlEFO+1ZhvEm3xFLyfmPZddGHrABcgKJIC4GVrSYcd8B1T8bqNU1W2M8
P7bdsiI8lDen4yMtCXAv2Ql8ce9+ADNF2MAke08a4XU5KzvC6JGumccKSvap+u21
7o+isyPLRW4CQWCMR2zrxLVa/ZPzPWtTrbkb5IogUaWJrasRe+t2iPmmknk+v811
UDg1EKNzMY5IfhUsjUOGraO5uMtaPbhd7e77lA8Lva+SErRqIs5nsFIrmXN9RvN/
oW8nH0cb+tGuTxsX+MuVEdI7U/YjkvSIl3aSw848WpTgdKIzd8dIgYUvbiY9Rsbi
IsvicKD/l28O5jVE8v3u0dM+A4JJF4Tv/cyy/cZLpEmKrx1vm08RqXhbD7taPFby
kBNqWzIIQKbQb2cw63VVTaiZfYT8K6iODbHK5M+231Udevx5rz1a53c8r7WycK5h
QYMaKFMfngZZTWyTphwxkXyHdtD2RyoXYsXT8YkwbAxuokZoQdd6uHbp9AeJ0r+O
Kox3Kr0Dt2nKbuyQFtDrc78nLv2zbyMslbGNhbyIc77pzo3YP5C03L5xrusaXyND
chYb7YOc0Rhf8TOpVTGgNmVtqB6tWLR7qOUP1t2GQ3TWRtIGm2BNLRDBNrYjIPdg
pgfEL9/CFXG0S534XCgEI5u2TUKpNi437jLArLjTZ13IMG58FJXmB15c3R/MXQ5D
jhhdOHYlYKCfzAf98WC7mEEgSnVLNB2F43h18HfVOZT48ALGgMITDQvwn0QB2xaO
KOlchGc8+BH3uSnoDJcuUIbbzTW5KPek1ZDz2I2JGiB/bDUTjxNJpWX0KgTr/mEw
n5NHwBNzUbSwUHJgGJul7QPEVz4ZzTpXY4bRCTISohw4HBd52t7+mHp3nwCQm4sO
K5YX34zdVLPN86acG0jMw0AyQ8BRvc6xJZ04rAUWf7Xu85t1SLoX5A0sY9fdedTG
7bwr9b5kOFUCc8W3YqW1pkaZmIzr4QHFcVA1LdxN29Z+lP673tzqgWq+aqUWsHyj
bEO2ho91MLlDgeeRiDvrXM5T+loLM0+Lb5nbfPriP7KGxHSjJP+Xa/uIfpezKmzl
YdgKHIGnTMdjTMtaImUSALtSK056sbdSl++CfNsvSgTEOZnZE3beD2FXfhRuAIpd
Wx+XaDIYYNCW6919nUGFW3y7oUvB3PZb5CUWYPwd+89EEmkEcNwSI9qaiS5YEF/Z
NSnzymaKC0d6vVmQRUdiLXKagG29z1WT/uKbvm1+y3d+5m3yWxq3BRvV6+wbFUyM
swPSntSCZ7vCNBuyS6ZNGD1xjBKKphob4crNiNufnQc4TpPk9VOvJ8eOckcXgqZF
m/0xTaWIJrdhRNkBr9q1H6o8n6+1MDT0mAUNNZE0ZB8aN1ZM2zzRLr5V6rtaIi44
YibpFx9rpB+vl7QW4rdO10HSBCo+pNS+B8J+vyAE7Vgu9kIHesmYMObZswAzFieF
po3M8oE7Xum+oUz2r9FCjG1Ij+Hxe+QS9Lk2LSKqMgKCaLiWUAizY2f/kepbRKX1
IAgPta+R+pdZkv7zQxcz/ijtQkl14hVP1b0XnARRYnMoxFOGHPYDnGY2G7Zrw33T
ZrFU2TmRNcPBcqxcyVTiEDs1P4DR6O6OxsuTvsHZltQTebNqeIeVzziMzb9egAsq
Mx5nFLyl3WktmNEx33BL4pz6vRJwHiOxSmzr2NTpgjXGc6tVVQpzN+H067tvpIKp
ZZov8SJnv46PZwBqofAMI+tzdv9nmo7GyuWhoYTWCUAonC+86EXjd/oNZ3p19016
O4L6nklPaty8LYqSDmoIc/FVexma4IDZUbma7IPlLaoVrw36j4IlLYKO7mExvkxX
t8bqaQtZJvO5hmNwELIy5ZYvu8NYme8g1qJcGBz14Yt4yUyfg94M3MSnUAAEN8eJ
bKv+VJxmzOMskY/gwnI6cJjPXt2DdMWYUODyq5WTeozUqwgClnYYcbLmnkg6UtHt
8HMATq9ekSjbCM7a9nwIjTnfJOsMSAQDqC6kPmpyKVjrBg425+HuWcdy+CFdH6++
/o94cInPdiK5gLNAITnQRqM5NNFklihQV4Lwer8L66mlxxkukWR9Y917HflGsxw1
sbrI0f6hGnjRLhXEOTA8w9RCopeEbKlhQW46JsMAxO5Mq9+hbHVXJhTUnaHvUCH4
rjgaWquawlyItcOz4fs/5m8VJn4gb61YY/nHyvk8OYdSgwh9ig2NbTUOPtM6pENu
P63zWDf4LQ190dErdU2/zwdzXbblagU1JU7BAkzP1nCbDqvdjEQhzzXwIeWvUYmf
a6IjmAf8sZ8GU5MKViZizD1cWcoWWSBHOqcl4La8UpHEt3dCV1OOTg4PW0WfcQkn
w9vGU5K4bSllflmMqX8dXDSWjjS0KokCjkD6uwEWgyx4SVhOP4uLGSVPO/rIyaxP
izGeRx17f+z2K4jFpaXTHQZTtoVB6v/ZvE4WzqqY8Oy95uPO49Mhidfyk6m9H4Ua
tM5ac2XGUgUPzNuo81pPODWbYyH0YrG0OqVJ6HkgD9PqXD2JXq1ck1godkSvBrDU
pXRHk1Jhk8fGUu150puzryi9hUF86qUzzVIYQYGVU5fXcX+9fMe7yC+O2ulslsLW
JCkHnDkdGrIMW0KMHzo6WmYqDTszbEAeIeV2E7GC5FF7lMCGKBuWzSMLOeSGo5Me
W4Lvr8KxTmugfkDyZEGnGZ6d/ijj44Mw7poQYSYAxgtnuESa8IMyvdIcQfHCE1EU
oMF0sJdGWnNyPsEXu7UFYo0RYMNr9x5wj0mu5KZCnpl2XvdQZKNzJcKkpimSn3HH
193hznVdx3Xtj/eur0Ycgen+k/he0/ITVvjwCyPVNKrIVVeBSzHr7z1wKYpTdpwv
3hV+G91uEA3bjwPmi3HzprmzSVeHBqxu/lj70uwdttCKn5S9L7RIrZB1m6ezhdcA
Ktyi/KjGDU2/lQAu3nDzq2b0fwh3z4ZB+y0HEoEo9aNFBCviYDLoOvumsfUayJG5
poYHgFbwkRsoN3ZqSMLH4lD/h+N+iqUJtKAZPjlPopfJIxCgpfdQToQzn7/F0Dbx
tctxhgpovu0wA87TMovdsknxzYt1z4wwPWss+PdlrRWefJOi2ESBdL04K1/DzIEh
/2Sok5eFwdwJS4o6MNtav+Gd1bbhxfNoHDFLOFe0vIqpidiDiJnBpQBfByYrBUID
Mi8qo55fWO9HsiSKR5PV1lfh8dlqEcmczdiPHDeyVZOWP/uGmdM988styZzXLHQk
3PKL8SukdllxZ6LX5ys9eSF7c4raPSAG3eqKdiOKEgdm+roTiGGkCpIJZHdhFrpW
+sZ/swSKkDpvyH/ZJSDq05Ea11H8kWAwwIz1M/Oo0H0P3dd6Qzs+IwGUyb8VELCg
P2NB3CVny/+PUUAhNQtRcrAQ1ycWapZQwsTUTwjlqVJhiNiF2dQmQfc3eGXSxxqS
YUWZAq+X0BGLngP3Nq3NFkwskTtepWDUXbBTHtSHvEZ2bOiZgU/P8wxJC6B9lOzi
Y30ZSO5MsruYc1cOlv1n3JdUaRZZBw75VxjHnVAYZuxHQwOsDlL2eakiBOJmwQZR
tFzkNihwyU4IuJRyPkzSzBxJFVVOhLaqGAR/Ud5Yta1U3IkFf+NgUSju7QpAvMNp
d3Inx0ala4YbVepZVkqi16DxYZcokVVLJnUCv8dVIpOZJQ4VthVxWPKhUdYCJI6g
D6qXrlomhKjocwweYCCtPAnP132JdbV889V9kxXDE2zjyJBQ5iq5rdxr/9tNBUqz
n6MvA6gfCsFhmr4396JhrYlBU0QYLdSwobzXCgF5thNwiYfBKyAKRmyd4kRvBsrz
1e6eTJ4xc1blkjGHSAPEGh8G5ceqFNRsOE6D3oG44VWEEA7g/vJ7zWJcg20fCqoo
KaTnLM8lY6RsHw07SdsMWQPfOnBgXXWwCU1G/E7rgIf35gk7dNt/twXkDxoLv445
CUilSgPloZon3SugJ+wIT86APXfTLBZPCFOs7DNUFhRC8wdtaNLqwkekEqGMagVl
ckBHIeeY6UFXIqfZdAkdEmsOnflSDjY1XSd2eZ52/GTmyxQHxCM2wW+ey6DsC3JD
+XfEJck4iy5+27DIUg0/NqLKMoJyvGIic7W8wNKAs986a4vC6imxtDF3n27P4rAc
rF4jtbeptMw8ssCEcPAfSk80c9uU0tr7b7slpfaEpeDn+afXwNHHzOCuEiKwouVE
G6mFNKmv0PL6XV+emZ0awiRfXM23Y0gR91t/YGoRE9XtNFKbd2yIswWhHEkl/j9x
JyOXhw1KDzsEzoreDEU+SmqAa3qGz6ETNUFpS8N5qePk3B8R0bv0c9aNNSSCSRPk
rNDr1VGNidnb3LNhivXS4kJEGL2rXDYeJdNetgnlKXt/6G2VHZZn3BPQSw2sw4PR
+XHP4wVjlkPGJdiVDnuw6bzqRM8BZNaQMXiQVWOO7u3CVKRwz2AWCReR3Ghtu9Cc
O80vVTYet+fsKPAD22vdDz7hXEdkAnJb6Qe8sREum6NLP+mO015EizjWLKSWbnDL
LpsZyvy2w8pXbtRsiKYTsmjV+kg/g5/wapBSDXpgJaU1BtXk0sbD4zggiJQgOf0y
K9xx2AaxYgvipiNFCNFOzyUOYD97ERoktjwGacyiGf9SWEPnpGGm215MGCurhM32
xtB51T5mA/BUPHwMsV16IyndzvY4trOWGotx7v1fD1ZQdPRQyxMDU3QZ2S9pOdBO
ToZOv4JNv4sTriRnxS0g96JaPVbLoEMX6k7YOftj/I2VSCk82g1JjLtSxxw4QwwF
qIT1lpeC9NIuamXViw/hvwz1cshWshKyLJdDrm9ZXtqxNnZVQ0svbrhdCNpmH22X
JOycMDmR8VQgY0lr1cPRVP9fUeZth7jE3zX3JB7KqkFc9pd1yeNuy3nexZRhqYyG
Tb19Q+FWfXg6NakYxzurIEbEOxrU9MTPXDjUlB3mfTZ1ds75k693ZZnTWloYu6es
RjNnQ+VtqqlCwL72VELp0Cgst2g2emX7RfaR2mEaafKXcx7YcJUau5cy5sJ7v96J
UfUZzw5SOhWW0zLORHVjIsCRoK8XsiGxZwGHvhvBwDHfqEe57CVe94XtoSULeK3M
TI4RcaGPsQ6LcxCm9xZs0oogzkXbHuDUwYiS7H5Ee4MBYgJFBirpyybLh+c/yyCd
ndmdtp1+03ECkN58kQgUjTuBbP/xnwhLPDXrhaQphbJieeCbn6K2AQfkH3PdEMTb
AsytdsU2ikgwHrhMVLmrhOzt/AS9j9Ya42CmY48T8vQI31CRBTrl4RuhMNo/06SQ
9RKzp4g+DXFE2cNcPmw1DEnr3hYgaMZl6NUnD6SqenDLyXdYImZ+eE4C91k37BQZ
FRmGtBkzYXMw4S/xlTZFS+y71ceLKGd80Tw/Gj5UPuJVILJx7yw9j0wCXi+BZbt8
SsRjqxlhT1ojtbDER2zINbJlWdi9F/kS2/cVffHp4zF421pWOuwxN9MYBfu5PMId
RZFY1oEqAEXAv6ldW++jITeAJ1NFMVMwP0posEVdZtTJZyWZRoDbGWQjWEj2W6gl
okOyPQy5G4PlpnFYZ+Zlctoj2wuNnylK7MdJb+CKnrViLeZ13uJwuNZvK6ke/HOe
KcczZey8oxl9MvRYbrdTbkyuumWy6EgxYih59vFntpnGx5BL9cB2kKQfsruFA5Tk
gsHKfmdEQMXulgxG5+vdfK2K7OShrjnhWInzBH7wnGeeyz0fI9Zj9KnBZfozySxR
lE83fHo/Zy2hi7XKZwswv3EXt+SBwo/MkaEjjeApZMxuov2WU2UazPKtIHIGqScu
maRSK+jh4Ep+/Sofc/5bAgFPeWMy9yDNfNz72oHgFYodr0cBEwx02PeEAd/j4CJi
hs7v6PX2c4yNhfKXVnISnQY/lF50robCKc7StStabhhtsS9vub9BdcNjUFqXjf1a
2iR5o4jLrOtekF0Dt9hDx10C0IfkWWgzze9sMaQwNIFno6bfrpZOVidM7TJjWpYq
LuJCYe7Jb612aUpmML8UluyTdsj/Z9+aJQbw8QABEgqAm0lXgO1uEmlKgWBQDs4F
MFTDhVZhjWNfFjm+wYssLimB94/7bUqchwGr3DQP6hbjmjTODwEfH3nnG18zJTO9
Skqw4YFasJcrXEKXHH8Lmc6iFZIadZ4gOA4fhJ3F6s8lw03Du66hxW4wRZ6aZIVq
L+6+K/4xrYy7ux/BJyP98B2gh1UwBp7DDJZYpt6kvuKPXisfPBOE05gsKQhU3Qii
ISQryBle0dnJPPp4ChJk0a0aTEmiKBfBRfquojM08n8mXGfmX7QwfTONzCqAFpD7
JcZvUY5gfmHYog13cj3zCXnDfWkkaW3F1FmSdoEkbFIkNb9GXvNlblk+xt46EjEU
NW/Xja+DCa6QJTFJv6tRmVzL2qEYbPSaHY9/c4iA4bRnOZlOIiX36YQIB+09QNiX
kYiVq45TbwVNyAg65bldI8SD+mEjdIvvNv2jEPjz1hm9l+P3lzkzo1PThY/cw4/a
GthUOk2yaMdrDz4KD8AnPtmZ9JJsbcdQL0mxSJr6UiQ0659lyxLAlEZpS8azaFzh
uNYSAPojK53b9GTKpAxRKrOxzG1KTtK3erNMhd/d67QHo80LxWWo8gtKoYgBAMGo
QEKzr9cnh7Wy3XP64+YSsZT9At6KuwdUOhpYmEtZguayBAVB3CkmsAklUHF1ysl/
NNx5IOhotlHNSRLSOe3HOj3/0hzfleHS8Lxs09ioj+ehejetvAc7MmRrG/xnIDQw
U1eW7UC7tJzUSuB+CxFAkfxcwgMAA55q8DcpoSI7NsgDC29jIEa7sy9XwhYvd08w
vG0TVGgy6YXW6tTQRGeFeMYxglWNfEJb4n3ye4uIc0ZrlUXDl/DVTbuVCgY05tLQ
uNK84NRnnppepJTIPZ40n/ATA+WeJq2k0FhK8T9IOFjgNmXhn/47a8jpZFqlTdR8
zdVppaxeX4ESJaGB2dbc4bNisUWkwMAytdeK2l3dGhazuuAeBA5yEaJOm8G01ZxB
RPCmrzhRnd3ixRtD4TYo7JKvA+NCgun3A3VVKMBO8pN32TDvFau9uar+YyhQ4+nf
XR2/rX8HFWXBTEo8oAKuvI6pIm8nr58zzEp8oDBnESdJyM0zUBxYyZ1OxpSzo//v
ZTMyHhqDgUYk6ookyNjvuTRxWukjq+Cu6hFPfsYwqrKXFpWNfukoSWlze0Dg1ci0
xDRBouEBSI44+2hfSAVLH5aWQwOG41UA6JwDgTikwb0NN7rySzmLQ1CE78pKa7/W
hgKumdTWSqX4zxprifL6M+r6cLEUMISk0Dckg4xeroT2ZXYxcns+qxwD+nyqaIlD
hHGxFgPXkM/6fTZbT4h8tyEKa7HDy4UhzJTxJGVfTxfoiVIEoM4YSyQ3Lg/jfGUq
bXRC/wCHUVgH3SWw0w9OqlvSFsP4AXyEI0ORa0T0ZRQgE7bPLHverWa5Q0rHKnST
H3koeuSRUw477oehqDXmfph2PdJhU2PAQfPMpLlAQ940/Vj8m9mlnSRCQ9ntL7VA
TE0djfRGZ+y5AuWN8enpynSR0n/Es3mxuZZNchLrfbeaNkztX7gicmUrvLyQ3Ur7
y2m9lkbBkDJlZjsbO2D2GWgVSrDJ5y9ELd3rgaCQ4c+DkLKKH6XNd+8JB1s5TYp9
59kRNtB6gL20rGimsVPyJ+wqw3OIyz+hik8Y/q1wnC8kwwb8h5GpZ14mMtlUIcnZ
qZT+P5OcD28dZSLdUswTI2aXqc4aJnPAzt8INeUtGY5y/X3lHt2J/xGV2cBOq5ci
BqzGnpz1YT5vb02lKRypOGBqdMBPwLI00Y412RivcC8RbjANuaE7a95+3sT/LHJb
cw/fJWFaOoOqU/KjHOH+NA8eEpkImwMmQtyc6IV2jenDzxXmfUy00FOsEjQimiaO
XCN/3Z3S+vKmb3j7n+N/3omFPUcVxm0wF642fwIftegp1mC7GTQyLOi7HuLOy+BO
faALlhihKQyECHMsrPPaaKGTVWSfCdpj9YiEYQOJ72jZq91BhHh6ie3YwriQz5F7
c8Uq83dCwm/MWmER7kWSIW5dq3SbtY0jSRWEgEC+ztzf73b9hOStJDkz1cuchme+
RDGDg1tz7CL/D3lCkpHI10riURKMM06qMcGEV75LmydE/zc4W9wjM9QxCM/HmPjq
RQz9cBTO8YZuXRQ8pgQTNA2A8CKP5CWkMnmWrd4DIbDUXgTdU+5TaMYJ9TlYY6qa
o1HeiLbwHdGX+cb9ARjuP7oERA483Scm+zFEL1kHLbJ86Nsd739Ew3WJ25RhYC+y
qzXAeOnICSjG25PkeZLff3CbJJUIt3hJ/JgyQjKmNdytGvNjHGfx8KoF6Y+IIfu5
z70EQCBNqbLTePb+TRK8IjY2NbCqF2j8E4YMOO3MGqOFEPLduzyR1kSBxn3n1QoH
J6DgjT2tebq9UzLBgUaF7OM3kxRwwOzWG7wF2Q4t6AS6nxp4TYqFupQNhYLHhrii
Z/8j+GumTyQFLgSxboWqD09P/1r7TFXfefw5rzzWA+JXKLpe3QZcXxc8/5l4ss+j
S7YNY+bEjYYMIPG9RM/eid+DcdejLHEdeFK0mdlCPjeUfbXthvkYuBnDhRtCWVcx
jOJ/9CbChDEXGB5Ns8Aw5+io5KOIMr3UPAL+X2Zs0AUByTbbyeLvUVVzLj7ABplx
nIF62f687WNVm4So4a9NtWAE1ZA855U0A9yCsfx8Nwgpn5bWAu6D0F0xVKhvZkbR
ZRu/kRJTzKVMWHEsmnpWHuTrY5uKTEWMT72dX1RjkWb5Dou8UHvVLhjaXZLLsO58
yiiyJTSKNoDxElGCkSP82k8I+2XHXSdKjGFhfKBh04DLVyMt9Oom0rEkGl57F0Sg
6lwxChpb92KCyVpTNLSmqaPbHFgRqTzKyYyi8R1WbGndnf9KDh3VP9cfr8C/pYuL
oVHb5OhVY/kXXZ63vuY8hMAvtZw+Jby87P1O7D9vYC5Y15pBBvl2uewLi/WuruhF
2VIybE3X9ApOazoj0yDfJQeg57kGI91AvAUSwn/42XIaXPup8Q1QhaglrZEiWgMU
wGGhv0mFVbKizd7vRSnuC+7X+wRS8GKROlfBl/fMlVfpreZhINWa1di7xGq3dabC
BQINrWKbp/0pPkjBH0QTRMouHz74VtwRVacPKTT0UxZT3yZwCSFS6vXoBnsHypQb
2knij7vjhl7QpicPj7eBZZwaXHIxGvqmAwORiLmwppXN7aUl04GPGNfyyQkcLOEA
9PPeWGAD9Cfxnta8ACSY5UdwUXO68vnPFNffvxDFpwMEnXsu7J9Za90rM5tBLIhW
g0KQRkKZ0eY1R8CSN1W3VKG9E64gFNi2RLgIQFpuMniHLJXZKDxftq1s2EAibBSU
l/Egs3O7826wJPrdwR9FDLsWNUnKFKhXal5ZwB5il9zsXSU8Eq8IxDrgYlWyOAV6
Z5ostCFWfO0rCbp3z6ZietJdXX/iTFYy95guNf3mB3MYUS5NMEhPgYGn+kb9OILN
`pragma protect end_protected
