// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:45 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pIU63A6B+nPHlPiVTH7rNLGMMLH8tfvTbA7Dskz04zJcKjMOpCWpizOlehBFWdL+
HouC/CHzOtm8yeN3EfClsxpaE+blpD/eTIOmyydrqXhfQ1kzpDy3gdKgu9OH8gvd
YqLU6n20bTfRDdL4TwpuYAFcoNVP2Nsd8lFDRLpGjCk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48608)
hlfwt3ANDeI0lejtnIbqu2HbvggijsfC3VaTQPp6KuYgnbeHVQnNX/LOE2uJf1Jr
oLfC9T/9nqjTJXMEBhZE/pJKdw7UIuhAvLeF+SkOVMTKcTu4n4MEyYegdHafk+hR
IXyAbu+Kj2ufGRQ55dfA0KNQa43keim43ibWCxwe0X7q5ffz1uLJvta5MNeMfF94
NKQxHHQ7lwi4oyuVeKtrF4n0nssFzs3gdSjpIFBggC61Wl4bjqlk7TQSuLgRu4wr
u7zzFhktq1QagW+HNCZBgt9hFsSoMFkS2Dlo906H1OJtz+/8TGVnJAceVA+AAwi8
5g9G4euGg8FHVvWfxionLIe7T3/ul67Th6BzkF6rTVzSmI2IQjLD7JogCiGQzWFt
dAMBNFbpou5liRpuCXwAyqFkchfh9BlBiLxND0QbEa5QqCAebfAe6JIhPSawZxWO
S811+Ra+GRvol+SHD1gKVezmihh8kl30jZTHuxMf2qpHG+FABk6ZLQY8NidzYmOw
YNC+MKkcS77cnBKJRoO5yFpBi4IwqJClFOhMV0S8Rbtf3DFyVlRlOQxF1J4yj3fp
l8xRiLZBOb4NVqh4Gd1piq4UNyxy1KjYkNMIoo8nelkuUl8nGUcsxMwe2oTh5xnM
30i7y+0MJSHNEdKAgIaHEYUrMeXd8Zp2C6yVXxh7OXRaSY3OoymR6EC/+bIrKECW
GYcwuX34gc6W4tBHijbAY60Z5VBjGLKEc9t3Jh9X2RmFqqzq7AZKBGNphEnFfgRg
q0XGkCFTcKxQDVWtJ/md7Qu+Yw3x6CFwhPLwj0nw2mUp7gPRA7F9W2A3p2PsNc3I
Zcj8zypC1vFzDJ5YrbxNuoGw2QJkQiZIvdDhpoUPbo5mdNrtywlhcay+FBpCab36
bw7x2x+zwWFtURdyEGSGvsmsoE518SD2ScjkFTvXsBUyjFjv9VduRn6auBmXH7/9
KCquyDvIBFKwVujF/o2AIenIvx3XoKXMtXA7fk0zYnaW4LWoHc8FjFl6Be9andR/
NYaV4pMniHaEvHWL0ljHwaS8dXSZ/oG0vteyA4yC3QYYVZ0GUKqpdut5suVKqux9
0/ACafm4WjwvLYnVukkYX+0YufKxsP3b6rLTn5Ccqs5G682c7zreUrsScmoTdmEX
Rm+TjElIc3qOvd793CKW0anbQ72Gkc5h4yQ4BbPkv1pzvbMuuw7EphMKCAM37TpS
8a4Ev4iQUpm9SXCF3jvqAhhnFPugzaYNi43fuARIqhV1TujLaaWEoAjWHrSaXvFC
/il1TXcBqwCHNYQCD0kwgDvqpi6hPRtwi0/ehskl/qffN6ESIDNegMTWdl+4i5D0
w5DcX2x2agveYLPYTeQc/YtNRgiFM93BIjHC5gekQs49rO6ni8DXfG9YLadlehTL
PF40veInCYnp+eMd2HIh8qhB9SRBYX03M2yVUBGmZI57a4W4lH9DqnLoFVhrPA1A
WMdr9QqkLarxfQH2WgBUdLKKRZ5zHpiulbgU7+wn8jeGBblU0+QVOv9RZU4a7cE0
wbbPIc3k4PWJUWRfvQaMYRgoZzWuRcxUTnap85Tzs3GEHdbiPCcScx+6wbi8nH6N
ipuH1d7qs2v79KL6IMo3H6a2S2XjFdxMpX/2bNHewGE1n2j9VDiETWM530AUYBk/
rJJI7iPbxlVuV851XB7Fc5J9gn4q3s77RKBV4C/S1fCuXsnWP1095vRuFZzEGoje
oTP5xV98MVDpLsIe6UDDwrb52faq3KqljqttoUdEZGGjWVJpA1brC6sf/FNDIKSP
nvsKAdoHAsW2XMeLSUZZP85755TKQE6gOZ6xOr3LZMGHk7bG86VwC9Odv4F1H8+A
J4m50YM936LcpVyuCRFOwxzWc3p4GzW087+uqB6IPs+pUWc5ppB3ehzW0JjoSglp
yNNgm4mzB1ns9CVUNb+pFUkVNunvexlZSOhAqUioLfyYpMxlfGOWmKBX8CrbXdTq
Ow9c7DnXZBde1RqBXCndQuFP49xo88xzYFvVP9RrGsTkUFobvQJbewMoja09fXPx
k9wfewVugIjWr9ghQ1fdwL8TEqC1S7P8CYSRJEj+B6DvSNCYy767ic1Y9mLLJOeu
xNGHG5n7TF68ll2TmdUIeD0tOEnZkodvGpk/LZx8eL+40u7PxKxYb76qRokD7mYW
pLctOPHv3Dcv4Pm7Lz0IB37cNGE00Y39f5Kdq/XMw8Eol9cNk1dQ+z3IEs4pBJwC
tOnctWVAkU4bnGzBVNhs9TlaEOZtZnvfPVJiTifdKd8q9OzOMAF6YeoACslbXnUb
MbJ6vZjBVtdC176CxvAE1aJ4t9WyfyCZpFE0tj3rTfSZfWJo6wWtsDCna1x/rDQI
2YAmh7mBNbITXXQ2B0Immi/XFrh95nvFZLxnI81MskKgynXfsEz7MuIcwYzr40RZ
djO3Mnq92FU+lFjqeq/3r8QLU3/UxPkkecCUTPEyOKHeMLnwSGu2TCqc2pQeMt1M
hQUA8IncJT5oce1Qjy9ezjz83UCWz+3uTd5ygIk6jTZoHL9Hr8IuFvNwKGjEVXyM
vcnQx4Uf3LatlbGdBXPx7WkI7C64vlel+cMV6qWFUQs7xDIF6/0ZqH6KHrZDmiOh
7bfcWi7wxNs907nH7oQwRlXggPKNcr8j5R4dcqG/8j1fIdZ2jPyvuxStkaF1ggPh
8cho0CjTfT0ikS/sh6ijiFZCdI0uLo7jb7DWtGaeF0vim/vagoSJx76CTl/PjxmM
2spAZsxogdnBEeXY5v8TuokBRe+gwu1E6QftMPvtNISVOkTZneiBIQe/4hFqdrQ3
zQxGuIjnh8OWckO0ehD9+HGjSlIav9RFuVPsx8Hv/QzQrAMhF2nObQsjxcoL2Qce
nnx5zbt68B6BWaDVM4+XFx5v+kRxugEhZPMjVN9vk0g4jspkRwfZsBud6I6JfNcA
thlzng1QoTYh3AjTzPFSAzJYcCM7ZdXssqVIONXev/BHsE9XeOagHlXJz+T9sgky
ZxarBOiRlMLZ9T95NZaTbR0eOX5dMDiKtUlE3KqpG87hIjYHfXNi/28OXYnE+fWK
jaCDx+XMf/fEe1IfQEsXwEI/qpEVjCtiZnNDk78zCMp5ZNjjq4MKOc5Rea7gGIWy
DfbFwwIaQGhEw5tGae+2yjxuUcD90rlkj5mDiZLhIh+/RXXrusSAIMVl+jRgU+ve
pagocJh+ivFbxcL+z06xUx6XzUkupl2SbT1nz2PYqIxWHMnX+CbWU91ZVJKa+Bgf
Wz4KS8tVg3Lk4ULC9N5GbJmNJwdkT4dmdcsIzfB+O9fZ2vnSYUKLThAFEIn72oHV
SfMfPD09WiyDPg7VV3e8E4yVeWFxto9D3wB/QzGuXa/pMncXFUfHqNCjBpL30V4+
mvrdbYd4ZHw9SMsirXyyHQOt+8xlA23GEflbn4OgxKLBVNijYxcFiydT/7eItmgO
TCJ132NuQaYVrkAgv1Tjt2iAFoqXoy1I9k710n08PvOcD32c5t0+Zr8Vy6A/FiLO
ZfyCNvkNBMrS4GzvCvNpAR9GAOd2uAcqVeNnNyBr0+40T6mX8odZfXvsbFmKtrGh
lZXTWtLvmwjvZSj4HzSDBH4YNZ4p4msmVC5fR5Cmy8f49rGt5RdqRGs+CJAdcR7u
DPdOIzOHniiqcqra2lOx/h0tDqS7gYTUOlc7RTjkb991lk4OF+ka3gJXLpOZQv2e
+mZ+uTQDAh0KdRcO8XE47iAUE/+zy8uHFB8oTVkh9F/JTsFtzOFo9fQXnrLz2/49
WGQj9Zag9HU/S6vmu0N1YRRlzldDP4EE5NNLMD1nvt6C+9H00wjt7Lr/CEX2E99l
xEGeObpO2CDMC2R9f6GmaGcyGkf6KxthGI66Qq5LcE/xlfiu7m7QUUj/emj68etv
NrSw1PNIT/KOhHZnEURwkmM898Yu4v0Dxm9sKKSIzTg94+CFPVn9CV4s9xKcdex/
i6TpSfPYu9JkoS7L4K/uNZfd9gKScWhV/pD5DYV8avODSrEAxktWqrGvHFlUo4k/
9qUf0LSvGQXHI7lE9GcrVGvRbF5RmM8yYvXr1Lupnb7FBMxfL6TGq+nIPZ+V+Ew0
2mIDJ4m9i05yxr0XIGyeGvXFKZnQNm69/GG/Jx+tXhiqmc31d8zp2L2xrHRcnzxu
bNlXBsPa4USQ0Z8/2FmJu+dqEqIWzKBZRSxaecWCvxLELa5blPOSpnRf8jSDh9Un
68ckNWPqcMMV3CttD8F+37auizoVB5NR8RP7tO8ZII40AGfuZiuV1wAErPV4LWa1
yq0K9laQhAYHThV9BfHrFGww7gb+c+H2Phblz9khyCfcR5LsEOhwgNsKuaykrYqV
Hgl8lo8ImFARqHL3m0QISDGLW5oWuuASBcc7YHxoq3TWU+w+ET0m65jq+HGjLRa8
RefZWOWIPEf9SQS9gU+RtU8iUUbq993AJzya9Zj3esasoQmyykjjU0dWRMlMWGNH
KQKloNUPxyX0BZOGllVWy6kyfsJ3tGERwsI21hxhXKMPjbjL+GjOJks7mHX05GM6
vWTam25U3cNOZgHszvLlhE3pa/Oy+BDrObDKoEzWf4wbyQ18FbDv6h/0mraQRsy/
p1Q6USpissAqNfBjrqn2ybKipr9xTEzuqDuavnZKqr6IdzlYhnnsZpsTNVk3KImu
rMB65utb12SaLUfvs9aQFc52ReWPEz2S0+xTali9IdULjqOtCwjY42CNkrswX4jF
qcjWr/i6x6PZ4vRWpOaQtDvJa/xCZszOtiGLV9G08zn5UA5Nf2CAvJQwxrhtAiru
the8E5SiY/5Wv7vBzrd57dhrIMmdvNeNhXLTpZ7Xavli1Ea9eOubjaxXXLwssDoR
zo9ueAtY1TlLNOumaQxk4XEANalm0FtDz1Ua5Sq4jZ866Trwjl3AMBpz3GUwiw4t
Ovg8L9lBwcwRVOTpZQ9N0z5r8th/WAFEOg4+sTQHRjV2BBKSgWsoGIO6kTIOIiXb
b80GMTdrzvtQGpGNtpeJG88hLaEPT609r3JwEd05Ow97JdqVk3jfiT4QejgDzSAK
sJSbAOhmgqnWV/oFCwRC7B2b8/NFQ9QHnDf/v0F0JAPBwABSPZdWJFTsA8zRvtIN
CJfX9IHyEtzZrzD+kFYPoZApRNUfS6D4uY9CakSIcqQRxJofYy0q3wAIMTAY31OS
bVsdMDbyNlzt8oKRVZU16Tki9zw8V4TsetxCsA+r1J7sPU95EFhB59jE1S4Ob1PL
qFVgC+Wi71yNGWvg981Cl5q3546ayw6keWV5FYnY1sc0HBEHPWh0fLDGqoPrTlxT
1LgB+muGRstHUZ+4nY6e4zaksxaDy2nekc6FPIfV4a9h61JKOwpvseFnxhw1SKfC
r1FXEz09FNWVmL3VBDi4F1gkoGp/WcBoMhuCZL6IvpdCnfODwae++Y3gHgG6SmiO
0JHNicYS7UkSkeI7GU7FVKXJ7+ioFQ8aTik4VecxTOx7E8YC9SCEhI0zAdUnBh26
lAgMSn85VCZajr4J5/VWAQedzN8Hk8Qxx7IetP08Xk+Fm8kV0BGd+poooS+IvFqX
rEYNwNPYMDuOWFkFZ+GMb/fpXAafoIzCbIjggDP3RVOl/PKQvXhk8w84NYd4o2vB
B0CFJONddEqF6v8mbF9IWtEiZr/o0+Cb+p7EqWg5FE10ZHLYdS5yHs98WfaHHCF6
pYNLhlRvJHGll9tJFF6UpgKo2pSAveFtVqnWBy7NoR8e5Qg1XqAaRJ5/dYgkux1w
av2ejjvHzgpoNMOgIuuZjHDwIz5n4pfIwrnJ+xnSsXPjvMRvDu05o05eJ0L5l+1c
fVIenhnJWclFYQZvFguNyndpb/QpvLYZWl6AvKhKtlMtxnz4HezumzXnVpg6t9Bc
pyrPYyYgdUZVrVJr4IxYYRArPQvw41e/qaY/o2ngwxOga85QMyd82wCSf8xngn1Q
anwjJvpOHw9sCCrkWIBqqDvp9mE+CX6xWwl/n6N0HVR9lMh8fG/nO0QikvXH/2r2
Zt5W4jS4Fmj/ecfCtrxzB5DpqHww4odXkqkvjhGo5FKZXVUK23ImqPcJbEh65olJ
uKrTk7Er9PB5KnHUSKmjeEx0gD6CUr3cjA4dh6smGrQXaoLL9GXWTxFHRuaNZ/NJ
fvNJuS8oOB8MheOYCAK3wk7lTLemP7MHiSMM7Fbo+k1goH9PtM4lIhs1qP9TeZ4b
36COuebl3aoleWcAB+IKKOoD8/iBfeHz2wD3wNzDUggR2G6cYsphYOTGlRGJ5v+Q
6ozzNil90F3AkxY0hHNUP/RfrJzFiLLUAQGHqhS5h2lwq5im9TPOdP32aKoCzfqz
qmAiET8mo87EKgiOAsz9GiGGLDnkJJ2crOWM9Tlo4/NEZpPzQ1wu6mR+xjk4ca0E
D37Mt0rJV8zANq6wiLhyp2M5o5x14NSGrB3Zd0k+/0OGNn/rR7+YOWw1Xu4/NNl1
TfBZSBwbgJe6V1dtcjCByyrEnU00ZTU+mDKnlESaXy2NkErFmAP0NjjvvZ1T2CxJ
Xib6AkvziE6h0D5fZBoxyhCZuBO6xvQDsmX1eIRY/0Lkw6fNiZpU4FGl3S7aDys4
4zz4N5xq49aDMXIaLFd2pt4GN5XYnD0i+ne4LBjBkPVGmNftXIvh3ZHqQRDn7t5Y
Qq4ALxz5ZSILx0MHNR4OKr4QTEaDMMyFKM6r+6PSPW08+KRyfTv6ElA+0op/Kjy+
wEXek2adsckpyJkweVCuTJc/g5ksYFCECgbef6go9BrMRjPtRFTlzBrtZv/V7cW7
xah7nTV/tJGQHPLXRwcPciD2aSe+pXvKJKXhnlUvWZ3FWFuEUu/KiLZnbyDFHzLy
tXmbGpQx2HGXdHlRjhVNWGUViK3KgENGn651vZxb9TTAF7rGQdKEpbakV0nkEXCV
ttFm97N5Zgy22Pnp/fKOXi0KNxECiqDUID/5MwOhQHQ52VZ0pcglQ1757KAHg5S9
H/0QfFcQ0YUwUMbBxwzVL0LL2QL3r1eRS8W3AzW8Bl+v+DVG21hbNFKMZuqXDJdu
o0bNPEGvSht6G/nDHA2PJQsX/nzLoMR28ZZuWB6SRBMcJYHI6QljN3C7XiDrUqAc
/0YuiuLNH6XxRnh9i4aHL68Pe6E4M2gkPlTKniJEn65IrNQgLr1PwkXiob4e0EX1
8JDyoUYnI/LRs6kCnZk29G2WB5uSWymDWcaBL7JpVk/ipseJhlfCcvspL/uPRNQx
zFyxzy+64PPpVrGEnRjwtb9OK/4edKJQY6en/nedllu183hSE2LFrHLkjtKhFfvo
ZVNSN+Alqw8Y5O7FRC2jIMPIzmyPoxKMKAHhfSbRboJslyQ1mtyCmMtdnjovZBm8
v3GuVEZeM4viQ5gwpFobUpATcpldC+oRGfAYuEzy0SaIHmdeQywcyMi5jGbsRTuA
lEpyohTPbNeTjkCIJDE01LMf+1fAy6Q2ha++zMusiBg4s4AWrVrKNWRK732QJLVX
NS5dtfkDMQ2RpT5LncwkHEmE85AeEhMjacP14Q+zQ0UcfUekg0zTFYflYKYcONwE
fXJX/AAfLDNSA0FjMYB4NCHwSu2EdIh2kpol80lmggdOqGl2zqiJllpELHMY8v58
5SWnTt4R+Odid6U+X5kyOai8/8Z2WF2+ctGuIHLJnA9oNXxVs9myrXQMKyXQEYiJ
L0+qDJDT7dg+eT253Afju6ZRMHpxPJfKayTZNHoCci3IpeXJS/nn7oagLStrJIFw
Kozi25eTx2g8z4UMyyvK8R/CsobD7okwl1EhTcMa+3hZCJOXaD204M5vlOXYZAI3
M7J/5lKKFxh+eNzLR3r/MFmuF9uPKKjU4yyXLxRxLU94gSOLUbVA2a4xEzKYzAcf
1SUijrU63UIdBsVHPNwtuRnnhBvVXbGkDmTESFcBKdmnf8eROugbE7AcqYnk+u/O
zP4+W8aSQAxyGrhn6xlKjYya3IqhV2diL1yy2KFjd9sm1/MN/B3/qw2rVNLakemp
NZksy1oUVXlxMrIeDvzBvG0MIcCFNm1axtNAINno2G/0fztnAx+IINvneoUAEymc
KK9ZJ5pAryXSgqxAx+DmI0CdwKIqDZPtPL61SWwm190bZV+69MI6bi9ZGQemdM+M
zi6TtqPedeyKwDb3//7b3N+1PkjUgljlclsntXKUkuboVadC9Xx6nYjV7r+M3sZL
rEqA3/1qAui48tsnZAKKqwS+iVENQCy3d2J5iX9WkmmhAb/8ZTl9QHiK/zPb4A/z
Dxl4I/5FxxgO2Sk7EUOGH91N1b42LCNkNAfvEX7WJk9H9CkrlE8ZXp3k4EVu+swN
fC1ePFuSxg7adh6R8O3C+c62XmiNg9T0kxkBhoz0uQXyr2vL2CprNWsD0pJdBzqO
X7eS9iyW0nWNyn/24oHpAV7tfYupcOf68s5K756bpCd1TlIjnTJcf8lXdEu4eci0
ImovRBpQytv/gxwcmbd55subuwlU3Wa+BZUluZhbrOLF1Eb0PT+fkTc03FOKaIfr
SitX3P6S/3oZOOSz10CCNjbHLEqaXy62PfjyomchWSLJkovlJMwmfONiEaS3jACj
T3QR6dhFb4tMGK2F6nUSx5HQBXpA5qqQU8gxybPoaESOG90r08C2Ipsi+j4jncio
2qPY2cYA2MucRWvyNjd+gQiRR/B/yq9+V+jfpUrvu3z8F/idRYUeBt7Fif6lJ6cK
CwWUZpvLHEAt/JkPGtpMF1sE0JJsRR4u57i5g2RCK3Z3BKsHy3VfSEehs4dVRt23
Uq2ln8stYxtDyZ8hc5sY51L1gUt/d1hpPJbrrdk9e8G1RXmuvvLGPYUEpFYzbun0
oNqAH8GCd8qXVVG8Cv1Brc6z9j/3Y/qA/lh8m4YBMc+/zjX1U0nJ/Wl72oAWg3N2
Kq8wzmexuxU1AWO0q3NgyDboHw++uJLUV/R9cPYxrJrOSNn6ojjXnsJ+uk4B27JQ
8HplfXR89x1kJE1UAKK46/SnFHr7SPxSGkweyZKfgRryzEcFq19CBeban33WuixF
gEM6/eEr1XpI+jnCXd7Drblqo5EtkhBAIcA3em3pirD4hq9VFjXwHKDGUIGiWNXS
D/p/OCgWwfo/pI5j+FaficmlErdpqUfs0YZQdSZD4JS4ULeziRiF9L1emqCli0bH
suOEcjnSJYjsSuRfl9m/0SbRWmAj916q/pAy02M4IJ4+TT7lsRl4hLV024Angnrt
XOzEOsgGpbhEqDIyiCqLfz+EifIp2zLmIzuob/zA/5Y2eGcnL8ZaRbkv4mxPtrnK
ACBEeBAhUI14r/JfsgYXsAcm3uZjRhFL6eXcbsHa9vEjlT9EReGsRhXJ5iSR3tNY
rIg7Ao5qdswwBA/VuYrlB7suD8aYH1MmiPhdRLYxYdbeLIgwgbVjoe2sxQJMgC5B
mlj/3M/MaY2J2+RRmE5mUwPEO4rRzbVspNcorG31zlbRurE+DJcdzkhbyPtCnm/I
YOzEMZZHBWA4yyztTirwPQw7Q1xPcVQZR0Umw26140+KLwODB9q070UTPOX19WE7
mExsIer4pbKBnnrl82Gya2/HD7AUCWd1xwWicNQQbSITtr37l55ko3p+FcMh9vkv
RvVeMASiXni9SZ3Kgi7x5Io413TcI+E2DXIwF9eA+oZsgAEHsIJPP38duWyDQB9w
wCm/r0GjWbTd+LepN1JrJDLIaIawERneDJchV42pzRmk1gQmzTWkex8ljJm3JRB8
mkmCqS+hlNn/8vxvPYrPBra/Xw3JVoyLr37hVmazlp6sNNxmfFlxtOeznoWYQF+b
wHTQlhRLaqPxK/tga+EqieW49QsIoiklFjH1CzdzlJ2uL8egjp4SLsbSRo182QRD
7tBZ9JKjFJp1Abl2mKBK2whWlLdq6xOk6eqyM44LiXMW1Hm+2MU25zQCbp1BDvNA
eXYNCnLMonPh+vQvilSuWVqehe0dD8nAFPqJ36443idq/1KU/PRqSpMxe4JQn8/J
NtdhgBCKIIgSjgBGKHQeWt5PJeDInH9PgxGIOI4zP7rnqa2P55BCcMXbspLtHTgL
iRinpjYAAJCMmBVTZ4fk5xP3QWRZ6gVec7gKXUhH5Dm2cxz6CpdACRLx+nV2QZ/0
D/bq6xK/vneTrRqyVwan+V7x/LZuQN5dOF03MfB0jPe7IJrckVS1R84KeCtIMana
/Q4hr/ROmckYc8MsdUdDF1FKx6SLRxghqvN8dmaq4Pn+cDhOkPT0Lpc2ZM6wWdFn
PtKnRcu7PWvzdDyHQKGCWBZ0ovGawWzrM53dW4cnK8zbhPvvneifE3pb9ozfvpts
ebcBUPmJ/Cgv4/XAYW5u02OGKSvKh6rXv24GihHGukH0NpTbr72DGsICWeuPbITD
bmGOEHFbEhypNpIFtJ7D091kOjjOOaJoFZQkJiz4BtahrlNGV3uj/J5VCHnCBFpC
JkkkJgvT0nk5rUMaYTUbK+cktsgT3+QMhDzzJCZdr/lXA5Uk6Xje/osfhyFyirMo
4Mjfl34u0stJiptIIEjn6QMyN6Rc+HOhXNvBpynXghYj5lfoYV4PZb01uOK27kMN
q5BeQztYpj0nMIe6zHHWY0zjkMRcwfUEqrM/TKN+N+6AybKt2PZlEMDXUC4JymFO
F2Bo1DUGDLfnMYCylPMEQdBZ7EyGFyqfH3cCh9WcZLroc+mNVApBv/9DAIAD4rTo
I/7CN5V8eHrnXQl9xycagZQ7psCMIwfnBf4QqB8+jmwjpu4IOFsn9+6+LHe65SDJ
2yimfT19EluOq4D35L060pz2z99jfnUUSPNSrSaKmRn8ybcGIKKmgDVPT5i+RXuI
mtCPyoKyhftoAnPaebc9jjKPcTAGhEtkqaA22nsIh3acnq+1ejMZAAuM6EWOiiVP
itUQGU36X+Iqcy7SI4OF8LmRK5ONmguLL079tkEiVEI4d2PsESZMNGs38tEWYivs
3OQphdJvxh1nz8FeZoeyf4Dcqy+Pvc6erPVEk/xpxCtvCyBgrah060uE6/KBMqag
6pr0HUcgak/o+HLwQtHNYEBI+zHnvikHzD9K0a7Tfo/RU9JZ9e5SfbwpuESeN7RL
tHgpeFW0sdyIZqO3v6+eZob3tY6+WoNP3zVoBAPcv8VIgnHnOWKxmHIdUAit6FqF
QLg0S1jqKTszZVb/vFO53nZoBUmFPL5euprksHBgSTWYCMEKv3UAI6DbwI8GzDiF
D74TSE+kB7U1g/tifPEcvlRocsYodldbDGJWJyF4vEf7UYrfPrHaEHJTmSjqKm30
2neB04lFiFzhnlSY+cHlBq/18Jx/jL0hHpsiLD/B5v5bdWXnz+N31NXYNDcMoxIg
WFnAgEDLW/SvjOOzHMRW03nSQXeHzjZ6Zppf7tOR1gxJY4QKPVOez9ca5pbi5BvF
yLZkBZ2GnI0DJYDH60+A+ltMqrokOlFUhRSOl8N/Hjm0WgdjPqHgO52qZ6nOnSHf
19CQhzwJZhWcMSOnMG4YLrNAZoOomJIXteMvuF/n60bRJMaxJYen+4VnXOm4QBAw
1Ri2zxU48tS6jhtdBF+K2rU1Ayu3Ujtzp/veXA7jx5EJfu4P3qNFWb2Yk/zuzWtl
BvjYmT0HFjyty2pF52iuQjRFaceCEOXthGrl33oGCIXc4to2KMbMhYchRN+Vxb4w
HnrWx+Cq3S4MvqMmJ63KJo8fYifnOCoaxpjE3JGk0A/k4XN/RZDISNM4dwxm0k5F
t4vf8xTssYo2PMm1VPGiZeTyUsWXiu4IhX9HmEVgWTyoMH4LutZqY4qKizfaREBF
Opz5yfTfjQ93i21Vsa+8MfQNs+e53tqk7pw3aRpoRF1Tqi9TQIlTx1ALd9AyYFWa
YkX+OuABUT6TrYQw539DpaXewwAZ1NtQMkri+u+ss2Nwu+y9az+B0RqvmLXWtno5
YJ79506Zo2eQbZswF8KSOXJQOWoxEl/7X4IpdQhy1gXdYJDgsgbLXSvTxVu+yKiS
61mHRFPjOijElOdadHGs5JbqZFbwwmspbhcauC73dXorIQffkEvgkeB/+H7guptD
o3lR74e1Sq2iKAW1o83FD04XEWNMT8rPDWV2zQ3Yrtm3lWX+Svrz+lxlXGBBEd27
a9W24wtKdt+7rM7Kv/6E/87R+USpoG+F+YPl1Cw4SKJ6euBusBh//uYZ4TLGIfE8
Z1SNa/tFSAmR9/cs/vmVTXOp9qQudZRXOO3Zxyd/xtUC2C1PZJo8cfs+wMtLpmEN
iP1tcAsXHqd3ZW67+IYpLTDsNcDlcyFwHyL3o3V1QIpUwxOEzZpipJZdrDbt8Pkr
CP6irYrZ35nlGC6GnAuSLnL7JOylBoz/eWXb/kLj8xgdI3nir6yGSWpe2ym4bZkU
Ec4qTPK1m2DA8aitZhuJezNfN6yxwUb52NUJ4B+kEO2SfhR2u2C1gVeOWxFg+LiO
LffJlOUD4GY+Pez+IhtUMLshV2MdphNVbu1EI4+zX86roZrmk6gh3cfgK5Kw3jqG
/QsZDXrsH0NekD+fJc2r5wZUzvip0eEhXe2F1pythmX8YdQHuvZV3ckOxL+p+Wpv
g159UHTiaVJmoHVUXh3NAqGauZCoRo7SY3+o9Tc5otU2WQTTI4annZ9aWOoIs0Z6
zLISFZnR5an1UiKODk/7p1o8tILOgnBSB/tpIQZZ2R/+uxqhMvU+3jNoSF2GP8xO
opggO3ffr2z0V8R78BUbUhM7ZChr1Zi+N11DpSqAmxKB2SGkd7whvDEhgGklumCp
cHTtZTvBciy35laFf9l5iJK9ai6dAPbidxa88rie1yh9PPZhn6XT98v1nrLlxrSF
FY2DYLPNwHtjM6iNm33nmWe/PMPGBWUOgnilAJhrBuWe9z6JHGR007m2LIJLgj/F
gf2GpdwD/Xm3J72BMrMtNd2oDn7ChNWnk2JtvND8pN+BIUSiryh7ls1x5hCZ+9Cc
30UfZ2orzPVM8nSa1CTxrTpMD5pSs2VqujAzpkZ1ru5SZmEvPqAPyK78ccQCy8HQ
LZW0jqFDSFbuc/Ysk44KhHH6LTVEf4yc1in3brXJU0nTgTgMG3aDqexplP6Hheaa
8L+5mtvXJ+kd148SY0HNacf+17xB87AFrXKJ3dx9kDHYzJro72VlvluNuxORvIQi
GIteXaGSQz0oTyTDftooo825KOEt73dcXIuQDIavMF1xJaDb1siYJdpPKLraUxsP
VwzM8zsyoyHt7hZf+SdLgXsFKaOSdESSYh5ASeMxO8fPcO3DXeaDfWaKSJ7dsR8R
UMvOPgxX2FRGE/cqzL+oteZ4UYw6SjOj3XEp9YhHY01dB3yIiqLqzH4bOoitHoBZ
es9/SXixD5ZAFN6eQu07vBQ5DgDAQR5J3MpjnaAy821PbPom532Wk6wTBuW4ADC0
iHrhGjY7J/QqT8ewK3LDhAuIpc5c57k1uI8ngJ3ywrB1cJ+e8dXZkzfvxWMHksgQ
1e7q+9/kmmkUFStk3n3nWrlqvj0KM644u/W3mqO0hxwzht4lZFPqSweuhvSA55vX
R6qTWjaFSuc2kuZQ7nhoXYAOG8Aae2ckGsQUu8oZz1Sxl6P/9QT65Vnn2woay4YX
Cx5RdocwkQSjZZPJ0P52N8b7CLYsAzyn+ritVNfmsmDuIvLlkZLiU5vyZLNRtvgv
fSroIhUmbIoo64W9An/Dg/qKtgHHYSayzyKd1DlAfxadPwSkrAboxTu42e6jsiSv
gCCUEmXR1vmypSltqPGhNfVRS+c2ns6HyxLHXVU08/LVNOjJy9zJnNuwsiPxs+9D
zA/pDH+MQWisdNRI2ClqaXIm6FIfsx/QGe8W+AL7SCWKGrcjy/7aZTw0oKDZLh2Q
uB3CjQGz3LjsBvFXHhRRKRnCXB1LBVR3H5IVRcb63PDTC6Qe1b9V5SNYp25b/LsY
SwOWIbDn1284+kc/frfMuO/WYohK6PxbsM/cKRP62NvzCxjjBAJ//umMDOLwxumH
wvMOnBNiMryAmB/zGyWPFW++kaRLjJ4RXoaEmpJQViUauN86O18REyGdryMMdCHK
7jIlMzFc+Q4HcpD5//Owx1HIkRJNyaH+LeTyhnxiM0ZGBjTDAHACE3Sc5XmTrPwZ
FNeinCVv+95gYiQF4MHyMaBLZYaFRlGRaBhgYXQsltAPYkOWccv9eM2bnDf/WDSb
bt6qHFUrHdmpjMjCs+CxSV2NEqw9TaM5DsNGzRbp+vAP7bDISrsZYW3R3vErTDrE
VnVBjuQDlrurDnTpgCwC4yBIc0Y6RkXgaJKunxHC/H7rqppIRuRJw2sbN+S1Ult5
gFGqdMb5HLfYB3H4Y/dujJNg9D5kpmJfmcLSkASn+OI0MXyg9ksc7cUczlRB+85D
xCnMsBQpOirTh+UaHKPD0YwfH7bI6Lz/keDtRXMm5zFrTacUKq1a1h6aTAw3oo6a
gwxmKb9a0eD5GNH3rqi4Yh2srUHgB93F76Sfl3XplipLsKzGHaJeSU4OS2ciNi8B
Yn9GgH7olpiJqiVaxu+sJFc2tzokynflpq3SEgiTFedgzLuL3H8ZoD1k5/kkAVfy
ZZRcKCwtXHff6sozd+mwv+1tXF979cXQU8e25+c9yyEWovpKhXObo5wJc8rQTF0y
kb3XJfRuXzNz5fcFyNzBD4oLCn0cf/ZY2gYXfiCm0ZJByGkHWaUppbr0JHC3A52P
AD7/ATZDCaSJpYceM1Rcz8UK12bcobTKpDl+KrNS0mp6sNQma77vJn6wJwCNfRls
Ci2V5mOskbTrtTFbz0PStjWUvmSh8Q7YM/39U3O188L2TYlXrJ4NM9df4IKUd9NN
e6ORFLbbZPFqfQZDkPW9/i8U7zglcnF7i9DGKlTADlr2sG4qf1yXaQKIWupXYuPs
6WzIcmlxecgV6LjKvCf8AxTho86Uz/BE52KYH31+yX4PpCIR25gGXRzIlJw25eza
lNH856GYbaPbe40Ybc2MNllPsOoV5mpQdoPJfBwOywQElOBhyDfEwx9vx/UghS4g
IBvVF/Cxlqy5g9gTj6pswIdjJ062x0JJgq3Sgs0RSbGhRzWIgqFBG+DfYodnCIpq
BNa6b6y6EqNLcW9bvSFPvTCZABswVpfOu+u6Xtq2bI22lDP4ioyWzBSl00R6Cbb2
AAIQ9YXZZv9LnDUfvMqcYNraHU8h6Gw+3FD9TBMvAKb2Tfqw3gZ7L2qKRCa2bD28
bL4+05Cc8NZyV5Q1cC4JqG6jTq4wCDpfM0qjz5sJZSbMr7cBjzSYKXV+zuSFjhY2
ajGq+KBsdH2BmzE008cJEN6UzSWGAMUTz9kJt8v80e6WSD2+DnB8N8bKtZRgXykg
8b/dO6cQfWK+1zJz6LjuWuj6+wcAzUdwIMtfPgpkJ7cZ7sLhBipAu6DLBDBn+Fmc
1ZqlCBObGWhjyD1P8NSbW8eYQ33WnPWXhPCJXerMrmr3wv1wTd7+z6YX6jKfqXbo
5cCwOpm3mT+lOqT7J7cOVG4iAE7We3LJZI54VjejMjPF2u2LaVAJi/6/LADk9HDR
t+Ar7AkaYiGXDLBEfwPMv5EGyq8ziGe9MgJt+0nFc9XHdQoF6Yare1WGBjaZ+dst
gdb4nAdDyrEGeNcbnnaONgEb20LuNjucfHkdA+uQfH7iw02VQh8A4+ToimMY8hjT
0ikeS4UaL7JCTpbVwF8z7qgNIqKttOeFGsfSf4nhabFsOZ0KsrD06B+7F0q/Fifp
QwTZkFLhat1ggzzSfMWjOv6/XXiOkq/jgurH3sE1POGCY5yXnrpwg1S/F1z/BRlt
2pWh+bOUNaDiIhPi/HBbRcGKlhijqF/6cqb/R45zT56mDuiUDp2gfDHq3FPTpJnX
cytTAkwLOG5YgwfNR6baFaSCrjiVsY4oxQItAn+fm59Ce4uzyhcVxZ+cnuR9HLo+
33e+4N7iD1MQ4xNm3G9R6+dI6aceuOPygOg+WU6/s8Ff8eHBX8VRxwkqfRfTsTb2
ExbJqChyB+90HJ0ekvo/7JgtCIKGDJrjtbtp3ygpiw0VHGkV10IlLeIfoVplIDqA
nz+hRITHG/GOrYmqVS7e2Hen/vRAbaeEyqUcjeJeKv+glVCg/thyu2bpotKQXsIZ
GYah6V4IuQ+Jq7SV+XS8CsXfWFTKsetQbO2zDLdPFuegmAIDp/j4haAUPeyjLxui
4y5Vzu253ySTJzwberrQTF8DOg3N9Osus8sMSm9akppoyI4u65zTuGHjP7daf9Jf
TLY1MQ8bewax5B0fGpFsObu8pPYZrlLqhS71ceA4TSXnq3ZfUf19rSBC9FxilGP9
ZyzIEKbU0oZHrBLL/dA/gMgZLa8zKgmiJZmd0+K3kLwfIHaDcT9QXaOCXTL4WCdI
JzD9FhOy5+7NczU7jRbw+HTCc3AaxfJ0FfqMHsJn3vi1OWXuzlDZEisaefqXsyK9
Ds4Wll3o0OWBrXZG/knaaLWfl0TCxLZucwJMAjr2zoM72YcRw0jYEJ7Fkmy1wuZR
vAov5fmqOcgKREsQ42IY2xFDwe4JVBRQYL9wkFdMyYROa7d/AuHbftuL9DaUjwBb
oDzDZrnHcQCiazCpoFmDXvLeCvau+rf2kOjn/+t7+0/jcHhnecd1dkICUUdd7TEi
AVODZltXH/LNt37kixtUXXwmrum6S9kYyuI1kLhVEw9TrGPddGEQPn5P/tYvymlW
NoqZSrMazH4to2OfVVd9eQ6CVprbVkE3LbI34iI45XXxQXm7KwR7U6Mdf4HfxeMj
0cnQGyg7f4T+fSzgEJE132cf/VGsc6pdk2Hz5CxDs6xrOAjTh/n+pk7xmp1FkIZx
ayT+zuGQrkGkmWgrdpn8PvrdtSVuLQDvEtodfgyTem1HWXMVGEUzLv34FU3puvNv
UiNY68FjnwhjKEMgpaUwHwUnWB0gq3c3SVN5/aqGJ3iOInPwusB9mBIORLzBgDOt
1p5Zx3JNwXwoszWa61xcUZDfgzjOosyA4vSxnxCpv+S+wfpGCbE5UC/QxKWkKSJz
ck6FLqXKDroocUmiVcHdxFgHuXXy5+nPxJ+KOYvAEOEzphZg6aLzz/A1VnK7xai6
rHfT23snTuGhGk71UXjKt8eSL6AcvpPI3olJJIUJwXmzkIWGIFuCQL4qdEdguWN4
I3zVFKAZ3S/d81RTPKKFog905PRNHYIedAt8PMgqTwplRsLthpeNwZffuRrjulPO
KalvlcDbvc6n5Ab7PO1ojK7zG9g9HIRnRFvAQXrbkicapoPtte8QKjdfrKH0eO4B
ceNQ1SPiCCHMvbnSpQD+Dm01UCde06ZVD6QA1gCGWkDxPa+LjwoIfkWqg9IsuAhu
rI1TwPLq+TsZKsUXVWbkq4ouafZgnwGBEpyNlxva57bOAQFCJXs4hnyA4IKcq3t/
7sJ1wCjaa3/CXFspnzrvja8mdNlbdnTBGlYKwaZdrFnijroqmVgmWIZj4tZo31Lx
uKm5nBARtbfRzZcMd3RJlV3LbDThkz9OIAxLa01sERU9NIP8dRd0sqfLcr/Lkv4m
x68YlaowYpJlCtX4bKfH/FG82DYez7PAkGfk4psU7lhzgSaaEKswoC+rDea2lnsk
rZnV3VSLbAlShhMIx18q5enGBc7QuuiaaJocU14ACKs/ekpdpi9sxeUQwbMjTuYv
z9iWhGjqvcTErmjy7JlykSoY6M2vAicBSapPbJHG4cKL/FgI7e8507zuPXs6lxoD
bbWAI1grFBfMqvO/96ir1jkv1iQg932FRxXGTFO86Ktujr37JHnEuP6nFSmlZ3J3
BcY6lWWj87ClC1fcuHFuOEY3K7ShAo9Kaii7d/bTZEBM8vobUlSDa5uV4nr2Nsmn
gxch52OWun0i9IiE/DlUpLAhfaC14rvcg7NOQtEme8bwHTncFuptSJE3REgCx6G2
Rc28E1wzRzLW8U0OaQ80d+AzcIZehhtBa4dcP7+Vhsfv81ZzpXnWMxL1VZtd0mgs
eAAqxn0dOxY/Tn80crTWqlkb50qDOk78dPhs0qR0NbjGac+Ki2CS07/IzpCA8+9B
W3YLc47Jldau3o0h2StncTJzEvxKSVC9+IvYx6dlASyW45Om1LjE0YSkUilNXgjY
PutSxp6pKyW/OKfxgjv/WGY4X79aEQMlcBskGIqzNLIyTSU5k8X08+nDtLBklm5S
pa2Pvcfre8OjgLZPOzOwC+XntIimWwqOt9EQ2m2iQt0KWdUlgG9QnLUFVaWcozCf
Xj6Zye26k4BEOOM1X2b8LtXs607CS499de+AkCJAej8BtFtmgZLYeHZftneChpQq
/3f5QfT443+pnRf7yCUqfmrtGCki+JcimbgOZgA9G3puIJxDsgRrVT5wVT7aUods
3ief/olNS6FPlD4BXDSmZuot2JHrcEN/YKYPVEGsYDyZnvhD1hjbS7IpFCPpsLhp
Fu45RDb0XOLLFacas63+wXC5KOZ4zYfLJ6LB2aOeJOT+FJYjkc58BLEPlGQLph6M
mnzRKzHokp02S5APr94TgFC/pRSBE9yBDMcNBohX6VtNzWQF9NHMeKl2CZGXRA7A
HUnBhfuiQdrA2wpMeZy8vWIzKJL4bxq0aupHsUiCCgrROAjjzHMptx1N/RE9Zak9
NmYQidDmsbxYJ0fu4thJ3ZFXjG1uEIa1j1UPZazE6YLu/Ub4IROOBhZbneYegtgw
cN8td5r+AldS60UPGi10HAnGwRsf7HgwQ1CwQm4EIxNysuVbONpYNF7NIy9bKKjE
Cr98cbXmvQSUQMaKakuLkYbGgF5xa2zs0P0ABn1bW93BkB1wmjcexs8akuIChxF0
GWYsSAGneM55xb4ZogX1QkUYLyJQRiGWtPvcRDwBBg2BgwLxYU3OXD2OKR129qzW
CIac/hgJf3XPKAr6LZFZrS5JBq5DrOoHg4PwoFutZo3I0mzXGnqWJP7Wuc8qGnyI
oKXOC48WchWBn9auDlfSWsaz4+VVDQYT8bG6XjAj73U9qBaAKHxL2ZijldXreYy4
XdvhgNn9PY3gcGBfrwyj7TOgJtuZRZIUvU/+LlctHfwUTQG8F5jCMtouAo8TUBE9
8pd9SllCsiDE95gOJqsn42ddYnx+k9NXRGkkRMeNoEw5ON98xYYL6/IxGjYAVrBQ
gA0gtA3ORpILLfLfhCEhkg+i/xbHguadUIZ1CL9DMTCm81i4/zbfed3Xq3f+89PG
qFEhL6rx82lnkF73L5zvyoa8BBTFt7M8IZGbxekWDP7OIdJ9nd632UKFoicg95PI
sXrRV6B68rdg/SOIFgBjyyl2ddms5JzlEO/o4tS6Q2sQx4hvFKNkB0Nzbz6dqMGY
RwptcuhyUJNWBo8CZxXGf0uY0DaejYhd2rqmV2P7RYIcm9RgCdfOx/ZE5kp12vsT
0kRDZL9edTrpkKwzYn8pSJ4u8wPfwEZGYowCUzsLXdXEKX3r37hHm0MqZ55gTXXu
0ehh55ooJOB7F+BaJ99h6fHv8RlseWlICBdkxZ/Fx+b4fjvE7c40MnA7yUuT/Vby
wyT1Uk1vBKD5/UciOSROgzB482Tksb42qSMJQLbCLorySDbdcf/002GzihTMgQN6
+3TLOWx8gJ/JvOQ1UaOvfSJlmAU4j6Y8ClEi8pNVJI9gdZ4rAV9Q3lxqyiUjTyXh
Oi03AiVaR0c332iKcERWSnG5epOhWv9z6iD+HDYgFQOVzPwqsQH+qhowZUkpTPRT
s6RkRvnbdil3WovulnjrXM5ZpWmWhKZCGMj3TNC8I5ijpZp+yAgcbSjPm07FRkKz
9sJ3N7S1seUh5wtCR17wWSpQ35KrcXk/TpzEcR58U16qkj5NKcIDY5C6zKNlpGRY
/f1TxI/niBzo7vasdJ/0Bx/CDA5PXIM2xAuRBYOyp+EqF8kxG0MjOh8r+8IBOT8p
r/AzWz8rxg9VWBXyG4tAPhqNatLf+ZK/MPclBJGPKiglyO0yvp04RUo+hP0icD90
Ib36Wi4vFgb1EQo3LOoeL+3mN2nsR28/Jvkdz1lDZg0c83XldNFlZ6ts5gW4nfvR
Nli7mqBG1GUXRRAp/Z5XF3LZ13ngl0jhpyKlMMejNhqK5/17aWNV9MCbTEoIQeyI
BVAC8q/JhWq3NUG9/3I4tqzWAJgnuJc5ZWyJANnem3Kn297kFTKk95e0wPdLblnh
Jz3kI9rWvY8OpiSwbrtdbOvsHlg+5Me0SOsWabox+ftiS6XBMBjIMKYTpHPw7jQP
75Imr3GOWBscivy/P2iHqDA3ws6KbD7BtOCem+N9qObg6tM/SYQBOcoiDnuQ2g0H
dlNghHBd3WS1j19h1crdtWjqHrcFiiSZRJaPyA7Od/9bLPi4XBJ+g9oKbSLHWUYb
LWW+YAEwg2/1TpNTZD0yqFrOy4TYSNuOQMEM//URNkthJXgDfXWiamxS3hiRNcpD
PDL66GdWv9g9BQi4QEJTXEpnbVD/EFkRm0AKlE+tgtKwaiL/JqCYMRXd9UK4hH2o
uoJqfhXNlxyi8JZghCFw1676rMTOgxUuNSZBpFvXhwAgdjTWM89wlTzPJx+9pFH6
TrKU78B+8Te8Q19tdxaVKsUapnceimabWBVbKqlt38JEOSzDiL6fRtIjXofDESvU
36X8Q9IWEFu0tLD9FrGyfU82HJjTAqMARbjxMG6lVDSDcOm7ibWEuinnawZxyGiw
K7Gf0sNuuUQcMwhLHcumZD4zDcvX6EvBGqGRj43inTS/+MmcDAVe5Wb3h27Lb+gs
hFGaURH5gfOWAoLN40oy/fVd5epgKeTwei+E4hITdYfQKe0jRLpg62TccaFyo1uy
1ml7FbdA99veKCror0kpj1iowraxnMHEMmFCRynAvxpxLCvqXpwZ2nVm7snNwq1v
OXYtT2/n38Z7+kz9aG1y3cDRahRAL7rKTudqGdrChlMmv8QsRQctayNIxjKkfwzT
Ymzx6dNlQ5wFi7J6SuRly5MzCzFBnYLbo8ffm1klwFnulNwAj/LtBBTOsl3BjeWj
WJt5WFhhsQDKL9eA8/IQIkwR3YZ5V/aOCbD/BvGsaNrB+Je704w8j41D7qx9/y68
mi6ZWvpY2epIUQTxztDPKxm2r9LcVxCj8E9NLaog16dgtG8UcBbyc4/cZDpE6mD2
/DWIArSYc/NcGp8ScE2lEqYROV8pn62G9qzIkZH+R0qahL4cj6/4FsfdcH0Y5Z68
2joeMneE3XvI4Cb7vYOaFetuNUUvjP3LwWAl7C08O+DaDHL0J3b/+vRpIOOeQiJl
FdETGZy7oowMqFSIx08mfxeC4u5BGtjjPAKmKI3dOgKHJ4KaYVI0T3dAYMlbcyb1
4MZdeyVZdmpNwfpUeaPt8KhrZR/d45upAXBzlZ9j2JAT9u0QH+3jrZocbHS7fsKq
mOJGUqEKn56NfSC/jICubc3r+uagrV/yazktaE46Oz4eLUnRJGySfKIwAgCigBmp
b3YsyRR3Uljjs2E1zswOFBRVLQbfmE716K/IDukc3pQK0tcEcER0EbWHHN07Af0T
517tqJh421RUuzNvYdXhOAFIBuVEjdW5q00PqdXhPtgB5zUOKee45j3xKeBk/GpE
kWuXp3/7zo/7cPosYB7hC6OFBo97aKZ4rRUwmkpGsDvzto2RXC5Usa0neDBevX2X
WAbMrY7hWD1UcHUEoZooSRvH+j7AGHRxOtx9ufVgSIX1ZymyHQep6sDtWg2y2kH6
36Z5Xz++KGRAWGj4iCXIPeGTjHZ8lU9+Tk489wSvk8KzH0FzxycHPjkknRJHxiOv
+YM8RslZt47Om4VPXGrTG7mNTFgFLoTfQK029Hl2BVYWSXv3CBZWpOM/3lqzy9ki
ZakatMHF6iwoSmD/K7hw+28ffTOIcbN/Isx8bGdRvM5G7idafP3dptyxgNqo7/Gh
BhUEnAQIIu3KwBASKYvMe2e8uXg6un35C7xGiDN87hpZoCcwW0gUR+AM0a4OUkZb
GLRqZa7ksKF6WPqlPxCbsD2gkX1/7gOlbwgi08lqPkljcmILImkKt1N761WS9/qS
o46hN6ujf7uHz/3rwodddu5FRSHsieNcisdUVtMpPiF17jlWRMPhdfpZinuAU9Nr
kUKX+F1+ozHAG50Hp/dJOt4VKG05pxMoPHJOga11ZX0ONa34TP5fWJ61bJ13tuP7
OVQZR7iiCj9JzcK+BVTeRuXrJUlfQ3XaOoXnfiDN2VTjLGYSTNJQIo7fOq0yxDm0
vW/Rk1xRzowji+Che0oy6NfiKeQA1GNvYlJCZtGwJYWUqzU02PVByc/P2DsFPOsx
qkylr/C8a81XDGHV/CFSgC9tyqai9NWhD/W9pLb3b/KBhq16dzTHSsacg8DMPIv7
ttti/Aku3BoNXumDuA0XUioTUOTlM+ErzBOHkLVTJ4yc7kf3q2JRqv4KXuwMrHtl
y+yuoZlQNFMBFbn2Z7Mscjq2wlNJGVH/bgNAzlHjUoC6OML/vbk15rHhHCgIrLQc
B3SI+A7fGz3ksDrV6fFJywkWVsoYNBojJ65WaF5dp2/4at+LCfoGCegacGfLEd42
NM3Sdn8RBfjqOSE//w1DaKkKohpqKFVTll+YrNLvgI5ITEulCEE8DJddyQw5mSNp
hH46JmxJPYGWQ+bvao9MvCxVLz3pubO2IBvN34616/OgIuK/1HC6w3+kMS7mXkHi
4y5xMpeZq21Oqtbt898vAFnKWVTwwpUV/0DYdEkEKC542C4EG1ATRxGe99/zk/Ul
kIhaeAQNteAtVcfTo4egDTDlJkLEJ0xdJuJE5PI/uEdT9f3HcWPkBKjsbrmN7Txs
W3BNxLzhfAbrCwR6j/ZyszKUCJ0mHo3cBLgO3483+k1pPCYjNx2TFrthTrDJDfWO
5I1iQK13vWfyGrHWPaZuNhkviIuxiK2gcJWj/O7IVcUCrhE+oWngFY0vUbGDwFqQ
XfsFGUOIpCnUGB2B97fkhsBHh9E14UHrbsyy4yf9krKAo6jX2GlsPBbZ0VFQHTuv
NfFpZyzm1Vrr2m8EcWyciI57nqXRCI7iWlS7V/ljYopYcnJrPrzXQWnM3lYjRxJB
VqSA9lkLaXzFCi5kBKUyaQDaisbxc3AN2If/ktRvpPy1c1xz4HPKi/goJulD4eiv
rNUZ/7c4Sz+1NvdcPBFrWErcU9b97WoiY8LQ1CqE3f6+/KiCOvS7w3SAoLsdxaHM
0U//wpxWccHTawYwjVeG+UJwst8YzIfvEfrcKzleMP1OKfkNhC04IXgmnlNy/qTk
NaedjlhYx7vWfJTe2jafzxmJvLMxBYKXk24Cy2gDhSmXE0i0hIpmkYH1D8/ti4Z7
5Y7GXxrdxehVlyQl0pguDKLdN76mrDMwGlYFgf5zGaI7ELrKNA3BIt9wxkjSUrlQ
t1M5kwRosazaCpQgab+Px81gTNiT0xfATJsqYRCHmWWwE/mpAaKxdEIJ6f/Ea26j
gPlT0qIOUKV9TAqgfBqksu+4sqdENHoo2VYI8IXpuCrXCnLTP9g53X0pjNZBLcyL
Q2O8rl+Hla1ripltBHQza+86KsWHwPuPtJi2FhAy/fK/2L/YYPGE4P09IUf5GrM8
GTq0eLvZqY12ACMKEOR5v5BC9zfMOQ1iu0Ab6hiohbisHrmD1IT5uQuwfW/xkFLU
Tcj6ENkwXlmHFlTmDeSH3qH1A6tDOP9c7ALvrvcG+RdzTOEQeCyY+pjA1JyH0hFx
t+OM4Z+TTO4HlKcpT8RpETxxs+P/4WhslVO0lwsU8WaA/0FUKIc2VU+vF4U9QT1o
UppqtPxN3VKa9+vzcac8NE8R9mcNF/H4UBBOSiBvXn2rtf4iY/JrE5JIRCa3EVY8
JAF4IJtn0SDrm8j+Syoi2jfSDb6ihgAPCccku6VRwDjAHnn6oRFXH3IPkBTOzi8o
vSCW8WbVCk4Xbh8/4w6Pk54CdbAncC/dKyhPs8v7B+U4guMLujeaigDDR4/JvWO3
TIFjSWITjjC8CVe9pA5/bD0e8qe4lWAMQ8GFJdKhwIuAfLgpP8/lLd7+8jCrBCJa
LAWqYlVwJ9GUPx0Y4qnyM+QxqmKiKzNHmgsZXs0BuAlkCNGv7fblW4XU+9Hz1QVm
6zXVkrRdpC5b/bBvzYXuTBMwlC0Tl2KQ4C1yyFvExQTU9rCThLwQkOcHxzt/Xwaz
Zx0HJInWEea2lQ8THffRKUWhJxucyGsO2+k5/bHlfG8Ral6rm/l6IJz53mLPrHhS
iOuhfoBHJm1GUSrgTKV7Mxzmbmq+ZScC1OGAWlfhsNoVA9xgyyR619bjTRTPto9l
Y9cBjZyxlNJTqQ7nCOzjKFlmgfMauNqg2Cxz7jlT87/lsz6SYwG3IlfEeGyZojmf
H9iJ6gNF116l7FRibsrbsSn9sbwTMFUvYitAfUzHEjt53X7uqujqFppIqVTNeQYn
a2kDrN+uk/sVvJIhDG33p1hwD+FzfMHCZvoCl0pDEAeAM1tdHNEz4sFa0hapdZWY
v27v4glvrA353xXqDlq0/rKVcn5PUhsR4HPLHpd3g+WuFoyx3T19Oq/0gzxJjaYk
yKWGxQgws45PjJWtxTqUeVljin6CYWouqAhUClZC8uMRvmmgl5TZ565sQI2JhfcP
Qg2cEjFMedzLXAUGBGLcNWTeC0HHcEisl/1GzAb0TW5+PoKNXKuJteQUERHNio+u
RqSRIvA1BDCxjAxDFmh5z7lXvj0skhpYicEPuxvSnLVq4hndGckeU3xpdlZscPWP
CvWHb52zwEPNPpOl7CjHykwLY/cUZ/TcmcPwbtsBGyCkM6EYZa+mpb6HTNc4GO4w
428Z6rN1c6OS4aK2VF4G19FOv3mVNZ3/7dPfKTictOsB3jmgDdmrELUTF/0WUOW7
Jn9PQNp9CEh/ZADyIYV7l2iU+ZAZnQn9vB3+ZylHBvbPkltfRDPYc2D3WJoHrmeQ
B7vCz8TZVnwH8ZdXaGdYQ1+bGioPHP+vLEfbBu2p3mFyti0mqHoE/hBcl9Ycuy/n
4goegomibs8++DxCwPkHUNpF+dN9fK1p1oENAaiJsfHP5666APEdWZLPQbPN0tG0
s4Zzzgn2ReyAPTtwVPsWCiVgiVju+w3HIqw+4b+hgxUkEdpCAIhWGreB6qedFQXA
e4A0YCByz+TIjTY++eqA3mM3Ft0YJmBMjlw9l49vmM7ugSh6C1SvmtDZo6bTXpxE
ctsWZ7ildbYRdQyeP585omBvibmL/59aeQR5Ps2hWJmnaid3OmIEW6NXWs8m5OO+
1cdO13XHbr5jjMAthSPEkd/H/N3nk8KmyG0f9PhiWROtrhgXOzVEzeLSyaJmHuRA
BlyOgi9pE07NURrQQlG3TcNu1p7WN1T8Jws1NfSqHoCDDv+C40WoscQ9YDg/jtyY
RbXls7YwQJ9Td41bJFSyOgQfQY2vHjqsxYsq82kg+dPbiIhKc10kOvLkRwh6eBa9
Iqp0HMd3auuaxVYLSEYAbJBL/snD6Q9TOeOpmStbAoeAk7Q75fDUn7h5Nvn++27d
zSFxqFwDJq2iQ9Kk3CIvhUb0uOmRB5U3GB0urETrieMygPTJsY3Xp18YtnuXMDOe
qqvdHoFaDPivI4aSL2cIeMXUgBLhk6IueOJRAjaFQZJTpK1t7/fgIXcYAvXUMdk5
VABWWY9ErTAs4RyQMaXnb0vDzqYDCaiHkjyaf1cp2yg0dzU/wExj9/14xvvfwsqp
069tSwy7eb36osESZQJE8jQ7QWi+x0Vt3QKrz+bp2xAVRtpWsUJecSdsj2yE616H
Er/t+CMjdSLQEN9aEYMTqKojT1pAajcL/Dr/EBFKMLwWjTUgRFU9eOH9Zfnvghm8
qeUu1VUbqs9bJo/MzMp0J0MwZ8xWNiDDKgVnN0+YuDwKAZas+5E62mkQJn7S/AbY
+r2C3/WIR0QnXXB2j1e6quEiW0uTUxOeX88OVfXtIWFAxOEw3XjmqfBW+OVgFsEZ
y7s6qnzHXVP6ZrtVzwQEr0l3WEk96KOcf4Ps6BjNEaFb1c001UI9KkBsLNm3+8YO
/PjNf/usIbeUHxycm4o6mpg+LZTS3NjcvvkQZiOnlVlXzrkVfZraHEm3MB5IMIVt
hYNv8fB6ROg8MXEjOGEsmII0masmquPqxRvI3G/dqZ4K9OuYbeVNr+ndzpPNDF9y
yPoBLqTsS8yFw+JPLPEUd89TyucY24keinu6SnLcj9fFxjOfxoR2aEjQrHsYQuba
D32q+U3hClrnmj2ziW7cbdfxo4mJDa1Re0RJzVqT4TZ39bQhQWL9ErHU4NMI199X
hW2KaG1BG1QU70dqgC6vOpnlxCyXe9tzhm3dCJsaECR1B00t6vflAyKY8m1J/Jlq
CovJPyu3fXTZwmo4A5uX8v2V8sUi//toPEjNMTJg37XIM0tfFSMehEHiWkUJazrV
cnfvTist8xqFSW6C43kjXnJ0bDDvysAGZLeQBDFNc67PaG/MP7Gg3WXvy9zctz7N
gxOBGLfZCFXI1Kvw9Me2jlv9Ub58EWxTRY3aXXgSnOKgjLTQAHsxYFXCbQjAfvEV
iZGRCbTi2MCNslnJSoROaHsSDxkm2qd0N+kF2AkclGJDvfGDMsozqM9sJF5G2Pfb
C6ioIFxrp6wE658u6Rd7w5QAfpAmMRFr7/n2MrYIHFxBhEymeIyItXWUvGVhDQCh
XcVfAvIjNnPoeP+7v1jpZ4rUBABtN+Eb9IUgGf8DvRB+Zdk3l2UnPxEbz0ZugVMT
jzpcm3bY1UhTSL8pg3kPaUGPsYBr/QT38BAeV8eY3AxebAjF4bnbJUtlnE6/hYUf
MNdkDKsBBjXuMD/Q+74IGVyULlv+0Sfzni6C4WlZcA/KeuC9aQvRts4T+rXC86YB
rLFPirlq7Rb9H4r+R9mtw5xlh16wXwYVI/FoVd7sBQMF2gNIwtCWpX4EA6GUTAFb
byIBNtFUcl/EcaKuw3Xf0FfqWk+AO0x4NNy13o1uSU63BtGeNPfPdSsp3D9Dmstm
h9HPhvS01lBcHD97gViVtIJba4OVSJYynhwAVv+w80dpKxUV6oCDauc+InqJbU1D
FL4Lb4f8QtzbpUnSwRsjn5KYtzIF/WyCZQETzvwenZWjviQ9oykue3GElydc05iR
qFr3kY1Scxn8gTi3HbPy+jJcVqzsJUOVbzrXghrsKrVzy9jtL7IKRUuZAnNSawCN
U9L5hCptxzfB5fNG2kd190dkJEpulRLyfkpO1N+J85eY2HFeB/WxdfEwaHFnXXrg
C0ZDylSI/zKVZbPBTfcqSxNMQgOKpOCo86JM8vqtnuxbho4M16EVuJQeDfOR1b0N
2KiCpTobkUXcmCKVslX+Va865LDAejuADDehfAFqP30B4n4y4nbFyrDUxKz8Mo3I
me8qSZ7/A8CCWH11r27LwIUH/icEVrOGmkbEZK0EnSJ3rtwfB5IuedAwy6hqhWzX
KUigjKJiEBUaTuDk5pJfcEVDqyy0AcR1HBglgVM5G46IEvcVj+Vy9Ox+XaYSB/KZ
BDi8D8EYhzeYdk1APuPievduDDC+yDdJGYdc5J0APCpUsUn8Znfgi1kaBcTazrUX
sZhelyOHhGwmNV02dd3iSH08claXMp6umBJ2tEHMM1GWA5mF7QCTD8YKcfbnvErB
VzP4oAUUa8OsGgzjE1SO/FbnB6C72dOTqF5WIzTynaXNw7rhJaPmWsNlwhYO/uui
l+hpKR74Il3jlpHlOpi3j9yx6pzJowHijb56JFXvxrD7IgPCENnur82KJmNSSpOR
rDls3SgfbWcmCeprC29MC9ByYzvJEoM2RV7Q061cXMMdidCgqbcTEamk9tFryq+t
BKpobPhcn2puQJ9BkfVQR5eLzRqWEVs/nrqyT9x1O/9ho/UtXZKdNBjfiCxtJnSw
qVYo55BKOOzCMIGnMJ/XBxV2SNT4jRZVyr+BFGwmSWBNhHOV6MiZ/FbsQbJR+QQJ
zPV6yxjpfbEjCGvn+yfdAxdcUXm4QAXII9Jo5/ejW1qlebMtcNSyM5+VUITQQ6yD
DZpApQOWpJBVxSGo7u+DceoZxVy/8e7+1n+PJc8oWfae69tXDkjg/Ik7eseAQ4Tl
AxQDscBkgqgG5hJRCxCOFBcu/I27/LPWogZH0datKpUYVH5eY/XrKcHhyGDhjv9O
+oXBudd6B2vd+yrgh/yIQPeME0BW9wAo67s6jvAYI4iERxQReSs2YSorgP4LdybZ
SNGJg4UJUvSaW05Kc0KTmi27gIgI8FFSHZeuA9lCDCNM4YBCut89mWHpLhz69QDo
ivPUogvlUJQ7hURjmdKtbD4rkiLV4dl7W5sMc4jlrkRvDSBkF3t9qn1FYGwZR6VG
CLqH31IjEKPYcsPEPJuJ/KNTfd7aaPctyLzlJgPnTCuq2e+hWUqLpd7F4wKXZOIU
9Um08+DOE1ygUJjX6w6Dk3H4CPqStHz4p2KvGaDzq1yWdMBCAWGlKb4uoeMegqK7
WmcLJpdiAGjpCLLquPo0lPyq3S2XHT61EBJqDil12rGq06R/WPeakfhVrvoDOS71
ASUcubxohTgkzSwDxVkZc7aWgPd/nW6LcpyJXju/OF8ZK6NjzoBxAFrvOVUd9dIW
qc9FpOCRvv9SUJCewYqPnw+ggFD25M6/yFmWbQwJYzauNe2hyQnxTv8G86k+FKlm
QnG2++B2/aeZi2UEUGCUQD0kUS8gJbptzw8bFCkrYyGK2OKzEYKk3DUFkGBvSA6T
ao5lL3ZIs762J1fB8Ql4S3j13EK2vLBVCIZ04tR92gKdbm5nYMFeFRLkGFXx/eyG
wSOYAz0BWYhYhlP1FfX7t9AulX88hBgsfU7YULbQ5uI5sDd9lhbEi16zcaS1vqM9
e0csOvzQy8zNiBFe74R503x+79CUljfWUpak5woK2lpsDa2q8fs52MTZLyCAsAhH
tQcStidOVQPnT0XDUk/Wt0blRiG1j2gc/ruviE9uAOWJC4HDNTSvFEiKOKV9QCco
ZRI+bmiK9QgF5jb4ySBHp+OiUQKy6qphRjtdMfTyNxM4JdTRv4EuIs9y4lugqdAN
zyJYsMNbvlBdbMOGejcoRTPFmHSGBzWR0bpFiwk6/xpsP6Fi10m5S58KvwyM+AWP
0OA0JvewIVe5Aoaztq0O/iaLFoUCEXYjpT47UGVvZbrJImi89m/BJWnAHRv/vSxo
UpeIV+8f5H5Ga8dWv9Eo3pGf8PXN2zxx6BsgqVXuj6ZWe0pb4WlXFZeRKDe+h1Sc
Dlt1Dkgc/mZ4nSlbw11X0ntdf0JoqL70NQrBb3Sob7m3eCsZ5p5gCatluiysW46o
Erijtbb58x2Jg3jNvS6tTUh5SaZF2QdYdE8mNduoW0cSmm4jo8Nk6JvuQI+ZVSse
3oYa6EK7NbcxpsgXrye8A08h1vDnDJaP55GmY2ApVuNn7CxCtr1hnchjScQX1ASv
4z592cMC6C7ZY6GaftoVNvn2KVZNQrHnnIm27xanmt8KQrgbDpPJtwwiIvNVnBMm
tVhTaht9wjhx62+KY6cM6qVvSLCVgQjVc8HZ+KTeCcU2GI/F66/Q8GjKxD1sz7V0
NqBhZRs8ZcOud+k4OmKrf7OM+hAurUWDIcEuQ/yg6x4r9+WiV55Hvb3BA1NlGQt0
bwImgyq5I09ACYK3Lrwe2DEE/yRzg3HJjZZE7GIDRxUvBxYAJKCDlQ8yTVmRZCqY
RaS8b8rYfNcA97cQHmLQwxX6bs+m72Td79SP+hBKgHgrvh5KChfsUUuHehdnr18i
GpV1o89YY0tiUlff4KIYVfdLgBA8NU5kLjWmnL6Is24FIeuGLilFH/qJQRo/tu7V
vdC4wJUcHZuG6A+D6VvUzMLVqhDinSbHNmk2phJKK0vUhEUOQfePT8+DGLMJw7cO
PhyWYiosnmhT3I5Jq9nATjtJAehw1kzm+FblJTEX8TSqIjXpwKwdJrKROO75bN2o
zbzkELsfjndt8vqLLgTKFv0Q6ePepnuhhRWvkqmxRwugPRa7xnQGq922qRvjr9XE
QtFVK6VlNgDe7w0Qd8XW0MzC3BpSIM+q5q2QiHJ5uVhoVd5f07XPUrKHiG7MLWda
iM820zSLVRmVrHe/2ScPGNzidPZOrFcDuFqocX7QcUWzX6SefqEL7wsTM6cqMKHY
pUiNgCy+ayxwJPSW/Msd9/azzbHyR5G8nfeUyVin+JoDGjqTVSFKTpcqMNP96EVr
fGtQ6CeVoaWNL5v1Fe3qnVmsHVongQnu9a5I74pBsTQT/YebwJobg8/zlK+mcWpM
WaalbcScUQlZaa9Sv0+LinT5rzbp+Gd+3eCkZ1jkjHI0k91sppaEPs/xJ5nO9ORK
zqgUD3uluPcLEFRes1QbOtevYAoRFY3daYgtYYpqvenB/KHQSTB9vEiJI3mCl55Z
svahdN9qOYypapkNNWHwr66ygmSHsWkG/evXg5xZSclko6WQnyoX/rlgISIX7BJw
OQXjRL7KhvXe7r+BKonnmZli5OCkHv0c4S38aDqWO1TwCquxBtsNIejJCZdi3ADq
+nldUT/SwX+xDvyOWummdiFO3BRmFJzBo72memKJ2IJ9CYxY4fhTrsxwqzSHWtCV
0tcgbqC3y8s4cWfO5cCiryRfcwwpNMBEWDCnoyEZMsyB4+ggQzA8PuknMlh6mK31
2Xn22WGAriyoNZyxf968dCaWrl9WA6PXgJahJ5uwfrYLTJ1jh4DkeaQm3h3dOMEb
LLxdtxCAR9/QvhQVxhPxioBWJKWxRU6O4BmPwzC2qdOWK2cWZ3nAzG+E6p79EyeT
Gu21PALPjlvzYByzmX6mpkEa+G4mVReDBBhdQZvjt6w/uXaYO1Wtzo4bKlT9q+bi
mGUtNCItIup7wHWeLW9ws13TxUytFiG+gkpE8dlETPcR/6ovj3xA2aGJvOOl6AXB
BGNBfVJboZ5xcmKcgV49KBQTAnRseBG2UEbz2T/dpwCJpz38KUaoKgkNKH58NeTe
sTXy4H+igLomgvv3v/gEoIa+EIuH6PAUFfmtVHG0S+3CI7yivIhItn2guJxnIQ51
1Eo2a7x7Nu6tvKVimszTtbAK/++3IaZLnWS4XAmFk0Q8wBIx4tphbCPRVeiQ0pVt
Gf9ZioPfN3Ct554csgy2dxh0PbSTWw2b/lR4ow3RIwNq4C2r1f+FFrGJcPlA2ShL
Fca0NVlCo3gAGDOzVKUAJpUD24zCKGhNguWG6P2wfisMJaN3sxNdudVPNfCWG6nf
Z/rTIB+egiKCvP1J+0sTsantVGt1FNjofGpUqFBlUIO48sDcRGgOdLa6LeF4I3gl
OqCorJ/CLyBL016BNt9mT8IA4QE2xGFtxRZsVxIaoiGh47924TkwfvejiklZycMM
RNlm4Lkw/WHpwSxY6oTtFah7GSAg9ranz6Lel9hngxfTbrYieFv8gQqgy//yo3mv
ic5MF3gVjsdlEfIe49J8o8Ktmd3xa2cvtr0rEBnrn6W/fK95hAiMfFSWkqRxBh0U
i0BrR51jBKFghq29AoIrTQWaWg43o6kMEOiD0AbcA8JiIoGeat17PJ8fhQaMGfjI
uIIBZsggE99UcDaxNjHFWFtYPZV9MHd57ukFS/pOiuejGwQYr6kiiqACyZLEkfZr
44CIDnzGP72q/CpnAbI7qV+GIMSR7zMueIXv9IASe7+YJSt/tWEMjdMxFKS9C8TU
X2VeotAEEzZz5v/SQmcuivxhEnmKvFW5pF/FiTsdkdxi/Ov6VLuMggAlHXINWYhB
WI4m16UUWVAw8+jlMnsExfCz5w9InsV2U8RKNcsoNWyo0tFehAKex2ByIlr82qRB
uOg6+oC7mGNHBL5/SvlqcnLCG2r9SuHr53w0e/C71rVyOlrJwQ1AXZexwiWNjS9i
GLTYKcRzLZEWvzm6SNTqXdvh1r4T94cIi0hSAcVQ7n2I49fwsnG8a61jizpV8gHX
A1d9XYhXox9gPKIjGeUYppBz6GrdibO2FCAXXMUlN6/VI3NLFLRRsm8UEffi/vHh
XcbGs+lDab283w6wDklXcktxdDGVIAldmIra63Nfrd1luQiutLmkon/BuDT8dRsb
g2LhtkdTH/rUUqtpNXS3Ymi6bK+gv4hKNqXeCNQciBHJ3ibSdWrIVTJBS6OUuJ5i
li9S9uhrTSf5xd1ChHOse/7epq0PSq9y2PQ4LX2vHxEQcTtoZARA1+6idC4Nz+Zo
08syH/hSNhr+YfFUAT6aNLAmgt0HWmd8hVTswyB1FRkB6nUS3VfGtUW9oA5ZIMV5
qDMoDn2ToTzmyPtahvMsIRVxdFyDhNZ+w0AbZRBuuRNAleDy7QRBrszC+8ui6yzs
qKwicnjrPNzTS8qAL0FjpaYyRwATq45+g0DsPCfYWocYj/q/qgLclkD4Z45m42eZ
3TyvNtqZ3hv3C0EJ49rXG7BbamY4zU3dPi9uScy7gaOdg2diI/qRu+2Cc7wkQ4fy
y29vE+r+Z6/hzdNGeGn6W2Zl1/+UBQYKlsd+gKJTlzvw3e3ZofB7ZQOAFEa+1lgU
YU/c42Y78U8O2Wy8H6rKxh7VATEtUvlwHY/BxbHu9tRkWi43bw3sr5Bd77+GZCdT
sSBW9emEHlJASUKztmtQBSLZwmJKUjtzmGeN7FqG5fr2VSGFnhpiouSI3QgaRoD1
yprMgTwVmSy9dzQ1bPtcuyTPpQKAAI/Pz7+xbDbcXh99+sYnOc6B59YTPWgF9Zsx
x21EscP0qJNnIHzwdpyKzdS48W92tJ8Z+6XmdO27664tTvIC2MWWBZEpDuuBw5Ke
DwSGnn0RvC44YIQ3jDtx7UOCC3HEA3MBi52iNy7JKp32aWWNej1qRHD3vFE4SL0m
P291Z/BkLmpkiPULqFytQ9nN1kzF43StanocGFn+HKv8ocl6faukVSwZpey9DtO1
P56vkyhcbKbQv4lrmW5K2cie+AUxLAv5F20ftjZDTHC8O0IUOiSqcT5MPtf0urCO
RsMQoTdxjh0TERFfvGUQAFIpxWOTCtkoQkSOp1oQvMXhDAQYrw2zV8lY+ZqE99E6
7tOAtDlzSQX6ubd/aACB8rfdbj/BOQdL1CQMxgcJdK0HEmNPg3+apWyieHyfxRtO
RdpdTS6DYIa0LMyb6wYnihozImvAEDJUWlcEXpU5UISHjxMek1f+HsHiMqYr13Wl
Suqy9D8ywF4FXO6lNi4Ae3e9QYYYLBYN0+zhqvl+zVJLGRc96IrfdZV5EC86s8ij
PvGToWQZn4X3SF7DWz/BOSk3EfzQEGIPTa3kHlyTqKWlPnomM5LpWu7G8/vBm8O8
QdkRvcParbLeaRB8HFZ8jXqLfoi974BoC7xTWwRhY2s3fmo9mAbJBuqjPhh992Dp
AR2Jl+BsKo87AT6UIxKVtqWwimpYYuL5Nj0QE99i9Qj/3rbKfHXhlYt/LOWrt17q
Hg5hrHpEp4cAPApox+qFdWLaKXbKjhlAeaGUQHQXWySX769JLUV4mZotoE4AogiQ
mXLmdOzqc1HS/9arP2FMxtmt0dcV0XONrwEvhgcFwkrcgi2zFKjt4ZatgBXIMYVY
P7w6Cz7y5pgwLv3jDDDqCUksxCLWKBGBWFekyprT+cW4W/UTGtdIOPSeBYl7YZHM
k7RVVb4dNVqWl9xNh7TVWBzDfsSwjS7oXtUTAURI1V44r8Zx8ODhCHe7hgPKKjan
cZhnHTXlVUbYj7HA/NKiT7tRNyhyKRYlxpgemlFa7yAZSUdrt0RYXjhSj9Y0AQ+3
Ntc2FSB/YXm6IA5v4xxeHJPt0+3eKf4mxvxbPOGARKna5frUpKbFLlpCbuwlhRd6
ZM5Xdmh5S5HwVs/hWN8mXUPmoiNzLC/j7tzEKMcvZb6GX8bYQ5uyaZBUAHvyoB0F
+JW/04lD/Qcnnbnd+PsfbGXTX/vOQsqiQoEzbqUIyTo8YvnD+tEszxfCBC7PoNVI
ZwgQQzm3vTp/pkJRBalMpIsVddRcC495+U5FIYG6jQL88NeWn3OYir9RfYb7jpzz
LjtNv+6v0Y/vkQC51XifAMbV+jINTMCXtv4UWfB8uH3JEP8fzwPUrhdcrCD67WcH
AjjVaUMLUxFRjImnr5hEgghWHc60Q4bvb8upHGKdLxVOG0W9NC52fyH2jK1lk5gr
jc8dQ68Wvz3tF/CHXUJQsarN20eAeufDy73BlNgC4cOxAn29YQRkaGhvd4vqalPK
dA5TuKvOwapByylfhIlK8QH1DkiqOCSkuWvsK8oW9dakd/ju5Y5jaFoIY0/ezuA+
LoHqpUdeqfM/rIEp1F+qCSBxh48p7ORo28ZoOui3xNp/wwyoW3rMz2K0R/4r+sH/
oL7ssBS3C44NbnsRTkavVwVcYk2UOe23mooxbEIBsmFgHLb0xnX+Z3M2JAORB7Q1
P18InkZd/ecJyO6qmt3wBOLsHHhiRC6d+4r9oxdA05K4w9pfL+BzIbBN2USpklLt
fxGcVwh9UbE1zytdBb7rTJ7/zWNigJRilDuYWPy/oWhwjgrVGnMHuUI/QaldydKO
yO6Er2Hejj86N4gWWJu8W7K7qLboZQqDAnSjluzprAbrUFVUlPO+NMz540ZtUZYi
Be3SRuyPblr1xf9eEU82KQNn9n/9OyG8Jxe/ZQj7s7piniwVv6cn2Uq32D+Mj+Yn
6lEZt0k+AWDkaOWsciDm13l+Q51zqkqfcjQL1tE6tcXuGuTtNiYJNIdvovUNAt6V
Wwt4hqNTyguB1igkQvZuIMaQ1jb212EDMMYLzFB45VDdAqOabcjF2dwY+0tUDdBz
e87n34mnM3ffMjrPqYFUWZmjI8oSHD4qPjoyuy+5IzLdM8749yIZ4fmvCwsUh5rz
jZnafRBtCEfUo5eRuFlXfS1MTkfDxidbkB9aEpE0dTEAFUH0qSGHnJ4eHPH1kKrs
591ArgCTFOMYzLUH8l+iK4UeaXNLYKCi1/du5xuc0/oG0Ex9PiLw0LuahCA6wa2E
JkMl6aQn7pZev38Fv6MMINWeQ58JhfMxnhFsJ2rP/hbmtVI4eG4I/5JI6qFaOjc+
dL5YheVkpn+P5uYXM7PjPfx46PwNGavLG5bc6zOCZuwzXJTBDC94oMpslnKHhFL+
j9cf4eT2Z6mmdfv98LOxNatUX6EBgg2CdnhmBi/1O2cT2CEKBpwWWtZK2dZJ0xPD
p1SJDy/WTiHagOyGHCUK+YErYHygyYH1gBFLRjAhkuwnXvRF5pmxaVvOlFaDy6fi
dWsXdT2IOJ2d3ns/LFXbhSi9y+/bO2o8io8YmLiL+4t/CBn9a5Fgpte9SIZ2Dad8
dBQpge3HNCrzcNQuArFCV05IGHi4ogEAWnP72kHxxj9y3gevH+qeJ04JSnbQ4Spz
vX/C4Hlq7iBOWtAkZKuYn00+iaHaSi60G34nBQBhwq4Hsi13F7QcHsmw5ldZ+j0L
vaaKjI0/H6E9CqgSQNqST1hYDrRhWlwQFikuAvgEXASl10HFIoi4NGVdWXB+5GTO
VUJd6uzDEzQd/bahl1v7uWfzu68Lae1/Ap/TGITMMs5pIjifQk4ZoXg60Lsg1ff2
2mWHqJUKgTwsjWhh4TBSBUb3lExoFIFbfIXTCNNYU+CYBMjJeGmwAYp3OZlGZAix
sN8BB0gjnjAE7EDxi6vMZirpIWA+WsEh79vbrv42dK3dw8/225uYaP/u69qm4E66
NcYD3igBwpR3b78ozyrpzZGPkXH5U+rG1rS8U3YfO5BGr7KcEbj8TaqBbFxob149
yuoMw8b4oLBsgTSEED142iM0SXdCH5jL6WAWGnXnNY2jwc0dhT5Kj/nIClBEsQwU
zZ1Sla+Iqx2zTmfMBlae5N5daWz8ZilqHszwOBBBICDaTp0v3J38H9gFYgaar+TZ
Sv/NJq91jWPngKbRLnw77gJzDKegVbEO8feKyW0zDhhsF0RXb09X7kUCpFEsrtlT
pVx6COnks65hnmIc/WklLmbyM6kp6TTrAGshMjfBg/lj+4sft4rPafe6HeyuQLu+
rLAiuIuqrpiFchc86L8ti25O28c3Mzg0G+IOernxxwk0FoIAEufsL39zc33saoup
RN8/YON7iHVjXgmooUTh/mSf28Aza9h+zUB97ZaogtugtBG+c5jWvgL6kQp8fVVv
pBNzsOiM77tkWZ9L7/6YUALnIUZTvaGros68DRRPRY87gTFANSb5NBr6LrNo0DQ9
OWgLWLWc7sNz9OHHKayOWHtygFYSw2CbqTG75wjT0EwAg33oOWsgL0M0RVBdUTtk
Vb/4XtK/929HOjpiTnRVdpqcASYXp4lujEQCORtfI2qaM2lFZn250RZ7WP999K1q
BWwTrytiVMKAm0+hm4trjR1VIxkqLMeyrWBzXdx5AHTTgo8VL3HGMcHhusbGNk0J
tpAEksD1K8Aaurx7NUCI0IaQsmBdIV95bvnBhUtB938qADzVDKvFpDYeKCYEaV9C
tYOqRuQAHB+xdm5WfKEMOiSX/nbaRldO0rUGmx2+373HCS8oP6jZxIKbnGHpOok6
1d0JRX+r7jm7+YkGyVoK4Lf+/JqG7KurcYqhkHf+SKES3vZr/Q1KIEV811X9VZj6
XqTkERbzWpQtPJiVXG4AKofdl0m5fl9c5wA5VtPi+/xN1vfICZXpXmRzjByDgYwf
4TgwaCzQEVdfoALODQcu53Nb+4g6dx01jZZ7rEJsHZVjyelp0dS49nBx/eoUqTtk
fjzvVpsB0cT9dnUCK5JnHUuZbX+1bp2a9ENKPxIiiCAwehATd8Z6RTLU7kfK4p/5
Xk3D/sIfUao7jdS5Li0Kqy4xm/XtLyaF2LlGtW7tZ0zX0SxaOzy0mHa6v22+VmBl
Xob4GgKi7uJZ51xKxdkQTXeW1/HNEhenFLI0X9fGfEax5xt/LU0h7CFNeRiucTlD
NP6T6FL+7UKVCjppAY6TM8EybpTLvpL60YxkC2LIIc3oCLFzLmyBcG7kxk3ysSRu
LQoW3uTfSTs62RsxiwrE6UOvw/bWQzjBVrSNb4+8Go195rnh8vzqruyEHWFLI1Ib
hW9kmUdhOrR/LzKQvemnjlS2BZy/CTbNSyJBZLIXUiq1XodJ1j+wiCL+8jtgSkcU
ulWxOKRwVoGENpCX2KEyIAIU8o40gqz65pVwGGfFt+oVsW98psnZLyvA9LADMlhY
JB7yHZrdX5mjkqQ93d1nma67w2E+tqNg22K3ZRf3wiUfw1d7G8l8jAeJhBCDqosH
uezwll7WDfeZE0mWlXZAE0AChibhafV8oLmsHDY5T+BTlI1hN6A8GkZaR5nXSHVC
CPOYC4RpKH6fWRpfHkRwd6BBwMgyT4YUM75m2jE+P14pLEYULW+eZykysqC2YxhL
id8f+10qZhKrOkMwCkaFJIFT2uTbxk35FGi8s+acodvFxE/yTIDwDuGGJgQtVjNH
hUxgP6QSpGgWhAiSPJbG/C+6Il5JN9tdgynscAetrG/vCR7cxeDJvbu2RTa0SOdT
YeQT/upDDdx0ZWbINO8LKlGC/M5YAcUcdylVo9H1QFZCJ7DxlNNa+B5UlSMm7sbA
osPrRdRQkEKBgb4tGAgXvoKKdItA5ostUoaHIyJencIBflJIHeadJqzj6I/PiXqm
0r+sIconfeCfu4tvN6YRH4vWbKqsnesr9I+8F+Y4ri1QdBvPkkDhnk51N4+2GTXg
VDRdJy0EY8er2uyC1V+r3YiP5zdFyG9bCm11GSusYua4UXZsNn53SAPXy++3h3+H
ijbY/kJK1w9qdlOoVF0Pd0gKyJ5HonPg33RPm1JRRysMxtaRO2oSUTMIz5v5d76q
1q6r8dmnRCWymmkzsMXarFD3ES+ZaDi35/0fMGGgfmyffjh4k7+bi4TgYd9MT0PD
z7aTKlEVkXPhaMV6fq9GyIOUuJtzpfUAbuyfF4xkeQq3GQh2XgCEFV3RUsZCpsLl
CJItSsnlyy19fsFwrpHbH5R2Wz4lXAgih6gNKaktrHt9DMZ1PbTO161HxSsYtP0u
e3QSsqCYOQ+briL+8zBI49mJ48As+Gr5JjitOR8PYtorMqJmoKSki2/rrPVk6YnT
O+KxghjItyaAf7beGGTsKHbJ9kfZ586T3qU8aRGXdLBgskMOoWlrm2bOBVeAz2kg
L1AygWgzEqUCcgCo4eiZ0xFq1YgSuH6SPBMYigUlxH7hmXUgtHSNJCK3n++fCL3R
G9wsbAmYdXAZuTuOAMJzfFSL2XwRxnKFouWrZm+G5T9xthJu1le/8reVP+OgOXZo
FoPWfwBvqUklkW1zLkDMOerfTRdqFljA0P8oycplq7TqqGRXWUEuJmNQ4/0qvH6W
3N+L29doL1OGVmkaDVWcVBby3dyQ6epJ/9o+KOpvP+8yFIILnmVmBuwNqvk6fogB
nUu7qKZglp4YXtca3a0eEsNXb59q8ByjdhPhCzAHcAzwzss0fdHQM5GbvgQ2yHy1
S7oCQufP9OWcrPunJ5PPK/2PoYLDCyLUMg/WIG/UriuPJkdS8BRf40zpwAb1rWQK
GbO+UTiqu0PsM6cBOWci2RTzK+m2G0BcWWqsIZzJ7NSQLyiw9dELOR/kD/lDHyZU
lDf/wsT67ma8Kb4JrC/YR0fIxM/gdtcB+butO7ESVOmjH5Y9079zCEWfPy7y8OXe
Z7A2K+NN2CrH2Gcvazrra9oSG9gBRWJpXgs+7ZYXaE2xYJ4JQ0Eu9XQ5J85Yh489
Vsc35CeMFrYCVfRbmDQKOAJ/qFa8R7Fl03vexDoignpce0ZVhQH1NcGJ0J4Vw1ft
9iF+J2KyshiVBEwO7Gi+HvrA84/6g9nLqwyqkC/qCVpQj38J0dKjt8/IfMDSmfer
UAHXDbHzDCLnKhEj8wVOXYgVeALSxz3WEe7Gt1OgVSy+T6D3XE617V5Yn9+66gx1
LZDKj1Oa5Jg8+1T/4b2VrU6/s8Wkco9JdNoylu/pBOuzsNgtxjee0heZ2ghRGlAp
8btdd/7xEBTRudxlFKBj24Afsd8LzF6aoKK6xoHNVoaESXMUBfNm0awWH3qmp27J
pMM9M65Kr4lrHpYTGEF8P87UUkQ8k22BAGTVdrqa7j1kNuBxensnn6Tl3uN3Q1By
SK9d2uQ8ZTk6yvh2ZQseW3Ili2T3PEE6kU46pGHs4gtDgaeV4Ek+Ldk/JIHUuvP5
vvBljMxVlH+ZK+m8fVaeDrO7Q/fY10DoFVWZeCbS4Tj9v7xnmG7kGsRdEm7Rxqi6
LfQwQ54xCxRYMeTMpz4dSBjP05C2CACbwofCbhIflhXh/I4DFxz6cXrUNDjalAEG
ZVPKNHYlZj7E3WsthUFVjHLIaLwrvhyDDtRCYefEpm3FehKWTakAg1tKtAEvoGnn
2qpY72fplPWav+Oeunf5ibORKEJRO2ywT3Qg0l1buWWgHfxqYLyYOZfbu2Kxs9mq
f6q2HU9k8vlAsglfsmHs0MLZQayQeG41O8k+hg3jzLAW57PqVStCNQoWBznI7Rtw
NlauwwV9F9ch1IP3CyfWb5zc6b+rhtoxHGa5jAgeuxNSVpdHWh8l7HOhqyydB6YE
eNBJhcW9txfBQ73iQWfQSzOML6j9wKwJEalXWXuZ7ldly7XN/7kQ0XAG4avOQKCe
T0TYnaOELFIKMbE8p49rPInTGOYh3kAoB3bZQN0CmKk2kgS28MazqcyvC4hw/ave
l5FJic/tfCJYuj/K49ET3VBPYmLXN1cW8ybNj0UrbbYn61CoOOR3P5m1Qwu2pa4R
QCdAoz0TF6UYmsZWEKxll/xJmv4RcMeyQ5bzl5xcRLuCwvInc0GF5cfVcXcJld+G
NFxeY1Hq95XaVnhOZ4SjTUm+bi9CukBpMsVcHePD94Oz+b7WVBtIKAxd11yPCF2X
j2ipLnv9uwK4mFIDb7P6y6HRnIux1SNGUh5tDCqc88wUq6Sa4eLfhYSoMa5UJ61g
23P85bpv3LEWpjzqQ4NVjz6CIPBpNo0QDr8/ptXkZWMd0XB5r7rAYVGzFe2UbNjP
LlJuc86SaX21RFwEauAp8Fbt5bRvbr7ZIytd5xK7ODlK/pmT/Oxcjee3gJDe++Il
YajvS5dvTRtZgq05i5zT2WUXcXDF4fACMLHgnxoPbsq4szVFUjpdrzt3xmoQgHgH
+zEceye9tz2nRH3Qr63Z2Km0tbYntmqcBjQi4rH4Ct1pJoZYO7ytUVbTMEHtq/yH
bvhJ5Jt3ZodhRRGKZwv8uBp3zjxicsAW/PAcqu0+dF53yLTv7aWPU487E1k8N6t5
rtDqRgwyLJiPwANcYiTPFVXWqaRhr5LykQVVvCEwef4g0SrfmajEtTRhmisboKqa
dSLrDIE49Bu3OAJdzLkLvgM/UFLpAIRjAhHYkRZ5BqbNwBMzqGYrdADv9Pm7hjxd
VvnSUGT/xTs2miMhJZpLEwxH1l8Phl4fMf8cK4Q6uF0NWkb4aysaHS+xxU3JeRUD
+Hw8vYWuUsjO6ter9l/TEsUdIQXB7HFQ2p0mGyJHeNMVMm9p5aycNzRbbvuVFBV7
bsPXflwR2jgoiOWerZliQ2adTxwFNO7lHuhAYSaJW/3WjZFg5YKPde25lVwmjCyG
H/0saf0JmEWKHpj3c2ImX+YbOFLdMroajWTydi8v4pWYcjdSUK0bGzb8Aly3+sWg
d8e7TgyhZStarjA6bizv+3W+XQUHnFPZ2lmrlhBcvPUoeOMVNs0QK/vhR1c4N0wv
0aH0KdOiauNQW5H6lCzSVnAG1ABjAI5rsq9FbNlXA9/J/w7uTnMaax6CJWeTuTo8
c6H7pfwURAfzm+4pjKWMlSqUJe0ircIt4dEbSEswhXfz/JVlUdHxP2AVNCueE2gG
T3OpOgs2Pv0VK2DgdtaveUr3TyFPZRfKCLK6jaq7zamJrcXrzm3VRAiqCNRkLKJa
3SRL9+Sn/1sVGGKczktRbGgErj/Fz7foWZO/ZsF7AY4W+qpdjVkIJOl6eVoS9duJ
/ErybvVLM+BfplftR2hRZmxsZdjfdzmUHbZDriJWSxhwryfeZaWWbfaIXESukju5
tucfeyheE71UmgHcggToO3cxTLjDJfrRuurphEVIskWHY3HE2qsWrKHZYg4Wwmcy
4lES5DwV41Gsu6YjGhLnWJWDgKweRV4uVSjPD0ciXtPrv7hJPxh24gy9YYUCmKT7
UrjTQnAIm8gKdiE9uCe3Qp4Sr+8//YxKh7rmnKWXIbm+NRPUOfuAX3V6l1Lq/FSt
HEDIFqQMuLEo7OsWAlTlN3nuPDFQSeG/9ln9H/MatstFHz1P7Dwo6IMh2ZHLleG8
jZM/cDHfwLSRxHsCIBppU6eSnDaBbVTAawnMEMlMsgcgrhCIgJz03ookncf4Lt0A
z9I01OFsjxtJSPJbAj6dWQl6Q0YQBf2AZveeLQ/boohFWkjpQLKrxZtTH6zhfJof
sA7NzGKMcmnztKwvIR5ovvijr+VT6E+7nT4QYtPQb0dnX4/9icd1gh6iJaY9SpAg
bV/ZFihYAOVyWi2+VQpoXhy4piPoUYErHPk2aO++zPHJIgXAaMJSer+Q9St0Dof3
9xVPXpjfltpovHj1z1EueRTQ9KfmPxDaH9JEXj0yPzLmSC1FTD4a8yT9KJlrjWmA
pIyXOjCOEZ5BOX2na3fbtQFnc7NPpjOWSenswc8kiGo0Mw1AMDRBx5K4ILPvhHVP
mUTHQy4c6RxLN9mi5tpKT+c4VVTEMtOVm+tL6TNrGmauvHWR6+gL5WJdoK7YSQ2B
s7YXTfhFyYA/k6kmOphvIQNhvuHwX+Z1EPxP5Juw/okufSnzi8j2eOrAcMDHy+p9
uWV4BwTS/X1ljGQyw2W9s1UyegqbpR8uwudRbmq8rbQ1aL5YJ/7iF2h6nT9BzURb
JeIlma1XEGhjQ/gR2LFY8rnEk1doZ4Oi0jjKYPnOA+q6savGNly+43KT2CBdSYfo
YLv5tMqQCoZ9ITzClch1jzaNoe9iQ4DnKHv1pQqrPopT6IJdnJUP5vph6g/qFsDx
eS0ts8GmfnF8ijNwoqWs5zRAJoGLJxZpswWpD4QKbztmG+1X3NfM2E1pzIlwOkVu
LX2sdkOKZCd9tqrs1ANOdU9+MOyHdsciSykinuQRU/kXlbi8GuLNfrACibNw4YQO
Cfyc9XBcqEjMuCXcF0/FSzEK49P+PD8AFKyinKUNHt74IYzaaT98yGiLGV4YOBeF
XlcOVUBHF3lgPXdGaDtZ8h5mfHZmmhE6JZ/xsH6VUsmfwUBDuyQC6ZSDduzR/dep
zyKDkJq2E2bdtoD4O0vNRRqp2+yZgZgfUrMZZYYkb7HK2negrrRsrWeY0CJZW2jt
0fN2+aF40PX1eQI56NKCEZDL8JtU8+iAwSzgJgyXt2sgySrUzaR1XhhPWZACD5zL
nIIA6SovNlOSXtCi3XCDgt450FKIh6pZyg554tme5IXWDnAdvchoWjoc+IPDY0Sb
U+TiCsA9wNDV0yynFR480FYpF3xTmz86SDU6gq1Nvq3ZwYwPZyNr3N/z028gs4pN
eT4jWwAUL8DbdEBmabCYKU2DNi/6Wv2P29j65INSNN7n0QnLedqM6mehn9ICAxFG
tV/hbCQtYld9Dq4B4hryOlzPMEeRPwX2pgo32Dq7o7W76C4HxIONq3lvFbnntB1p
4D4Ki5UqecGkiwkZaUBVLcX04qicxQ6OvFKSZeY9gbiUa3zyozg9LsjnQck1Mjlk
xvak8IrvpTh5v5/fscarny69EqdWCO3ODECKFUl/TOELmFGuZRz0rxHPKIVOpfKt
6dXFTuaOIxLv7zr1mk5h/1mzDlNEWqym4cfWGBMSNwO9mIwtCE6tiPa7/TulT0tl
nv/aeE1ihcqmA9rj41Aag861dQtCa/9dyTWhwqSBFOQiPLRYi8hS9EAlebaywews
f5MUsi32ZQZWAicqP8PtAuOwNu+NN08rBzNSduOrM++Md+oHd527LLPaCRJxe5W7
WKYY0EZl6sgILyAfEhzKxfYem62hp8gkCm5qv2RyK0VAhGB4u19pbZr/PyBlF/lC
LBC+KyvtXm7TiVlJEoNG+ey2gBLOpegiekjfOtSyAiTWPOLgHEdNZhRYluqs7hIq
WF+qgiJcd6ebaZRdeXQuMoZzrwHkii+0y6Tel2o9/oaJ08E+clmQwQNFxXRkK6GX
JSoMQO2JLdlP+QyDirAq+US1sBMHqfB1NmodG6L4acXO39BAeChpwIeFRU7c7qUd
Ej2xzyt6DR8rrBDvKhPkDWa+HEKv/pySY67IJnrqohPeUt4qizbQ5pMC4JjvbjYs
bGJGzuuwY7cQY6q9JBcOJ7pjwfDdkA46lsOF0q7wcRhsTbdMhXJhe6nno3p/nY9C
Npr71bVlr5DzPRT2zHlnXjw+gNRfH3zh2Ibf/GVusy5X8Qp15hejb7PRWjM3C1YK
oYZfFF72rA9Wr/4HdeHwdzP/l6aXlH2yOWb0LZvSUlqsB1+6FcvZc5Igyjm0halz
cwVHEf1aLe+/B7cLgplUZsPKbAZnOWNt44kk1th5XGpgyLSlpRuuOd800jyAvzU9
gRq18xBHM+UT+eiRnohqZovGjgWK/BzPxMSa8+nGd4C/TciI8023BL/goIcRXNJy
LRUFk4hHe+WVRkjgmyC5waPwzVC6HfpAQuZnQkxG4iAT5nFnd4fa/43/s+iLxza7
1fEeY2mIlFP15ndFEqr8NLiIDKG4UYcocZJ31autQBqeNOKWMDsp3+Aqh0NyxVR/
w9mgL4bFbGz3q/npb0HE0CZarOZM48cI4Gz3sXnuv++s0NEPAfNNFDvfkjeWzb0x
KJt89Ux1STiJr9Da3hbJ/4xjRfZpfCiRzu4s68A/AEIt6a/vj0UPETaK7nGLPQx8
NKImMv48Dt/nxubwyorH4+lgRUrT8ZFVoahxl7NeIwiqe8wi2q5lneVvTw/m2H0e
9LVvKW8XCMaI9pZIME4bdiTkxoJJtM7fxqFqnl8BNxdyylOUaO2d7fBiLCs2fhBc
wN6SsXOi9F/5qFh3uAA6CYOcvxfWqMVPe55VPzcU9R8nG0l2mhsk0/Idqhb8NasO
kcNbKaKLj4igdis/HEHrW9eBz1I8V3VkOPH5pMuv0TqJS7S2aNHfB6X6M+TihZ1Q
W+H9Odq/gmYmJkBLyF2mwDK/Vw0iO0MpQ19jAhtsO5LPBd/cUhIEjKf3kcvQpW8K
fOBARNGZdyDbPqM+9o/Zy4hUX2d6SKZ8kjqSee5n+YpD5bMA0xX6W86F1RnWfcXe
ALWqhzOQmYcdgv2xua8a4MgnOP0b96DetbbXqjqL9I42S4Qd+Um/z0tmAEyjAnxl
n67Z5COSzuKA1aEWo471OGLozzIVEChoHPtyC7ROXnLbdMbIY87yKLZ6y2w49zQn
Zq7VAZb+/RA91E2hBpCtAsh8Yqdz0r1mlFlIGlWD/Pb29/qwM+eeQ88JRX0fZyOS
A+Bgq0rgr0ItGoJkuZeazmgEgWfI/nuj5MdK2+VmbVCDlADmZwX6keGq8tap3vLu
P9oNosbERWMDBfK7D8utHgxeXXG+jgHpkj51k7Cm8RupjQysf1KfpHNkEpXwWje/
/GCbZlMTyXmR6xIIIodPMNMOj3iGgVqIrZwUmBku9UBJXZALV7TVL/SoogDh1Zl+
MuISxQ1S8jV85+qYL1ZzcNs3dqpLsWjBMQvaqN0lJJ9LZDMHjIsSsRVjGFBkEUnm
9Hro8vUSksNH2buHiF4GvZRsc6bVEuPBiTh9a2g9M2SQEd98l/AoE2qhUiCo5OSG
+numjiVqqlPcA0NuBP1tgPLNIuqZjHsqGmbTEDbRfXnaleO4cwOiNDq/DghGeBkM
Bs+9awrAt58gv4uMoqpebZKaId6VW/cLJGUrrwCqaJ4fLTCT6Qe9YzFefmQmSH1k
X+lk3f6t/l0C3P6nKgRXKKo3wf25Unq0toh6DTbPCTyxzMuFp1SQxb4JaSY0kG/F
8nIct1i1VGa0nd1TrqQpc67aiP2hYV6nXuwVBZPRzeN2JE7nHcZet0aVI4eRz7BG
1uDozk35/5PaPO/qqQZwsZ3LuVT7a0yXmmSrNSt4yu6byak9vEJ4phF6pzKoNNcv
+TdkSlOD5Eo5bBY9evoF/tIy1q8Ksi2D73SQGuoRJ1K9XFN+Ix8ULzqMd6IchAd/
xe/BxXI3K2R53EXLmuLh5gQHWIXOhnLoV/eTnjj4NE4EQhevOQxFz7+crfuYkChc
Eo2BFAEDEUnqJuWUzpc6MBK5uG8OEKi/DcnJTozBl4veyoron41wHvOJyxV/wm3P
TMBvEn92SZkB4/FzLhErXZxrJB/ObJttbLAC4fOXqYfgLoUKZDEhRuDTh0MXltzf
tO3YIe6seaUKxIZtD9193H6VHR8DTg8G4oImRRZVsJfM9byUwJS9w13faELgC1xu
D0vUjTjli5NoEp2yXzCyWo6PbwogCq1+V823Yy8x2hIQgB0MIWtmzMpOBuUPdaHw
Nde26CwC40j9G7L/I30xPUCo3jHaITQzH1w9xrRAGDqglG3n43ffN568FCb/U6ww
lpYFAoZeBeBMprqxpRI0R40BSvHa8efGza5IKGXDHbIrqKzSS+NPCjuaNmsZuasx
40hde+c6PT19xakDk2l2C3P0dbSpiiKLXtxkmvaRxiMffBOvWDApHORu/+awFRAP
O/F/OvEd5SXqyCKHeM1oubSBWFDifMmGw+IbaEnaNM5VOFnyOO4tb4XlrMzTduuZ
sL4cnsAD821TScKxXlPu4uV2Bwr9Te8Em6xOCrj0JqVj/+wDlOPndx0zOnSXGPwF
Ltb/Mfsq5m0nxXHSSO2bdi6lWXH+WI0kf2AUlMV3tFzzb0O+KPP+gLNk9Qze40cB
klrkxO66aXGaWcnQytgfOQEsokXkhFY8r4Dnn95d0WBvICVJv7NXzQ7Ss8SQ+fsD
SVSpqjRNwhSE7JZ8/b7pD8ssHixgsGM9Kblt8sGHw75ZqCrk9inXRd56+aN4Fgae
dIlW4xhNuCJ9WNdG9Vqp9WA9JwWM2KHMQfB6/y4iTIzBoaAUbGBXFwMNQBFNq2j0
PRX7vVJuXxACguUUm1f95th5q1Ya8a+9yeh0DKecmGe+oJ3kYh7YtT7ybCYtXjeH
R2Pprf/zw3GyO6WRF8zvNll39JUQtnsyXK3HaWelPiXwusHLWcaMCbLdxF3Dl7au
Jqouu3/wYwpiquN5EFvPNs0qYUB0le3d9ZRDA41JlmSHKuDnI1j7QfhMdSxF31H+
HsDhiMU0SkIWE4V8RdFeo08DvUtDceh9J7T+NY+bMUMXxxzuQWEC0ny4tF9CDsev
fShPGwS6wyXVKiM30lRJPhxeZazEiU+dyk1DpDqjhmyB/H37b8q0iUuhIVf00TnQ
f80FExNP5njlMvbZyNIYqUrwzMYBE7FeAXFv2ud7ooOJuRuFg85trrqpCmUlGeha
L+tqKN/OIx0oTSqgLg4nsADBjPtd17ZGBkm/Lx6s69tlD2hmuwGmX7tMB9jUAzJX
mzYe2bmtb46ge/6R7iJF9NDYA74awPUKuqUT01y+WEo6Wk6foeAQT2WbMtWaKAl4
5SOAU+mt3QNMj7PFdY/0EHzTsFHjc6HVVGH48wvki8dkxCD9/9CSLumj++YJ3CZb
G+Mgr0GT6d4TINCH0al+fgGJMxhCnY4cJnwZXCIDJkNcoD0yeC4sKMG+YeTTg7Pm
doBLJDS+kbqbaYsZ7AOTHN2WlDztMTd+AyIXrPyNihdJjQ0aXoQbswwMyop0qeRL
ib2fzqW0+kA9JU30yZasQZN+2qOfE9bju0U9mCTEBNMY1l2D3qEVwhgzFy/v9xUJ
qMuOlm4wSwuGy23B8waAs8kiA4fge/qCqIrBbWPhOOQbtFTL8RWsbt3EW909T6Xy
bqrPCteW0ZHOekLGwqcPBhc/SqKDq4tbiziJutDzYO8agQYR9xlWcCo0l5bbMXMS
ewZkxeXZ1qltVWWuCC+0kwtW9SErRljJ8245ZyjFeNh0C1ETu2LBSFLcWvl8NB0v
IZIBZju/G8oIKXheHIf7pYEnjFHHYx6z4gG3Bn0LFiXf0G0izEwTxhBhqXfjQtH9
R5aYHlWVqQ9cw+vKu5nlbzEvMGLtbKVvYtg62X2pwsO1tWH5mccmEMMOkDEnhzAz
2+qnLi58spqDWOca6zM09n8AyyAB6VaLHvGzxotXQ8ZOEVDErAV8C2VF+QP4unBL
lviACdP+PEz2/agwA9d0njK18acyIOO6igTn5X1UY/EnyxWoaw9nqWlj3eg/Urfi
/eMS1afT0TY1cO19BXNPs870NGrdijcYp/WY04V+mxLHRtFc/Wpg3ryqcOdafgI7
oaEBp5zE2NN4QfsKmb/Wh+MjF7HfSI8GUEOhbC1GHL4Y376AJz+XD21pXpHIPWaD
KUWZRZREr/rUSQyG6VqyY9wZtflI2uTB/dLwsIkzfqqr+54ZnHwxHnsqPpth12lz
NxDj3a4++NhNtmNv9Ki+HHlzKSqTdjUwNMrv96WPMb+vH1B9BP6FENjYyGa4ZJj7
4pe3Th41l3nuIDnsQHQtmkquYvk1c2AGW3soD167a1XOZD1IwmKf/OcDwm91lp+W
Fdq1Pb/nu8H/YGc7xYnasJvbM8QIKV1925jz5bgkBzygGPqm9+N72dbBCbyYuXiv
o6jzj4P5lGerdf2Vn22hzcKlbkeVv2tJW7Xe5JQLOBBIOs/8Ccltek2gIBiR4ybl
tZ7RVWDpp8bqXFPpY8J02C/G1Tp/plBnvCf2Co+zW2XyewWdOkxEcbw6FXCFomM1
2YTxzErbh8elfuwjmiquW6SWCChPf3Suk0HTAfqTg/WN4GnRrAjDfO4ujmkkyhFV
no325QEdkKMV3C7KtfkJr8Xj1p4Szc0JCGDDz/JvusSet5JW0bG/J7zHugaa9bCV
tQM4lAOBUJnTqvCot11huBB86YoagDVRTdBeGuuMef7LLBuImaduY58p+TiWTb5R
+xcggQpuBWZCzqeW5ZW6L/mBM22QsjKMROgxORWGVfjdxQEgVN1yQ3BteL/l20QB
jghCpF83zr6oEbNWOyP/q3/y6E4AsIZD82iMLvvys1EOpDMhl2aV6wv8WQRJ3n1P
m2zmEoBtMQ09LQejhLi4c/cJx80iu5cXjfpDH4rsy6KEB7yjHM4I22c8ehBuMEHC
t1EB6uQWJ/WAKzoZt6lXno9uHMqpELyqdNiAjf959sjEk3Y5lKd+x3JGQAO2J+A9
X03Y/szCZ9J4FrUWdpKmeDTV1nShfPTUgkhEIbfGETx0Zkwwc9q0oH9LVeEgiVIG
V7UFHyk4aGNzSt7R3RRpWC4eeE2ogQZvPPGm7lINcY1zEFRV87TYkBnD1KD4jlqo
CCbSND4utzCFbTESWfeLNwVNOIx6Ym1Av0o1AHIixOVZ0dwolSR/F8M473rHEno2
TnifkKBzUPg0qTxBj1xaMDND05eeZ7KXquQ7ADUdxyg3sVPaN5TXR5Ou/IjTHwEi
ZWcMIuP+H5EDIBTCmQlMBuE827y9zK2uDoJrz1vKl/uw6wf2Q8gMB1CIkZiza5Ij
jtyMJu+1Zg7FGZ+dsjAfMF3RPmTFxyG6NDKci8vIkrM2loB+9JVmhdVtEMQSKm7+
ma+Rv2c6cg7pj3nrSJcg99lgr5vXIBeUI0OlV8wueYhs3Htk/Zyd4LEiQSD/FBBx
KZkqCu3V3N52OXWrgj/R4RkBYsX4lIfoFWd+OeInDO8e0vYvehTjlfaa4L2YxLZC
e9BdtgZ32amFWD/TzQbut1xzl7eAKOqBtocU1fDJoC/qgrG/GOwcbhui3lNQ1kss
7QN4gs784EYaFfDTDAM6GVs+FtuYD2WBkNF3kx3Vwz7YfYasUxexcrHM1vAFJJ+k
y2q0Bee3d1GzSGfeXJsdLGELYeKpLT6+WyDkf3x+e754ymYbKf9OkStwJT4V0iR8
c3OqkRHULw4WEHfJKPVMYtfrXmKY6rHZna+zXxYeMyiphYT2pHwir6EUxa/AJW82
Cm0d2jMncGS7xXC03ooh5jGCMQHmPgAIVcmPO/BX2ON6f9G+pcowZbTA7NhSugLW
uwGunBiA6C2Hsns3yVd+9WIjGtQdcBnZRfNNeLoyDSP4SFbHngZKZlJEJCvbWUmG
CqlRXSuxAWOEnGFbe9TY9Qdgz2k2ZpOTPJg1KRnFrRb0frrL2POZp/377hlFKh0K
7LdjgYNs0PRK4Q4nnThKtBBKUInhNbEIy+0GDGenxgtWIj0M/YJczR4GpCnOmVBe
5HF2dfQFYq2oFDKbOtJxpZNhreXIC0RWLGu5qX3h80UYeLosmhciOZvxFD3slAIm
xCapUusYNMm/kigDDMyG7+napcoqaBG3YAQ7Lypbhjl1FPnTwfaWndIFtZDVfYId
z/H+6k5MfcEjohFHT86gYK09HQ8wcAvjhKBwm/Q+ga2zfVmB1UNbgpJakQX9a+1N
alCbeDnK59+fKhZMr/rZPsUE4qG94APdF7EbxeZGw+I5XRdXCrdA/9VVVLYgI9Ei
LaTcp0it6Xz4JsrsuwxZRp/bEnqnJ+NQs/3BGcLsHdR0ptzsMZUOcyfo8l7sbEcY
VoJNSdzxgIe68ewHm/QU58shGk3Q1hhKsIsLTOzvXYz4POFz6GSCDe78ffmMO54y
7xXI/BGOjB9AbJBH8yiWmMoSzsz72cGUqFvbGfk8Y6khC7rgXngdfHEhIgsSVYFk
58ut2acjwBspt0GXuKo8yX5GYQRIzflAfkCnEBMC47WTWjWQH2RM0PVztGMnxCrz
Yc6CzhR6t/O0PMKJ6Z47dlF7XooOih5fnRFM/oa8yMqMgH3R1AO6g2BZwqTrYIiR
4gxTquAiuqrsHC3VAt9HkRO/nNHLIVqc+c6YhmPG7J3+vrXz8xxTRqj6t0mirVUb
NxE7/gpWYTQdZfgheFz7ru8TY87IV3UvVeADu86SK7Gzlg0PYIWTdRSNlQqo0AOv
ObHF65kNLI+A3nZsqXHmNd46JumeY3Kb6S5vZSh603Q89JSC8weXVvOScaffmGuk
R4XZdMYtZjVH20nSg+eCpnt8HRY3y89H8PYCKIvDwM/ivBzG0qqYCtQm7MYuJovY
gG2PXHWz9kCSpJaB3+zfYaUIPfBRUZjeRLow4DUy42lvsx6M2mWNdB2KTYA2cLZ8
813Xf/rafhpuS0ogyBC6ydUgB3RYhEKOJz34MJmhpb8VtUSoNKv2BI1Wfe9ZBsVD
5MbQxiEKPNde8O8G+wrxkV5zsTYbmzdRbVR8+epW//Qo6/FCSCc6v2LRwSlAVhnu
3aRc2NNGKgKZLLve6N3R9NfVHbPq72r3moddVJsAFqJlHOitWb2ekjKgNTmLB+SM
xgazW44oIPy+S4PdEZI91vuE3lqnhuDplI12mbULLUsdJUOGHJdJVw5qigypBvD2
l3zfD0FTeNzEbs2mE/LIyr5YKnrZu/dG9deHCweYL9J9xEMVWvhPvsdUHUecmiJ0
v5m9S7b7dG1M4fGG/F4BXT6/g4W8vMfkFk+hQWegeGt4UcvVFVbxvtbap698WAHi
BjS0Dt7J7Oc/ci16RHzAhiVFCsIbxfkgb2QYBQtuj6RXdykLMVF2yqMNPN4Tg5FB
ThzqSNg7yc01K2qscLyOiuiJ+AZGaVVY+ycVJMpfmPdArSj8+X8CYMca3+j1lxot
kzuIwPVEWrVT5RiNPZU7EMUD6WNXljbU631FVLO8rOnfZbM5JHHfbE/jwwovYj0C
p9hiwpOWUxYry19ZQXEG78JGdEj8CFf8sAmGVnv/TfCjuNQylrX3GFbybYBWnvIy
m8egfcvWPeDVzq+bR4l1TXZo8TX1MtQN6N+sdsFF1XrXKb8YAcdbZ74jMoEy1DfF
Bbym+m1deCvMM6TWLvKOT8Lhl3t5sQbveta55NbbYNt8EIOPEebP8ILTPusZ9uCe
iLrpoK0U/tjp4RA45Hng8cxeKKS1KxQUjr1HVv4ZMv+A6ik9uQHFq3BTLSEeJw80
qPgdd4R80Gyh2SOlhsHIftw6m9kdLnYmkM4wjplIQb4G/NQegUAbJUf5SNDKc55f
O6q2WhFQs+hTurXnBKe0NbIdZgrhSylE4cE4D0fRgzCjTdGiQzzgBROHhL1LhKFR
KP84jMe5+gy3BSBVuLrAQFvRKloafKuOUxynznSamO/XX3DZFJk2irbEhTofnFIO
rdWxGYsohq2fX81s+5GQb7VpCqQsADrINBxtqdrZv9CgAM0BmNRRXNGt6CcMkzmW
7d/1QApbc2FOkWg+LPwpIzTYJbX/Jlg32w7kXMaw0scm8b6WVsUXtiJScPJfk6Gt
2ylgAa/mo2936paSnYcT7xKvIwXWzl39Zj+/628jxEEsnz/ex2GKaoB8kKid5mBs
B5xB7WM3KcR6UrD94vy2XRUgOWD8bghX9RmxRBe0hOcWIsME/eRQzIaqh1qScq7q
DreiLOV0vv4klsQpflcOJz8ExNAGbwdYKXghsW0t2gHLM9t3qIhdcLkGKgO7TgFz
+MDXa/OAHO5b84wzjttGj3+kI6MSINGtMp/U6VIk/I2LjhZkHmq5Bi0rzweRZaGy
o3wfbU0azONjWryL95u+aFosBQF+oOPo/AJbkcegB8Y2I74uP126aIdNN/KmimzC
wihvFlfoR5imLzhHjYRhpzcaO/NGjRmSQmUxpYg5+zzFn8l79vOuu3+GZV5jhqS5
LuVNPomDXbN0yc3eVdJSpKmO8CUS4FH9tZxnYJUuskTDXyIM1eBBrrwCAotjyxzz
1msXZlIRNKEp7g2o+rJEnktYKCSmU0ksl1fZngLtiGNcIBj42sYtibfiqwD01Ovk
iik+LY7akF2jkNEvZa2K8gWVnKjO01eHTTLFW5XNKzQZxRHn9vPll9bvsiulklKo
DRmgG6+fXlXRtU8SclzM7GwAMEiI/Q4USZENP0wObBj/fE7d3XFk7sfB/gtFrtd0
LsVZyNr6heSdiM248idX0UGdiS8Zi7UAh2t+Djrj6HiOlNUJthZ/3lQBzgS0LQWT
q6gxsaG3Ah85RrwljoIvGneBIk7oHGlpuAyun3gmmv1cxxNCs/wKR3BtcEVGbf0F
BnADq1YjkSmylRhjBA/dxU2nNoYOHt1TwxB8BYNrpY/geGVxayHVrGVx6xOkmRMM
9dUXyLJYHIY+i+e7ymeVul71zWrj1c+ICsL5IJcph9wHqPgcohUoAONMnWAsZ7bh
IIq/+BrCqyBN4g65RH6oJ47gSL3ptk+rkNU9lTges8Cj3R9H5FlLyTqv2XwaVwhv
KLx204cd9EyxaCHsAatfyLxj1tP8Zo1RTKipp23FGhnKI7AlWiVT9saKqpR1eWv4
u0VLJEuG15+aBTDiViaViU5IKQuajwqBBsSTgMwzlQm/ba+BJaI0Q843XRaxlw1o
ZGd6gL5LA8q6cAQVQZEvun1wu43BB+plofAY4oZvSh3RXpRWgfbmyasginFLIEff
l8IzfzC/uehMOMXbguV73Ze1nnNs8VYxxpQqlRkqHqeGwO8dhE2SASn8RWhJ+YTO
u1g+oOZaQGv/XRfTSTDMQS2IOAIZjE+Oj8dtr6XEfHElue4OyKIyCPzYYWXay1yg
WzIXrf+0zdIBemkIxFPaYiXeN3KG6Dnzt3n0nEVbs85Eu5iQTN/ounBR7dNUPtlp
tDWwRlTozU+QI+nnwrZYQByKFrU/7rmV1S0LvOO3v9X0G2mZxCgvUMFMqAdKIB41
GnQJm8L+aCeUf2awAkcL+WhiotKzhs8iTr68TgvLLPwbTvc6n+YwwLZpAAQ2nDBE
edK09ZAcYE0fTsZtLsPsHRdC9GkOof67FpHJ4ouMuqMw7uYeRDLm9xuvEvmpVJqM
UFjYlxHeuKb1cRE9R9a6EPHQVTm4D7TWOCLkLEv/aPM9NLb8NexWhTvVm5EUI/iw
rYhjolSt16bFM4KvS1Pjm2F2GKkijSxLyok7C4Sb1pVDxZpSdRduJvALCZ8QIQyl
z4KyALl/96Ov1+63XolYnvMdPJ/zxqPiph+3dE00/4bthcrFoDVarmxwDWdd05cy
AsJULX30XItl3Mrx30vDuVYrLPlcEF3pWs73yV/t/fgf6tIj+TvNBliWRSI0Ayaw
JOqxdCf4iD/DAXtknzUzAj+hzsuUpNtRPhTS3I9VmVntnnqMxVl0sH/MMjuG2aUC
65aTqITU9uwUuxiFFJctA776CPl3eI8D3b3aww5ARVuY7xhnVc28QyR9izziLXV1
w/LD6u3LhsU31soVsMwaAXULCS8mGgYS+VT1dYbfg1UnlycOMgy1T4PmKAA/eltW
1zld80UQVP5RgKmt++eucceOVWawIqi98ou3LMEb34nBu2NRfRXegeREzV+37hMH
BbzveWKMHk5C1SXKT4O8IdbEwW9B7iVk4TFlE7z/EvVPRC795dciaRYJ8JijT0Tv
2a8mrI5qIlIiF8wHDd73xedBzAHtXRhVFn3dcwej7VdNFv8+S30gEz4iT1Vtvc1m
qgwXTanUakqx5vN/pdiEuADT7csIVxqm+Ree8Xnqk/1rYYCM9x6/aOTMfiXTJmQz
X8dIJrrE9FOVx0/gEoDzMEne14gXqVazxnzTTcIrslsDkoNv7lYXFPgOKQnPhKKe
4o4TiaKwGa8vWsV7LHGXZydtEt0QQ3Lo0zHKHeq45A0BZWik1mRR2kZSjM6oTQ5v
HGioxt/5FUNqc8JGuv9/l415vRMWI06zlVKWcutALMYfQN6RsgvftrO8SEW2fjGO
7mOna3z76bs2mVh5ZNvz8U4bmV7IVjtNxfNEjR7nlJECwMuaeAVznJ1cd/FFfuDs
3NkPzUbDvQR5DbzqV46Tm9bAmdy5QHdTWBMztxFrGVOl85d6Ce7nOW0DxOkdvIPi
k3mJUFGMkr0dZp3jIlsU2zsD/tpUQ9RyDxZvexLdzl4qgmBF0OZWZ1Jtym5aQSIF
HSH8CmfwbEuRECEzlFpteH/Iah81iDac4IpdCb5zwzUty9OS86Ved7Qmov6bdVaY
pA5whLGXPtl7W+3PQUsQLZH+0NLD2c/V1pT8nxvvwC9CmGqYuv7zg0fuG7quUYbN
N/jBUg3RYZro3ZaFbp20qYVoC2g8/COyA5AhFjMrQLzlw8seJKWEaxoTYJF3c4+a
PPKw471ynS2E+kHjD0hchkFTpr1n/EEchlex4rt89WyHsHXa73FMpIZOe1QU4fHl
jjRCxVz2nH/sMRxeKjkdnOffC16NIKzU+EFrG9DBBaQfRU/GP61IC2by8L8R02G/
wMaQ1m2TOV9q8sqZMvam0WnQmEIAoxY6Dfde+nb2Cg3Or9JOijjWeLS4+yDsdc+o
da+5S4gtaGatCXXrJOmb/Ge+IDavbTegoC/qj4VW5AHopaV2joT7/1z5yKZcrR6v
HEMJlk5S0H5rL1ZrDHm5/lgX9RXycZTCJMvKPF0P2FRS/t9MpMilq0fa2zLVMQwM
TZfvEwSr9foqYa+rw3ahuW5LxjqytUlGwNKxqb0/DylK9AEGQgcti8rFbytU5roa
/nALtY8AkQKsCO2hkcErra6aARMDrDSC55fahHX1fk2k9S1CANM377T3K81BBSoQ
DzIVgi8qJ6uVtL3LmBUb9IW6Emw4Wd/ydPEZgzI9LEUMD1IprcfUt9smSwjL5vGK
3GPIu4ohkBSHh+pJmOAX7IhB/SH2bKjZHzTtVS1F8ATCGkqDCixWMQ/BQkzVAy5H
5waE1P4TxPkrQSzUxxrgBirz0ZoyDY+d5HnHCEVw4KV10yWnmmTOuoIvB6YxAkil
IYQW94B2fYm8XRTPB5IAuCjG9Ff0eJ7ySSnuT0cTrCByRXYp/7HrujkN70oAMrO4
5Z913/js3Vp1C44xYzC9SWguYmD01VR2mUya3h/5vwvKEflnVLPan8lhIIaNoUb2
b4NqfCxtAAmTnIvnaJdSZSDnMUEo/qm/ne0eKKZoWJMvPSR59NTmTKI5HfUokgaG
MyhfIY+RPyiXSF8kwA7XNPhLzm32nw40F1ZYBh38W6UqagpPhFlqeoO8EGuFEALh
S4KFg7aUul/t+kyxLiM70GDs+tMMMrjwR1lXQHpCzqLEsl5ZVHJGQyIZ5yAtRyrZ
r+eGHRkimN5jDmNFKSbHaz73ac3mULLEqxJVup5oFoHLyoBo99qYScBup/0rwNZQ
hJs5Q7vU8qaXh7V/pwgVIcrEDnJ9zszHZL+Ccq/tpwCcudKF7QmfrPgMCD9ZC6oD
h66vunWXCd0+U3nj14QKPvOV7QSnpYhBsSmwHQXNE5PZTO9sx4mY4bpJgPmDMqog
MNFQtfPKkoTq0ZEFALTr5Dx+YNyKMAhAO8wgvx0FNl6xwHfPi79zBKKrD/HYcfsx
Us5gW5scBbCKr3MdPeUWikOYjc/FhDAGV7ov8LPcS96mvcIJ4GQ1SheZg6aTwgy9
HdLAz4C6WLozjMiRSDsY7KL6KrtW6Y1jg79iPwR4q7d6AmjoEZky3jThr4Qos7Cb
SZBu2CICM3wip6QcPnQwShNoi+m4uvV+NweT7JXYI17fk5UL4FEYaulwxpWQFQW8
KWhQT8x9tWAMi5YKFgOMKoNkhZPReJ6QRC+gw6dXC9KvwiW74+2lo+7kSuwG2cbS
ZFcnnxqnHQEYgIVtokofENr2Yne4YHqFKuudk/uiO8VzZlRdvTAdL73taWPIp1RU
Ano44YV3R8QYDR6UVSYUgN2S+tjoeCtq1z1a9xr2maSlD1mB80SOztfmZW06Qj8k
2PNnMXxQ9IjgdF2Vl6fsE2RhDI/3509VlFr4lvFLnubYDvuC8+dc7++sa0bys1D4
pVi3cFr7LkC6UBlt8qZ0tc2S0Z/jXQEdr+E7eyjSei9RFKfOrwKqmTGoI1rlKACF
ch3q3uB8YS4EFjEJW5QctLrlWRWA+Ax0rY+SAMZQEpVDdINQA/FvY9t65xOZ4h3q
gq9DQgMCG1Ug1tyqZ9/akjNWQxTJ3IHxsq423vrmnSeZfLtTKVz4LkjSikxKMwKB
w7biPiDeQhgLyvRhdL3Z2TYrHyFbb+xOqc/vu60d0zAY/bTMYRSIs7d8lqyaFjDV
UQUyZNVyj60m1RkX/OHzvqE+FdaVaaR23nHTnFj5542UtKj6pENXJTFH27A/xrql
7g6IL0ebjtE2dZclEyL0UvRI0FvXbNlsJLo920J1QmMg7Je5CuRwjguY0fAkJ3Gi
Kjxb5R8wF8V0daXjELk5O/fp7kEj0Y5dGEy+w5ALQz1LaxBBy1mgwgxRCeEce90g
LLUmNSCygxsmJHWjoqzgyajlM5HxefgvloONa7d8eOFwytZA46q5U59VUKZywLtr
/WoZHvvjNTPG8aiHq8dMccp8LGlaKD/0o6SX/6pXY1blRgSES9k+saKiaAlh/H4h
q1O+afftisUTFj+cz19FroGeDEpbGWHKLX0by4QcsagaHo8aD87yGXKEv9H9qI7O
p9Tic8q11D6j84AGEzDqCrhFJbyNYMV8s+dPoFAcvP1Cua/CSa0kM5wTyCdNmaH3
yC9U/4ad2SU9YDfRK9iBwcmUJvFa0zdzkNlR8yZW3pbWOv1/OHR8Wr03/EUG+M1G
3xgdizx46aXdyz+QpWp5ueulLvs1irS8Ttcq/TlcOLUyhl9ugT9TO32ZMN8vqbFN
SEfg1IXklWVJ5dAvHI9JY+T+dZTmxxvIPled1L3kSiYE3OhseRyxy+b7l8rWiK6I
pD2ggbZhYQFsa/4zzfZ1zrd6ZoNXQV/So6CHhzBiKjPrydZxZfgNyj9m7ktlZbmk
SkKQPIDDYVCc2X8EPMADDmc27YC200/DQ8p0+U/XsFNMysN/DB3FXzAYv27mVgOI
Fg8HHJRWhNAaA7Oc0sUqiU4C1SX8somtW81dPgP2LO8zj8pIhImncEqsd5JRPxdS
LRE2TaDpLW7u+kPOhImSlhQXgvDyHs7PO5Kpt3gzSvZlLkXDmPIx0Ux4CXr9CoUA
0tJtgP7zZ2lb+ue0vNh5uO6smSUglCvV+fOhbUlxcfxd6p7lDn+vFHH6qxlxNLe+
VVcd3oyjYsduniDdGkO/RFO+Rzso9qaL3gDzlB4DpYX5wthp7CO0R4V38JnK+N7l
voKcJ/BnzrCJviTu495yo5ZcU/s3ztn9LXsugB5GwbLr0BSs2ZRHoPGI/ochOdgI
z8da6PJ6ew20qVuKxkGJf71i3IS9Wk5G9d4RYe5Dmg8KkoaRnEF2x0ShitCIC+7M
k16KZb6aSMcEp5KeN6ofMYaW26lCF+l0YA11g+sdqlMuGFJU2FqPhodFkpQX2nzk
HB4gW/WoKOa6xFpblBp7CD4rOu9p+hsePeMwCoeLKvJWIkQxaAH/QKJtxyylF6aP
wTm8n8/V42GwyzEwAmIIsu5ZfoKUEby1Eu/O6bYXXZI6Hqu/jrzcJfB8UGPwo+Pf
PwC+WzLyA7YnV5S94pD11Tw8UFRcXz5+31jWfer2beP01x4Zyp+U5e3l5mVoUb2X
5sz6ptk1uFDYnkebFsb9MRWvN9138cXV+MgjLvC4Ys0l5kB/8lGDGwWagbC8BQnC
tcgcU4pSZ46dOfV5AMdzo/JPD1uAIRebNS/Y1HABTFBvb8fwhU9kQz2DTTmuj2nw
+siyg3IlRlLbEi5zTicCh2VBnlRpPyGHymkR8JgeEN3RuB7B22m+NtxiPQDmlsY5
Fzbey9ow1xWPqLGLQ9PlZ3TLM8vpk/FObyZpyuTzhqUUM7YpCeCjiz2GrRdqCDwy
LMdSc3ss1Q27fv94b+3ExqHp9ZrglVpNC5YDnEgNVU9tcDlmfILQm25Z3oxyv8Yt
97TG/QjAEDuuM8BL4FdSuEH2PDyi7CbzEDi5WXP6GtNB6NAbyLI3mCuQmDAppu+E
dmvEvvpsnjzPlKWbmxhj6aEGVzMRuk+hryojN8/2e70twhT05RT6kStxCbAOvFhm
iWq53+NOf9dO7oQORRPamtary0lA2MXAKdYhIFKEF/fHRYuFyV1yVeJt2DY9pzS5
VQl+hNXCqZ+tXybYTqCV4pKLPFHnq9ovzEWmKKpAIa1nEUFXTq83rVsz2GhQ+ZJp
dQsemLhirHJCjDXSESeCvLUOhU15Hycs0PPeqy2UmsdGyj3dRvgRVU4Bz8XvMbg0
wlNbFQSnm0JErGOAD93Vfbi56uGOUhZRI+0+AA4x89UsMmeZC+S3IaYTP4IF+yHx
Wv7EUzObBxmWVvBrW4cDof5nojjV+vfSjCjyZTp5FPkas2kIdI8q3rbgELC5F+Hs
nNy9CWnURhMdHIUG+BrkkAG0SHhz1+jQ4KQTQuWkCtg1hmyKwa7XKnndcSo12Q+A
nSIht8Bu+LgJK6JzL6MLdGKsyMMTKWeBrqE14Bnq3QXtHkYGrv6oiaRRmleS6yGL
VQcGs2t7Z0yV6+ZQGNI815/sEwVa9hGsqlYu+W26GPdipo7FKKhVXd6rl1PzxWCU
b94yJShSs9UhDolB4KeZwF1QxTJtna2nAnduRj156GGYtmrNMjxL2717TSqN8xv2
2pC6EgqUFpepVHUmov87XrohrZ2MAzSYCMehzs4iCUeeEWyRtsF9cSJcK4e4SzD9
85vZpwJIPRRwc9GdnzI9S3XAVUVjRdFXFJN26qmZorey8vWdvHFoJJilad39a04u
jI47XokXYAz/ygMvIGHX3K7oZledLtmL6sOgsGtbM9dqAKau11CPVg+Q6FiOfZqv
2Jr105db7a/CjOhrQLUheHiD8S03lk4Tx97fHKpPKa/wFs9x2kR/vzg7K+4U2YLu
K/8zhZ0GgKcX/WDJs+C49aQGl7GOF1yDi/10i4w+XA1XXgO8qwgwOoKXQZfQCEQ0
nF+Mlbawf2ybPA1XTXSi1lX5ncdRZezkOKt4uEOdC99BC7ooXAOR6x275xQN6Uft
VE2OSy4VRANJXCjiQN/l950ngYkWbqza2CosgnTT4SkW73EzNLDMyp1DXNV1T7F1
InCSFpg7MeQgLKAk0p1QsLNkSXRKtTL98CFblX1h8Asj1wrmIeuFafS1y2S/zbVf
7UrvI0mGJCBaBggTpmfalK3aWOf3g6r/45+Wh5JfAUjqHGxD/ARLoi5CoM42i8n4
B9Bd3Y/6QEC70j4vDK5J9yEey7HcYKBL00vq4Kfe3/EVGduxbHZcwEKMR8ti53K5
HOdtJJhxrp8e7IAJ/dP0NEVgM0kFl+qR/RVUROcf83v54LATj2w+V0TkzAkMyUpO
VpNivppac847rt5FmRnrxWzShLBYvKz7J1RtpJSd/qbmO4upgOYJK8iu6qxBxj4Q
KxbXkWZ2FCgcBOq4AGX1zfADclUxOrlo5LpI95+coGdRpQSxoMSTj8OKkhupOEfo
i6dTjTeBSofjGrGpuhc/OmEKuly1iuj9ZC+XtKkht0ORrkNff6lqfBSOdnHZ/z5o
5cRitgpSOzf6CFeesNbk19+uenudlgBRfQ/i40P4yRf9ciTqX6NXvVhui7dMUz5e
DJhW+soraIdiJDgFpFoDy3B++oY7owUIUXhyb1gfSC8hN/rqI36M2kPZruDfUuz3
Ipt/3hraznuHXvp+y9wuGQLRoKYR1GtTB/Vte4B8KDHXRz/2H2jcF3cSE0xpLmGF
KVkVFmdsQhdpWz8TWQxjiM5GP7Y23ibbDEr+RgUu7rgqlP62dcA0Oaj5/2lnIKTt
8QXoMJ7Hyg39YYl6FS4YCmelDsDbYIah8stCZJOw/sk+mR747/1H7oahmMIXFp1R
rKwIFna5mb9Zd1/6DQo+QUJRC9K97N3Ns6/HdJCDYlU/9DGXB5o+V7KTorRTEESA
1i37JvRvXSPVsmgvb6fA+ilzFaeDZcqhvxd8Znk9SaMQ5omMNURQ4TQdgsDrELDp
bG3auUYMkx4YIutZZLE8N36Veqlk0yovOL9duYHd5IrweNsaW2LNZRGNGSo575qD
Qafu2mxwjgWNGV7xkXwScM6knzuLh7MDE5UlQrzB7lkUqIivU0uBAbquCBCGNqgc
VPgtRFhkVpnexx8NlteuDNknM/eEeBOSULu2mmPKb34AvuJJ6gAJiqGP8YzBcfwy
zZh2rQ/XN7ExU3q1ug5/rxd6EUheiM9m9iW6Z9CpuPVn596ldpSW2edD7ZnmvPdo
nDr6XXRNsSmipa8uTFuLjrS3aKvdw6REhnTUylDH5sp/LQafC+sFUY6Zj4imnfXK
iznFziRW73YniDM8QWxDKq6mgI1m3BHrqXHwO+K788VoNiUqqh20df8M1ojgnoEQ
aV558DsFk6CCUydI0P5rDOhAPFbEREg5FiWwbdbyJQajSfPlU+t1Y1FOatLz3/a9
athJiN5Xxx7n3cL0N2u4ZnNqAWKlgUm9HCzES6aEES3Zg7SbcsF9TcX3O9/MYZTH
95YuEG6cp+1TyM67rCOWwxi24SBGZ5+HKw9XBJyygjVJnRQ0km8EIN14TloziBsW
WTiyS/rTAQJ1yHqPrI4bY/hOKcTY5sOpw//yteNlhCYWas3d+rH+b33qrN5Exg0t
iakG3MLy8CFfu08+XKoROWegqVmeXxRQZ0shMzlnUokpDn3n8uu9QHMKS9+BsIjX
kifiMAC+mrNQ6sz3MysM8sviwIMCrjhW+u4D8q0ccLtdP3anREzqVcKUI8Jof2Xl
cqhNSA+Y+O6PgN4i8cEH9RJ3YNn2VJFwLpasZAP0rFsYBoWLqMHnYmwRpZLovKja
q4/Lbqpiineqja/P7eU6Jl/dcHqEiB9is/S6CgDQqqxjVz6EWDUgv6I2Com2YxjM
kX+PECtMYx4zzU8Dp5b43md23Uw4t9lHvLNH7BpzMo49Gy7AC4uo6mfILplWUF9B
75gNQ1h/+OTuh48eF428pMoBZJOpE2NcE9vNJfdd2YTFtWeE2Oc/cUgUJdankNhi
64Rr/M8bUyO5/aaHZEY1mKWuL1FZITadkSoSi4ru/V+rNQFv/FaNQy1QghlWjB9K
BHevPmyG6DzNszNoyJaMWTTk64aTHY9r4aCJgK5yfglfWlxo2bPHQxQVVkgPVLz4
4XDnb94adv0jGfQucrAH22Uzy7MnOoBUK/K8+bu0uoXlezT5ZvYDMbRw+238+d96
zgkUoDh4rFN39S4v3StpK3zbG2ATANNL5UfonyyfeLDktyjhx56fdE9BVa1RKVqU
f0qbP+gRjggGznjJWS/iIy5S4ZrXnJ1r466yv53niLigIiNg/kFNOELsAVOlhCzg
cW1qrtZnse4btCI+zFbdr6apHJ6U+oHmDpWXDQ6OM997ZD2Em2CfD5N8H2cMtooG
/BVrEZAtfsYG1tj7t/2M3YEOAlyTaU6mWCnjzDiFoGU22uUJRB7TK5TbVuiEvDS8
LOA97pUV1C+PrM0UYQsYPKF1xqEVUBM40Q4s++/+J/XXQl9SFQfc31ql3/YCeQNI
STGj5JgN1DrxUUA0nmLKVt79qjIRpQcY9RwHYjXur5f/KeOMaLUr/VfJC6/W+mwx
viJwE0uSz3IlhgEfYvIOSndSNjuIfqBxt2FIYN/brLazLsD9pbAcNrfm274f47Oy
LWCKBxOzDH3WSws5386TpkjvDKW/VD5zWHB7XhjJHQqBkRp03XQdyJPaFd0TPaSU
3Bjsph5mcc+ae2Zvss9e+Fug6xtzVMXmo14/qYqhpgm8gDXiyYjxbpfBHDp12N4e
aceNRdICk7Njt2OwuC2R0nH5/2QJ3jjS8LTc+w8Nqrv7O0Zy4EISPH4klp5vK2Ox
Onth8nO/3PnnEDWRv2ri8OHFTR6jQCOSjdLyv0W/eDHzBAmAX1BAS5RZ2VUjrbKc
MwOk36TVefHah8IMoQMeXo8bCA1nDquON9YfUb1w05bRg/G5qUlLcilKnOa/eY7a
MlLbvs3ra49qKAIqp9+ND/VfpYO52Sexhvsre7fT8U2ehOm2IjUnK0/YdjPyoNj3
9DvPTQ2r/y4vFUeTEiPF7OmAHoh9sbqmRUAV8HY7ahOUDKIPjTVO5FLNMa8WgxwI
YZVIb9ZviBuXJYmaPHkPsnxqU1iYOBimEZ51miGz+QG8HZ8I+MGUE49RFL/lQIID
7a31fC2rEHhaGAziW4fLp+udPapP/DPa8Pfvj9CvSmLBnl/YXMUtNA45QQ6LL4OL
fy9Aa8jmflBct7NNDFdFCjguzGcBhDX9KkDbxe7rVrRrixydqsJpP5UsCSUFjnLS
4BN5rKoezAG/ZGwffa3CKblo7bisaTVppnq365LFLE21fe/xa986M9FdAtsp0U1P
7grGwzKv5EsFROkFGsybORwiUT3NIECdePyfzJ0BmgslqYEshI3AJA6BFJBiM33g
GuuS4Uk30owQoNQ5uI2HWoazZtUIBay4nA/HaNwjQdowC7uLVxGA6nFRYq6DdOf4
xk02hB9kGNniU7tZ9dPdIdhEW63wcRGPZwEVONFogXfNI3+mcpesTXHtzPHq5Xs/
aHuvkB0EtJCDH8xf9KdFlftGBvHqyPpmXkrjH3aAM73y8ABupF226Y5v2VIQfkrr
rpr5fOTcYVclam3+Xp1Zens8c8gv57VmJO9obIpV59D/CyCNmAiFIIoFjgNtaGKX
T6HzoV48tpASqQhyhaBdeyYjxSPx7VXKP2ck9QoQOyQEbWFcZ+e22/S0kX5evSS7
iLj3/xyNNhL9zONpNC7j+6WDPVoRNu153mdVZc7M3fYWhdPFOAH1KuNcxv0T8c8b
scd3nOeYrO1qXi+96if7+YWWtohhRuZ5NGwn4LYzQQ5XDzPW55rwGyy6eSa/7aSf
b6xL+pvHhFLMJuxdMTJStDckUdZnlFAKpcum8viyPM15Me9TIy5B3KxfzuGJwXAB
LUlX3wzEe652sw/d/zI5scG936eiddR9TrAj176Y2GQul1o9J2x7luGlIJ3IHFwB
AnYcY23E83V5k/Ed6T/ESkfVmzKYY6k64b0J9IAKDgxB+b+++UVvnP3MTei1ZiZG
eycL7BP7MOo+VNkGmqbjZnOHwX4pwqjIKesgDAc0SXJ+i+vBwh+BZ1knNDhD+yt9
L3OquIYU4fmKkZTuiHOjDllnk7e0T7K5KXf5ZUFbk2O+YfZ/sJ+EVRHVdzhGogAB
zTVnzO9j9VJjUASM4LHpW5rY1DXnJ9F/xoKsFvJ744GP5i24YVO3+/aGi6RvkzOv
4GnYbycX66ZDqWUl2W+/RAiPY3jT1P96hq+v4zjYPC0AIJsltMY5BVo9cr8dLz8Q
9ssOuY9EC2joeWebQbaJGY6imzU/0zn8/8wJubEkOO0vzw9cPBa18GFuvQKmr9sU
3X04CTG7TsyRCqwpIVUqjUwEwJPhB+rJxn1XIZ/rDhlckVtl+IAYQVDQjpqYuI4S
1/5rAQHWg3Lkq21c9XrRmOHTM8NXeCd3iKXl9dKMQBCN3Z2iopc8Me5O1IE1wlGn
dUM11lZhqivEQ326D+wRWA4PVH5+xF9MmIgONaKhzsF4NBamefs8kCO8HFmeUq7v
w8ioaKuhDN1Il84QF362lixhLA/U0CT6j7yVM8s1icuUpXBKUqJznQZP9tf9+e98
wg+23wBwEYFO90amOTiCw1qs0x7b6KcNmzZimG86lL8qgpX7QqwFpFv6UqJWYRSj
oH9W+gKzA3vvimA/ZKnpyEyZeW9nwblQ7D40bp5T25I6t/Xg8XPVCyKp6D8coaKe
93Iirvf+VETK4J0U3tSp1TfdOKL3BzjYs81ZpjmOv7tYEtM4kmwB4X3PEoH7XArl
O/ggy/mQ9fGULWSj4ToyI0bw5nr/I/P24MxdNFK+78FmpraqfELGuDceo2P0RlHA
PhqQ2wkCCzNj7GNpZD9MSIMN2/6FYvinf6K3pSi0uhcNd5C5f+UK3KcUwy3X9BTm
3ka+cNbH12AJmvFhNjGwxF1SnJ9A9dtCwJAC4sgGwn09faEpHN5wg4vDr/SFaNQk
fJFVxuE5CfJGSUuzFEVnB42qWeMDJzlo8Gsd2Islvq1ciVVGK/ZJrW4mC90NypYl
FOiuu0U9yez8UrWLfd4Cwj1LVvYdvGgdPKeFKVz9B3QO7/HoB5ZgAXVzwFivNrNx
myMqnEAmr61xDnBJr4Rxo63YwFmVBXoyAJEObOXcByPOBYmO0BFEuPlc1FFMT4Hq
Sc7Tzmkson6mNky4eOM6pzzBzxYSf5BCjZyyTIRXcywowZDV8ss5dm111Iyg1r75
NHYy7JwyDRkGMiFyKYU5JHTTKLsfuKOsvIx7gaFyXXfjjGsXZ35MNBMcKwagtMDD
hTmrlCWS2R0joQGtXZ0ls+O7HRy/qq4ms4N7pYnoTuJV2BX+/dViYDBJA9ugiw91
LHlvdMi70YSZyWfRYO3IZo7+XHDJy+aojrmR7Ou5oB839NNt7t0W5f4LkH4lLOlF
E+SmM/+5rkMvPAJzFx1AuU1wfQ0QF5q4o3PkdZzvkxeC8z2B00+MKFQ9iOmvyHxI
ObKgdzOa2lDr0B494r2vjcCS9h7gF5GBsUYDoLw01ZdZmULBsy8ImfNwBcUBSehU
EIvxytyvroc5WNe0D1BoXhRSIcnFk02IyZDkYOHTAIfv16WTdvfwZ0ZHhItCxa53
rXLhqlVdB602ccpPssbJEM0zSACtbdzt8Z1jlS8cO0kN/3uK9auBaMfM+ay2HW5R
7Sf8YSrTjKaCm5sok61QFxFo+4NC4OLpGrpOh6yMdzR6DVznEer3N9kzZAX5yIZv
VOwrnsGWLVG9QKuOalsDt0evVBlby2hs7psLHBQTzjWYviVgECbAAD6seV6VGETH
D4bvJPm/JgLrs4s45kDvlzNrCKd2lJ/ZNke0cdQNCqWloJf3wYLwi8b0qcDtu7jC
Gz0ImO98sSqJrqZ0TD8ZNDpqZaouOSeZrJVVW6plnGwQzBXE7+SRBqgvuEQwauEc
xgJZIfDU/8grGnJGC/f1KQOFeVPbQmE6CAPrhRjAGnIIK2VwA8aUb5bTEQ+qIrMZ
Gwfz5dhvv/1sjEi+DYTWXmlnmWuiHRa6E0KMMTGzVCNpnkyoFmV2KzS8kZ5xNVv6
oGF/eEgUFJ6jNM2cBgdZ7lHHRJcfL25la9jE9pvf1lUaDUKJJ9U6c8KgxYE0vTC9
HKFwQSi7xJRzbwOmqvJHM3ip8FPr3jVJ+irm/gAT1PM=
`pragma protect end_protected
