// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:33 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iVEIejW5755M5B3k13WUcBB2hUs4LuY7YM9pBMf6tD1q46qsN8RWx19JsIUd0KKD
Z/KOqX8DQktR+l+gBCbN8rVmHY8Sw3U5pNfsn6ak7bNnlTQU6naNJ7inWF3IaIV3
okObMftD9fAApvGft85p9UqH0G3osbJ5tsxVJ/4qE5M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5728)
HSJKCUb4wlEHKNRK7LYHW9RbmG7kiFoIQwyxP850IXWp5pG961IDVxDceCVLGSg9
4Qkkq0uKfSJfQtbLTIcT7eQ6ahIGbChIahWHlWypUhbvAuTvzJ1cjaV6a1PytbA9
6Wu84GJvHuMN6QU9/hDw3DDbTk4rYJKaynG8a9HQvT1D8y1m2phQA9i0pUQDmbuZ
pA5p9cYtRNCoh0tVsN56k66TQTFP+FCRLQthxPmnRxeP8ZPENMdpTv6z+SxH4Jxq
UjQiABJu0i8l2Bgql2gSx4ChztBZr2QyLH+pnIuSiwSmKZP77rTC4933AgJlAcAC
GHrq3XqncOWsFh/TRHowJK/O301S7NRjNm1/2aZ6mVvenvWOY6j93mvEQAuM0TrP
+fLLGG726x4YoDEPY73Lxw6Mfhh8GN4OLK98264J7qxsZgIkT1dMENQufAjNKdvm
za9eMLc1LxC/iRH4KFjtgPmf5KV6SEFgODtsEMg698sTcOwhpBqjfHIKZ7+hllvj
P8zPn7e5EWtYK5qKFMGcWXsCP60ODgYp6sw4rUy5zgE87OLgwt6p0HdA0KtvDUtH
r24btziOKhuc3rzNRuvYNHfdpr/MmOW/55CTBCH5SpbQe6DlirTomYc1SWC/Ekrs
1eLsxBzN6+tSQRiXORR/E6MIb+G7rJLIc5KuR9GUGUxrF9FhD3nAUJ/xCqff3ZPv
caDK6ZgJQ1RImTycvKR031BpuHtdIuZWSqDPtjNOnAzZDKMT+866flvdUK2TgAsP
FoxZL6dtIMXRmoWczroRNDQnRr8+mAGhUcWv5lZf8blmF6Dyfit5Kce+BrRuwq88
V/zTJ/TdtTHci7/hhrKMGYL5+pdpzFpzeg5EJqHxc0QMO+SMye5xEhFz8xRUkz+X
jrDK/uQZdvXsifCuuF/zPA3NsnD3u3zQIem4nvJXX1XFbBDL1iF2EngUQUruobYi
+r57eKgcSEXReZLP85zLZoGkUbzd5dPNO/lz/pvHEYu8i1kysVOeBXc6Z7aLrE7v
/IovlU6zHP96bnuf6Y85L2t+zGy0AEehN6x+npf4XJLCHsOn/C1Yva+SnCsRRsUv
XzwyGtb9LK6oeOpuFFSZTdCcLpcp/tf/UHFnjNbEvf52QUY/OosU4qaSAQx3rpxC
kmRoVnK/lK/oTezOi8n0UQzmPVhn6roZMhQR7W8PL2Pw0HvIGVnU08wd158E8QV5
ByR2sD9GZabBVQYniVxyfcRLnyYbtwJUCEIXoPerlsQVob/7qgeBOul9Y4B806Qf
xR4dfAHC5xfQkiVvg0+nF+78OLjM7o6VvzTyFdrZuvKf+r1Bqiu4C3lDon+mL5ch
dTUIGjBvLo4ffGP8TNemlGnZThyyVLZXYMGHNyO6wG1NQeYFRKPAPUovBmWJgFXb
DsFHv8aefYAk9csr86wYN6mHnFv5bifxOKdYLO+W5+N78EHXtAIi8v0/vZ5+78m4
npaomAl4MLLX8QcoHoaDff7UHfrqM9NDjjvmmmE+JPyDZnToT+HoMQe3SmjYmLcV
H8SiImALyrASKsrFIziL9fWYu5/a1zRTLSjdfYeWe9xuY/0/X6rgFrU9Owq7Mfxd
cV6n7/MIMLjgoXNRdcU9GNEStrwN1IdAVjoDZYkRbbBdf+BUbvCKXsQnVO+zstad
bxRQas8yAj1E0yCM5Cs7lo4XRzS5VCjHTQieVS/CmcQzIhlIQxU87FtRInPEBa+Y
ESLF9XWIowlOFgaXZZOtnxwg9mkEWUL1pOlni1YiVxqSBXGc5t0SyPyc1dpyv+cI
lFwg1HvrvjSu30F/wZyyT5owbQGYP4spAaN6lQS1G1fJ2V8ENKoJUF0tinmLZ2h8
5oFLM4HqnWgmc6u90SjlKwnu/nZK/XFx+OrgFRGaFp2ZtCWJImzMMaw5OyG3nOjX
Ow+N6TdprYN9S4ld2saGfOLKWLlZMSQYhDFhRs7lDJVxyNr4zkJfzCL0odMEFfOw
LpON0P+F3F//KDTUWg11W+UGLdYf0pDbzJwyeoOn/vwRwmVw4k3FwW9jHOrOgBU7
wCdltdHiYLGEEqllrnBWDUlb6T3mYiZkgihb2g2gYOjURb3VNsoyYtOaf3g5sSCu
A/5D3MxbmdsIHbu1MYO0R0rcGuE8c5Yj7KJomtvxpINN724KTn7xKNI3aMBfMlxU
6TOH3nTKBnwScbe8TJp/T8qTkpLSSE7VMStY3zpTa2NR6kpCK8sxetKGzVHa2C+s
sEU/5/kBUy/eHjccJkX9HDXAgj2EHKFRNKYjetE1JWtFSRpEodv1xE98k5znU9Fy
J+m++5TZ5j60xdFo9n7ZgpDzQ4cTAV5eNfSI9iDPcH3oETf0Vp9qd5/mpF68FGJT
3K2q2YwYtMRQWFWvq9Qj1oEuqXho1oSjrfqjp2VBef+xofBOzL85RICOtOt0GJwj
A/kqudY4CLcQl/guaqz5bn0Gqp3W23J7nDb2SBBdtasaYoMhVgokkOhr10ycnbhY
7A+rNPtOMFlFC59Ye9Zcx1ICxgyVE21ImjWPB7txqYZzviMgeY+B+Jmy+Pz06upK
vwddEVsd2Sejv8ScxjGcbYOnbGw/3Od0OubGG4ojQoIF5ZD78ZO8n4+O4AWPk6JT
r0PqS1PWLYBk1sRttaBq12W94R/8rHc8EnLVEU0NGjgj/7cHwslQ8d35rL/GakyX
Pn0Yh3a+29HLaiJqld6cQVt/4JPc0W4wr96TC51AmPd4rEFYULhqoEIQKTkFvBax
rJADaPkFJdOuTw6PxuSe0idH8CFdKsGGnTtR/8fOZ7Jw/pb41kDRR3/VuwCywHQv
u09i7caDFsvs8Q6DvdJMZqL0T2cSiMLAMlC+wyPq+FAZ99IzJG2tcgMdq0T3Q9Sl
ODo1VM34WRGw43iCtHNwU8zuvBSTXDnvxXvZBYuiQOSWgXcM+eiz3WoclrhXzTSP
wHah7LL6yOlFrCV5cc6K7xDdkJO9g0tSvSNymKWdupsnLH1FU28nOrFQV5Ac7X3B
TSZSfWGNyfOIS5LrHk6rd2/0Uudl3JuvtmJMr0isz6HQIkyJaGevAjr13LTj40MI
SzAq1+UUWxFmMjKNrPxwmqWXhr/PpFtjpmZeBnUz+LcGfjhhhsQ20Vi0S/XH7cuv
I3rnVf7eanw6+WLD+13CniZIOPx+Zaz79uPoHGyEhLHHzX5xwPkzP5QWQfKZtKeh
2Vgc/BdOfah4yNnLFqbQarrtVbGmZaTtwm+rqLp67z+sBH8Rz3esBSQNp7hGX5LD
K7Cw1p8Xym5cHcrsrFfWKGMxBCz6Ml9UKLnFSwqLtsaSEKKk8d5dbbx/ueyQCTnj
6ZYG1Vos7It9vzkiOFOWjiyXKj0CHl7iAml75dK/ZQ9Z7XwWGbXAnALKJHVyZuMm
X2niRC9ZpBB/Ton+l57/dLE0OmL3px7kiAfEdKlOyefmuQiDueVfPapbZIQSpDgn
uRgUzXa9XIZYRSD/fNFPtp9ZGk6CiQD48C6EYgYNq3yUEN8ZM+IV4EN6otsLCwRl
mP/9S9P3WmjpnOtBGWbLtqnW4XxRpttR0CntCvQ7TP52Z9nY6UWvK4QAWS374UMA
/bb24uHh67mmRS0CGPmc2rU/AuILEoW9i9SoTt2+whtur8BSck0qzNnbdZJd8pB3
YT5KsrrqcQMMxr2oR9aJj7aNGPyaRrST52aJup+xgnkW4lbfu3G4s33w4hDmjurg
qcB/xW8emm0hgifilRAIXrQpkAgsfDaHCBlwnZ6BMjf11tInBnOafJm9V4gc5aF+
5PMLfSHLzBbYOKjDZ7eAACjaPMLwYtAuoLU1E1IdJkai9y3aIz/UuC3X4frFSohY
3SZnXA0XmnbwkTD+FzkBUQHCDrWgQfbaXIGG8jF+xXzYF70w+AENZsKqHOr051Kd
/Ov5MOaB/bbHz86AhupryBKDvo+3RKm5EaDe4Kh0NZ9Ro/N9YdmUoZMzFKkIX5E0
PIEgN/g0lPGWiP5GMBRthXGgD+Gy2btUwmXp8aMZhnZoQYpZJv/Nef5A5GqOfQZs
af6cxRlOQECNzZu2PbfVZ2iwsbqD9d6+DtBWBaUb2EQeCEKxfV8+cuwxM8SCODFQ
uWPtZP/6TRH4vBKUJ1hvhgTpc3DsM/XRhpgiQFugdwlMsogzZ3fClYvd8TsWkSzO
rVVye7voKWtn2EIo9iSTTBaas0++RmeyudQtwKXpXJztDz/Bil4OfVWoszLS7tQq
byWwQZ3sVQG+sHyDYNNV+HFDjIQ2/8RjtPiajJR60QQe5f5B7/iHjTc9xob+sthR
FbZ1EgkbUwiRG6SuKlS531OIEibmtn0exTnsuNa+XnKAh989/bnD5wuU22E3lPDx
7V8bHxIHfLrUxbgMYypN0KSQkYYzILrMiNzncZ6rWWOgaAwVAKKdqUFg8BZPfkla
+BAtLAUIbt3crQuzaeJSSgyBZBNcPro8RnmvYm1ClGQproZE9AEhNHqbq7ePpy7T
x3uYh2HxOMVjJzQYYYhRGgJRQJCxleE89r6De+fdZhIT5j0ornLg52x4+u3Y0Vel
LEQVL/frKHcG7qgmsztsxO2K8piX7zWzjA4E3uSIpaTbQkDVdFx6/Rucc41lXbpP
2S+XYALdB09bvZALBYFQ9gul8JVm6TJeK92uQuXng3lrE0BkqRmgP6I5j0rwRaPj
8V/tA7QXt/khWdnIThKw8NxnERtusZYM60FC//bBuHnxFXSeFjfDJPMGdr7WVnat
Km4x2DR0u/UuQCxKc/smYXzBCYC3jKKaOfD9L2GnVUqWgfNrHsaN4QY2QenFLitX
2/Ptjpmmzl0/JVeS+A2DFDyumf+LmGwKsOKr9KEODy1b0TL3BwigmWmYEaLnxPB7
GziR8gfgUAvOooSZteg70dOf1BVSDBJSL2mpetuFiAhnBbbR/efWT/uNgrsunSDe
LJbLwL9hzLUx7IP6Ihg89QzT23xBeregVeU1+8bJIWDq2pbEgp3fej/H38VWpHdZ
7l6r55YRf6hHGsEuUPLwcXiwbu2XdI4DUefeDrOyV/W1qmmA4oySurIxB1rjwBFp
0U/r9/1ASCTRebXb3jhwsmENFFxSapJr8LKbJPRbYLfJ8aU0VTPCaAHi+cpsuLXb
et9WzrOPxUr9alHehdNMTpoQSsuMhXYSReEtDLO4nG3aFq5qHVBovuFbncTs5dsM
4VDNh9q084MfFB0t0ZobRpqS78t3THu/r41C/EjiwWTNtGzEDwhj+BLAUKOEQcYm
HXay48Qpl3JrQye1N12Etd2p0ClyeM8NJkYf8oBMsn5SYyhqqNdtx6HFsIMs8jfb
FauzM/BGLN6Yih9f8dC0RtW0O9t7dGhhFdCnaf6jCgDO89+zXWwT+exewOp96/6n
re/fSCvdK68C7AWXucbsiXeyr9FlVMqPFIGDInxSBD47JlIjHzI4+vwchuHtH+eE
oK0ZAj75sbw10GFXnxsB+Tj9itjZ4s6DNf+0N7UJwOuRm5eT4laO3hBRVHugWxWj
CKA/B0cpK4MS6gmQJV7OQukmMLmfzOph5DfnQz5oeCjVwoam8Y1a1G6BP9755kl2
PH/X3TrJAWV1OZZyPgiaW73ODj95edY399bpr3r1FE/VDB1/On0ohuGAG7msd6df
4OYQi4bdl1ibSu8d9hMaC+L4ZejiP0hciKjGiC0KB2IEp91mIBdE2m2GbIgZn/Y1
JMHNQ0TGE7GTHdToK5WB8FPC24GtlrNX8+Du1tA2tuB8An8n2h4P1MaY0Jnxxfwf
DhUDsJb7lIR7OEKmudE5yFBYpmfzTwfdQ+kFrcNnRDBOCTPWVDDTkOfpIelfr+Hk
enzIJi0xo3z1Wb6M38hZV2iK9pisy742c01MmOHaHfkow95/m9/pBSV+1d8sBosQ
NCk8Rrpdsz1nYaXNld2lE5/eV7YLvj0kHRzZKUBpKKyJbQpsslg595S5eUhTTN1X
nvabgNgbzahKXdjVxOs2WG6nE1fUn7yef3UHpfSn9SdyuBwjDhU8F2V0O3QFy39E
k69/xyAo0Rbt+de87jmiL4rVUF4spyPHXv9ycBE+ALvcGU2O1CwuuxcvPjWCzZMF
FG7gsDUyF9pewCjpy9cJ97vw+G9nuHTyFgsAuR5oO9puqQv3kK9/fo46e0Nx55yD
uylF4dpGOe/TGyQlkQTChbORID/R9QSZnUJ28qym4Wv0JT9mflJQcGx3vFNTUrHZ
Ax+ys/88rA67dnbTyw5xnjmYDWpvDTdA5Do4pPj2SwV9th+hfp2ziyj2GbuIQHfY
fWU8ChrCjlndaCoIhGqzh4i0XulhTdi/LkygIHFEIZJkfBaMpK0krKuaFzQWRqM3
Tj3lyZ3Lm3+aApwM9CDWN2lU3jyRMxD8jxjmSZMH5cuVa3EykHmqw2A/T+qwu8oT
zoOcGcsZPoo15ikX6ja9RzwDfcLWe1pP+xTh1PY1ZuQJoJkf79nARkynCCGLqzSx
SUqGzo61Y+7xbI5Q5B/dtYEGIuYs/kmwRXlTSAqMUPhjIOTK6srr8WAAIbeANFN2
O+R7dS6o4PTNRgNGXBqeZI06BjoI7c4Pt5pKXb9Ttw2kUxocALLgC8LZDoTMW96N
BdnarNp5Knss1XUp5p2GVoEApET4o0s/VP38tIUoI53K26XGO4PksNFt0GHlSxb2
1MO8G5p9wAeLdFPJokWlKnoHOJbiP5RnWMrX4zanJxhKMkfG2EDNN1JJxV9FXGSj
loZMu6sbShRiVpgw9f/WJHHShJUKyOGxalCedSKjY1p1/RrnMs/3VspULdr1aPlw
QkFksZsK0Te7zzT7chozOmVqrspV+D2QqJOxPSREOZSr80YS4SESJ32hy9ECYWCJ
umg0yY+7zRh+F8virDVpTAdD5DkJvyy8XPJo/1OcmXzRnCwxUAlPNegeyoIveTx9
bsBOnKZ7l5+cLFTQB1g45FfJDn1CIMQFIpeGHTH632Ib6gsbllvGy3ImqNViAis0
EyKPih9NixKFGj11u4O8j/0jbT8Hg0vSZVlIVXOOt30V3BTdn705fNcxwISicHoT
KXUQo75HfnxxjaIlczJwCAWu369CSoJQUzY1ol4MAhDIrVHqLLcn+MCgV8erezWa
HjtSJjqj0LSiTPDkouDW+TfHcOAGxxH+NtOp45WNdaJvMwcIIUW3pVXHaeJdI6EE
EmfqIbzvGWZ+RNo0+tW/k+7d0/ihRc5TDGOBdYbhVhOeoCEJQ/vaRLu5IiUuRguQ
WYlN1ve5ny4q8f14AgJoOEsVQg2cryl7cZ7zvdkBIBm13DHzyDJAdUrjDXV3DURK
x47onkN7eOsRJ3XKIMZBrTn9Uu8WdI/d9BiDXzD17blvulrv/mC67H6p7HS00QvL
H7aMc3y/tpdYNm1yCWwyTyeISfu8akipCWADCZI6VJdRgAOiYbMaMCm9jWUdYNI8
LZF3EojSyA3rcFe1glVFvCJyITUfFgVuHGo7YFT8ceoXg9I4AhhK1UJaWFCSvjyP
AVcc2ACdI1FuGuydFEx0YTJ7uLiEsXVQh1bs3ANHdffYpRuzbwtvgCoyRuIBgXVf
NwZxEhVW7XaIYSRiXqqdRlAyg8lGjsg7bZjA9CA/eH40lHWdQfpoVmuUrZuQA6aX
cvX41D7oTdtIW6PoXoLctA==
`pragma protect end_protected
