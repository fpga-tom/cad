// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sOqO0cN0s0KZnQ5hmiEZHl1ehLUrEFv+ng2FvzNwOisLBllZMUG1MR4UCgF4v6LZ
zPGyiLfHxSlRMQtl8YF4E1NkengbolE3443YVVpnGTvj9Mi3P0WmYZnj4L0SOgek
jT8N2enuOfQreHbk5Q5+0609bQnAAlNMIYJLWNjm/o4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12016)
MEvbEGgFRdRs3fikUDGzFW6RAA95dbBeMs/smLJ9qat4vVJ/GiktJ77D2+Y5Y0ts
jVhkOFo5tcFFFtt+DiUUPBqmckiq2VIfTVYYCMHpwg8gGK/05ISc6+n20mH+2W8H
L7cLEmM33rxztP48I8rja9uM0wJogumy18zQDI5DEsxJ6wT+SQRDrGx5a6PCQH16
EpZW9JqT+0od9wC47Bx6U36BBTDqYzLG0jI0GyTCmSPWIwumUwD4ZhrTgzaPOpTU
7PUsW2JVUrP3BBTs0knVMtO2yn2x1sIhlwq8Zlrd4CKnn4MLHjQhs/SBk1uByzJ+
bpZl49RAvd5JexvuSsd/GYlYKCbNz4sBq/jefU4Xnf1j1Witd+mCbDHcyji/N4n3
yINwcY7KZVXtEPwj4G1tzDjn/15yGnrt6yPi3UYjBNg2jIBC7IDpYpBftWYhe46t
RHc1urIoVWzVz1JneYq1XUDW76aFbePCqb7aXpEVbDSAM5VLkxKy5R6JxYDJa+AJ
gA/in4RJg4OiQhGd7L8Jr39QYiSCXD+0neEdEe/mm3jCJA/0BrgrVdJqDV5S5Fs8
muhhSWyNjmz9n5h1yFq0b4QnS60v3jDbtzIQEiyRXTlL1E5rrdQ/Y2g7hzpBMw+N
bZBakqVLShCcCbPS0m1ecHzeizuai4c8BNxQ619lzVRcmWiQ++pi12dXJKxYpGhp
KheQwXYjmt/SoMZY+4cpUQmNjfwe5JboIpnss9gnHjXg9l02Nlp7sOyHd4gIxNbw
nAWN+cFl/LfUrh8RZiVfitGAXWZWEx40bpGzQJsTlQMbR1f9OJFlpodvmsf3mK7y
wNWMVn0orJtAaWcVq1SN6Szq+SI1roFRt+8oIUh7mrzFJzMankrBeI+O1lIfrHfd
CIe1wHRVyE3LYv8DYMMU6x3ShGTVJyfhlxcy6VpaDctV7WCjU3NYw9AfaIuMwjnp
GQ1oAzl9H8Atv6YI9ftXO51sBTMfuSQHeJy2sqVBRkfJ4r8K7568GdBKZezwF78V
lLWpDNldMm7WcMhBN4zar0b98apiUkqibV2k3CR+eoUx6W5hgsaf2kzsGENvtO0e
5c9nhiS80+QBSlksMrjQU6qWR8FhwEOtWAuMDeuEe2eUXoRQArui6Vz4AWfwi116
1F3NNQYT+6yuU+GICFg2Y8nIYY2pZq04iDtR4CFN+7m+xaKAkDbFbtlJEjvVbaGd
JF+ze1k0710PzH8eoJ3eYrpz9Idk1YAqCmc9/exGNN2vFJmbFw0TEpGGMD6V/TRV
ZFm9CJw8lvPn5KvCMJ04cXG25EA7d6e57Rjf0DpY3ojwpr6/AUdWKRmTumZZHToT
mLUdr/gEg0w7nZvflGFBInwZ8TMmsEzXAqwh0GbKZ/swTbnFtQ24cGMUbdOy6geY
svvRf7X5a3tnspjMdhfYRBic9IYNP52rm1ZHZBEfnKbEYvdtA6FuA5vzFlIvPuoM
S7XqUKx13z3EtfQe037eSU/qIQruneWAjZ7HUUWI2+3z0k8VybYbREmfNYN6Ftal
PKx5Mu6zj9VBK3v7ayIQeRgqlL1lO9s4mKubS5YeemJV7829tyzwj0+9/sq7Fhrn
folCVkvJVkDcX3Tb3JHZ2RfhnUCTNmDYO8Jhji7WRKpsrVqLskNtKf+V6+etC3km
uCt9V6PbLIG+kKl1DFBp6reW9LTbY0U5OT2+VuoDd2kFQqVZA2awDlHLJvsKAVzU
awtBd7bswNgtqflMcUMF3dmEfDsLNxr3ip+aAri3zwvVRuAfSRNlfeJGR0rrwLdE
mH2ui+blZv4U606Y73iVPWyTwZiq3UD00Ms2UUBO4bCyixPRa5XZmvo5TKQdfZMe
XJ/ltbFIR39VezcwoLfY5EstboPrnpt1sOZEP2NYuknWzgbWxpPovBgDx/gBfDAd
zHgNMPW1SjWDLU5lKPzutipzE/3ARh5m+EGnLAav652wHuQckSzhGsHTDqXm1akc
jSpkRVUs8/toaJDhr1LEtQltIbwFZ56OBbIstyzUN1XFn2jhDXc7v2iOshA4VUVb
q+Xy9qZzzDXRBafOQNNJt+JThrnUc1w/tdDNEhA0Q2uVUpTI83ZHpjL7gW2ow+SR
vfR6evHwSQ7mPJOI3uWmkZ8iiUd6BYbKeec1hKRRTPMMUdB/ODt3BD/3QMJy4cFz
FTwkP3DT2EwxAstASJxvEE9auKf64Hs5wYk/IQ14sJ12kpm1ghSuAjR3gMonqXdj
kIkUpk88LS+xKzNOdlJy8T4YHfFcVQhBTsx5Tp8/2rnVZAyGeY4HM+vFCZIPLPG0
tqNa0fQqoKmYa0YjCPkRK7Ziop3Kba1SlyHHaBBV4jqJgyfuNPTI4Y/DGjqHAH42
EiWVpT0kOjCATqbSGKVCDj8tUwzbfpPBWJn3BTeOBkrIbSkUfzwvcTD6akOrxs+z
FJQ9EQcoVPNnZ+/gd//35MVax0EEKurCJmU2VLZawg8aFnN7WkJj+94GXeJQEPIs
tEOW4lvuc4pO36qb/A0ruPvXQ2udvkFEx3Y0rW/d4U0WYMhIwLoBuBaxp6o7uvio
wvvTb2Ps35HiC85VkVqFtZs/WC9gGUzarKKr61FKihZbMKwh0Yhsaufp5X9zNQOh
FZsrdox0ibdU2HBn+Qr3YRc0yxe6YqzZx49zk4j/bUgZlrPs2YP8EHYZ8Zy66u0Z
Agp89kNdouj5Sk72lRTsArX1A6FTEdQ1C/Z2aSlSInkivG0L0fAI5jpo7X1indgC
mLIIkUpIJweWau+anTXtsDKQJ2I3t1wmFgqPR1cPAZ5+Dzr+eqiLT2xZ/gwo4IyR
azXFJVW0fd+AY+1SR8GAijTSKeYb0jyP/WlirbgW1ljtoohURj6Zb+SZuQXLaidL
06yJKIxC/ASU9rrNFN57JST/GmAHzIlMQwgY7heabQKuVCAMYeZxoTkNBWBtbkXI
5vD7EQYVXQ5xVUbz4mn/Sl0mG/GWAYkf3Np7tPT4QAIA6ywddR1F4tzpulwmvszt
mxmpxl0vd1tj5SORqigG0zFjKkjSCjx2QH4tgPRlkcJ/9YXvyTWNOmumqzY0u6nx
mzOny1dc+FLEfWvGm279h1z2LD09+jBHWTprDW5+qc4WLoFoxu1cv6MsZEXXyHct
HWLPcmOvPczwk05UpJMwlFvh0u+MFcMOAqZqt9cT399UViGKPjDi/8Z/eq8T4CZq
CTJnK9iCk8n3hlPRgBBbBgvI026lbMYvliYhpPaA4GmI/lJMe7jO2tnE9d6o5ZWa
xpyPJfvt1qEvfRJDrAHCtEaa+s0S3H8eGPfb1dmVqaXKxCYwBdMt8R5AjekgoKwn
SUloRRgj6SYCfrdYf9lb7bmtRMOXkGcVZ6sglrxwtvsjWK17QY91JQbQ57m/5y81
3Bq5tKzZ5Q9RqNMaf1oWgY3cfGvOG/bD5rYTxmiBrzeFjd5auUstDyWFF6Rb0Jsf
YngPMbPxohPUQy+NvrHNQ+1JsxzAMm/4HNwcfn2euDehAYzMfG+8BhKkXIJBxDwf
zE3LfcRtT/qSmlyEwKMTOh+jWQe55URTKdWuXatMpXz/8z/1nLytBaNS+iEQaI9F
KATmBc2aQJ3iwuV40+Ph5fd8L8Q5yGEKPqL1RnsTt131K4Ws9xgbZpGWaZFxsRG7
/obRHM5+SjJB+AoPj6FPuaEvzc4UInJgXSQs6fqoh7MXw9yK/yywlcgrZ/rMBtUy
K0ajxg+Rr4zWO3cYlvhxJqvaTLsj9nJ1kFyl6iPtp1PN7tkEwBBJGnc4h7kKW9FF
+i7X3qNE9DqK3VgyCJB2aYy+9NWXS1oADSc0uJxv/oMwFJUtaFs4VBqMZ4XglRNi
d2fznpu85nao2gRIigremHCem8O91sS7A0deoM823aOsZ1nNcmks0upDJBjnWuet
ZtxDP2VelEd8krO6vabe9R6+wepk2zyCJGQjmJPjhP22cgbzuKTkoHPaGRz1ad7b
CyNDqkbCLo2GkVyfO37meO2mosHGPTwYvaaLEmonmIwlAGI+kWYfnvjAr70hD/6D
eOIAMaSzc8jJxbNw4RXYQk/Y17F456qw3DNzoBaGbyA9qZ+82ibSdq3r12SY89pK
WST09xYKQs6JcWngAueFlrta9Pf3JmJLOycAXAZf6qX6DFIxADD7tclaad/+gOul
oOnn2jPXxXcawhgwOHaWD2b1ocfXlcN11UYv5NqefFXK/GoFwz7qjpGFFOQW0Vb+
rpGnEgBNKerPiAXmxltZl7z6vDaRMhfANBPvvXRRg7H9xAmwX8Ln4+Q9uu8sGfGA
/tQQKxtIIcHZyh3TpqtTwncg35cfSZlgnpPAvHZPQ8KDeWbMOSizdBMKNJ/24bE2
eBKhJNfMAF9D9VF4iBY83nxUO97cySaM+GEXAtVTKwet2/KVQpH02S8NFI23gFFK
QS8E3BgkEDNU0HjzwYG2DG6YHgEYfVIFGZyqqB6trJ/VvKwp+NevjLi0HA1YnJzK
2pi9M1W/pSnC2DaT0Ps7EBXRJdHBCyQTW/jSnPjWH2BA8dcRLZKiUW5ulcpo/xeU
2WVXVXxgNzm9c02ymHTYsXHqWXnU6vRzBduJbAG85kiIyMcSYA/D/R0WdUd3xmt8
7kGMUVGS1RiDpqh7p+pbgt61/uw1e5uYaTBinmbVfeSSLhNJ5T8/JvSeQncWPd4q
CL1VxyEVu9NljfdSw/2LDRMmgGbmgvpd6k5SJNRxd32tDihq2U9ChlNuycxXGGZs
iFJp48U2kkGYbVBZkPVzqik132tEqBz8yr7RzmbdCIcsbnKRMNe0U9FJOEcos6/O
e39ch9LfYTnf8OUlVQDXXb2rdBMwui9ykaQuq6AhvEygkMsn+FBU+ws18Wr04DsD
1ER1wmJqXwgE0jw0c3SIeDagSPV9tEh6icgIFrAFQMexLMr6L+XAsfu2P+F47/Ek
O/nBBCxUQY9DxDCrg7mmBJjlRgxmRjaGHyqHhpeuDZ8stVwhPK44sNhY8S21sexX
56Tm6foe0zfrBkPlj2tfmlLERhcTW9H6p/938XmDtz+ojzuZM0jKSzo2bHrIzSe2
tTMDoMbKGucg60OE3Z7ALYgwzaDif5Hc8pkURfA/zMfh6sDm4/pjTpUlpFFmtZEz
vZBKxBU0cZ3qBYPBP3IUOdCBFE2q+DtjHOghCkA6xLXMdfRL4cA26NDz67vrD456
q03QxTmKNpgwte9iLj3nQkvRETOFaMb9rmpignLr9Frc4nQC6rVYU8hk2utA/e8b
5+fAC7hh08yuq/SDAeu2TBlVXpSbbkoH6AVGjt8iPYjdaEciH7PYUlPRsDJYVMRv
KkF+NquG2ExGUOs34J4VMNo1SOkOkSl0RjV1VmtSmqupLAT+koBiHFDXR0iD9Z2J
rrmI3+UujKN/y7Q0xIthEzLvejmXk/4b66fu0Fh7YP4fUF4otWyvfF0DXUGic3I8
bNJG0BdtisbuchBhksl1TnzzHYwu05A7861kn4+qT4GIc4mcPaNZseUtxrkiYyQE
csrvV7oesQSUIUhZDvpIh0/Biq4VUuxtH1iQsfajs6WSMtlK4jDxB9RhUmqmQ3wJ
2JZ/h6Nl53yZpzvmXJZj+C4afEv5aMOY+EjEokFua1BCprgoCn0Ol4ZvFOliYD+Z
WYIsQR/JQUbdCoqyeqv/4Ybbt6t0pmQamhn+k4hbsUlAw7F+SpAVE0K/7XbKdTzQ
SVKEWZx4LfFlebZud0W2ulYgFbpvwkQCpd4zKXtCCzWkxrChh50QJkkAUDStFJ8e
YQPbeVsJSG+bbQWtlu+tvK6/tH8khj06oW7t031RYgOHk7fa7QfK24KmKRMq+Hi6
xsveWWmpHxEEOOw+lywoVjFe2YvVqr7kCqPcGIyvGGkOSQ9SRqxl5+6ZxYed8lGy
Wkeo2yGEuAe+gfce9l8uJ4Tc9QrFcUgVRZ1x9yt+Ffxa3Aph9nYe3Uayym2fXkVv
4X1YWFysOQ88oiXCdoUMBoXw7CHHYwPVq8C1uYKqhiD1CGK8eiLfLY31TlkOo0SZ
yYxw1vImEkqVfSa5lxL3Iih5wpbTKNAmRmazTEHd3azo+hn7WMlfFIG56rOXY/j1
4tGXRBDRCPwHXcOFkHMHusJFgQCl0ntw1s4TyQD3NePWYNFHZsPLQAWh0Uqm6jDF
uLzRyiWaPiAtfQTe9HVtaAuo/c8hnceGG1PzFSFvtAopNrQvDN3LIT+vgApzBjnt
fgYw6D4C63bOIshlZJjKtwUFz67CzWHDTaSjHlibctNjhPmoMbDPLyR5F8ovtrcl
HY/2Drb4gDMGzOzEFoXxP5DHqAXWInSYDR4aM1tlpTN0W6tSEGvGlZASYykqu/kb
BYgXgC8pxP1ehvZpnR1Vtin/n+hlRIXY1T1YtE3CyLtf6v7/M8A3lBSWWhn0DJar
40Lhy9vW6DZgoNIEo9ZqqoAM2wLQih1c1Qu/N8yiBFpUCBXgkzNocQI6yqTQEZzo
gBEEwjDEddNMeyeWEkKC5HSqKZNZqbB6KN4W8240QERvtrz2yATeJmBAL7tc2bwV
KU0IqrYGqqNWBftakfp1vsPRuP5uEflqjyCwo/fXKh8B0GtA6mfE0kseeYXKCTBw
kkVzc5mmeA2icWzoujnb9sO/SaTVtmxZyxZLqFxA8ofmtBDuVoCcIFsAdMbguLNO
+FfgYrKll3L2Ub7tJOOmNovOSeTTJgT8V24SHVrdqu0NzwzrYYxnGRHG0Tfl7IHW
UzNwUU2KzcRWtNPI+wzSweFoeT2vHSIUQm8PGXDWFj+/xsBQfv52m5WPXn9ylx1V
Ah5AZfJQgEJqhpmrxG6L5WOmxj2tvqD8KwfMqxkyj0NM5hgF8XTfb+yr47kJ6Bdg
yBt5lwJuqTJEoGAYrwzD5qgiC8AHyIQEhM6uE/xgAxP7tLKLWPpirFKiShgG+KrM
fczudzVWfbz7UygFXRaCWahDZG4LIaBfHVgsNwS9zQG2PbeNi4Da+e1pzYyB90xd
FLBhuek/YEE2SbBwI2v/UGJEsPx+jJ/3Fl3w8nz5KnefxoPYuaSav7Ww7ggdDhKH
WbEvUMOaTgFg5v4LFK2eGG+bZ5mRN+Ty48zR/uKfJXHlPph2bsCUxuPsPuqV8tTo
zpSbtEHpCbpQSHIroF4yeeSyhGE23tlhXXJ2TEyOvDc9tqNBC2MC6Rmjds457pxK
fOZ+QxBqFWNK90LGZ+wcFQLH0R93hYKQIFrk4H56qxrPAtF9OE16+mHnVy+GEPPx
U43sBaOOuyAalSbfXlNjLOWOR7vgTv3MiwzQoWmRHY3+CTqM2r1JkbFpYGXMns4n
0mB5V03sLaY6GjeUDw+JyIQW0nfk2v5Hlf3DUM/hPhfO7mh/S1eDkiuRMeuPK8SU
Zxfqa1THIsBF8k5RNBVzrPVmDDChP9cvRvuWEG7pvIP4O+6AvJ9ZQ/HfsNGdJaYi
Du1yUAPUhMeamwcjVZU+RHNIGgxydsOzZ6p6ZnzU0DU5AUUDQPacpBOzuorccFB3
rOfeVOjQppgyIhwJvaaYS4tB2Zt4rEdqzB6fHiDLt2ItH0fIpG+oGD5330knhLDB
zZfyoleHPGz+H08M0tZsPVjZYGzlnVONxqw80hTk90LGF/nwi3y5ByFISJk4uedL
VGc23FN1Ro9qFwsC8b3Yt/j2c2x3G4fXXh+xSZxsK6m7INks7/6dpjpyEiXZZWGB
p1KSq7UNRtF9vAksqGfmOFVDx2mqJRnf4k4JhGNXZgo/u9TQ130+7kM3PDGZkB2i
EzjtH4yk49T7EqxRMxXoHcdxgUWwsu0g+srtu6jIdvUowV+c+PNIZuCHhg0vYMif
UQs52H6alf3y4fiTQpzSKUuOqyhimBFCMlnbNCCJFKI1a20xTVeBGfi2ovtSLsLg
HxzpKHm8GuMcUqTdHeAVCy4kwln1Sbp6Nn/SpFiavDndrHdxKN++NZpB4aUpLiBN
uBrFmHEUAV6JfgxNPTgZ0GoussOY6ZA2Hwv4WHrD+CEO9y4F2bJU3nvQJf/I74sR
go9JqvbTTHqqVwIRBiLHOIRfmS1bkqWMcuKrhueSWpGCvfiJz+ZKBoOEwgBBwz3r
jQzXoZoFRwtrAaO+kiy2ghDdggRWIRlVqNIjx3/74/jVVHyTjf0kjFyGANZ70ask
99Ju4GoKXTsrkevcy9OQuTxqKETYfVUY66utRlN2TkOARUsBNFrAvWVOjL+/uQ4A
aPZAJxrpasGYw8Pi8hj0V4xS0bS/Znjk+TFEmOzUcX2PciTOkDCXXuKPjpMsEPHc
n1+AtbHM7YHgcCpUpiiWuvRD6wNG9sF0A8/hEgKhFvHensvSwT71xvCCQnNaQeWX
QyFUDz3IVwe867n16nO1Q3xpqY/RnDFEJeOEfIX1ev0L2xUVr2iKpIGEczVQKi5N
QrG5sQm7aKkRzxircWSa+ArHcKbkhlyC6//D9h1WSLHPqRUNTfJObcUFPheG2dwy
dGaJaHVbiK5BCYAd7sIPJEl1v3VpfRrdWc6bIll+U22Fv712weDLUj0o1Ls3JslW
Op+Hw6SQ0zFtbs9K96wawflr4R20Rl18pZpJwcEg+Ra5cd3oHmvlH7RIUyakBC+W
JBQNkNnPcYk03vFztJdyqskJwAcTLzuBpJUJf+HmV/HSjW8lLVzfyX3EkhSAT7Ow
YqBIc0Lo51xTEGyNJX+Yn7l/9dAd/rGfah1hVaSSpqkGJzbOavA6+I9Mr11EmjRG
dL/MIM2rSmHikWW1LmAoGcSDv8HmOOYHUtRsyylbkn+EX5n54p8X1b6hML9vFGup
h30ackauv8qhSeIEcH4griB9Exztf/paLy9zMseBnfyaYzeSUpjivdXNtK2Hz4Pw
bCKbrzcJq0bbbn38OeC1vdFufpB/3ZVNN+L+2R8VcZE02mBR49uhBzGZpJcvWxXp
NF+RyTDj6B2GnnFG5SEhyxd+fOHaq+y6dSpGRe7NSOBS4cjIE/HnHyPtrGi46q5V
QUJWnTwQJrFkxwM4tJhOT0/0A5d4SFda+vKh6lxERueub0f6p60oz6V/kw2vv4PU
aoRc8QO4cq3oX/aXuHi4NLonXtJt1Idfh8h1sBHLWS+npV+4jVITLbFXUNwH6aGi
h1xkdhmPhDsKYn3cKs4s+3LHDALHwJfpdloLiM41o+1Kf+p7uZgdzPuQOSwmhYbx
PU0HB71W3Zg54RsNEXrKom47XGOEU+RDeosUsjqTqTCWGK8mCCSlperp2KYBpU/5
SFDEiJEshxIHGyR5dPHTs+EnogLWhSs6iQChx3K6Zr36ejZ3aqLl6X+Ij8N/8SWJ
o7XFztLw/nq9rLSm0JbtbBUdrDsvWdd88GKULYTeqHURRZhT3PFAnSWDwd8u5vh8
8kzHdvR2qrbm5oyxme4V3J9CgFrerewRNIlfopNwBxE/r249AoaGpdxp4EttTni1
DJ/0/pmQRpdIg0KHrVh3kcttfFUie/jS6e+3/DX0VFl6qopTSQaVWIRkrN8GOGE1
rlOIP5xy8yarIsMsoD3y+0CZTEd1JEtmqojeoY7SKaC3pIiKOjP/JgmE1ZcB+tcc
dN0zTp6aU5zNw2aRuCqq72z+AmBMwQdM+E5V7O0+s8KTPZAnw6FgpzAe0Nvkr80I
HvNAX3R/W6uYs3lw79YyD1tUxsuf8VZLYxZccqT5HO5JjzefyTpqZqmarRIwjpuV
4onmo0Kund4id68Ubfi97nfeeEGGcN4AgztNeHzWJUVeP27t1gAXaOmX8LWWnwk0
uQd2vCfzAX4qHxEcm9juGh0J0VuMQOyB80XElED+tNJz1VW4wg1i4MM5PJDguoj6
cU26naz2yRuct2mp8pmxN+4H8vxM9iZOqdRJiPXhYDtBpVxI73PIntvWhuUSsijr
neX2uCUVWTNuLYa6qT899OOjAcCwWbjH2zhCajvMUMoib/SN0n3MV4RD3prBBpDC
SKHD7VOTXzhiupH2WwsS4QLjLYChjyhxAGJyrJaFIg2kDKZCWnd7AquAbFNcnISY
UPI9KVwjc54R0q8/uzg7Po9pWj0I+bTfbIMqgrFTqqBVCyYyfuX2RgNGWCB4EF6R
PrlowzfSDGuSwdBfhXQhlPdlsv+XJ9Ii5Md54u6lbzJ13kHN8joDRssXrO5Yhxqm
bMfdQxsrwiDBkfOhh6YXzsMiPFTo3LnfTtAyUO21yrLatP4KT29CUf5ol7RhXv2f
wnMQ8x8a0Yl2Dp86deUJz5Lvm/VF8QFBRT2phcUX4yG/AEB17jjv/9I2/7gwxiLR
wM56IaNfgQHk1jl22On79sdpQetaC4HwgFfjApHtpusYI5fQtzhZw6O+PmMHF/I+
nj7i+R2vnb/5UTU2F8o/UlMfU6tE4A3C4NkYwBdzLlRnehHXaePCp0TRrucsuinr
2+18GsgRTDmwbaF67wLPNMiDU3dmB6LT8DMY6OCk80aiYEbIu1LhLsHDTTpQ6GGp
qJ8e79H5YOzUJRf7xFI/UYtZkVVGGopE9PSs73HZKhR4IaQtHMZ+DZJtRQJcxbYH
hV9PNuclCLEO8tL7hB7DeJXErD71BP5P49Icy/g3L4+IR248EKE3XwdKQcAjfB8A
4OhMO5SZ4pCmpx1mUhlQ9ywvFN32Zd96C/Z4y4Pfy9cfGqKLle/b1p0QleWamWX4
vIBbknjb6n5xEpxeBiBdKbEEworbPtRiRLcyW+MrqhTlhrwcHoNaHnTGLD/bO+jQ
0qHTKiXY0rcCOMc5IB4buAJ9k7RKt/ix1inOipR7ZyFWdFPJhY5txUnlUfTSAtGH
N0q9c+ZyVf8s+RTdlq1Hx2VWsL2E3DftOAEQlxJzrB/dNohjFXpxGbwHK11x6ec5
cLpKzWi2LF5uDcYccs8oTNNqPuMcS1Zlv3IzxkDLGK/QBttBiQEuB+TfSfCQXi7J
+AVOF8pGGhySDfjEBPnkXzyM7YvrOLSU7NHT6uMtycW60lEHoYCkwMki3N2rTuHq
6HregktLt/5qN12eeMTIkdreJk/NmoUm3En6GJr4qnbwNQL1V36RYHFEqnRDxkfu
1GvRwu5aMCyX+jtgHn5hgbtoywqLXQHAa/+6V2RMJIqNdqVLMjMfab9jHFxgyyNZ
efztah+9v/xf4EyjP3Mkk66fimgOygF0+4pqzoSTrZYnRysf68a7kCDMDH98mEPp
k5Wvm0jBNBJNh7OcCxtV2YgRXWwsgwKtr82CvXmOXALUfgLbLqJwsSA86/FR1qUM
1VCw33x2hoKBYEpSqBZjjvp6JHK19BeIv3XCb97H9p7DizXsxOrRVPXUXon9pa15
z9r5qOzXrUD9SrfGMY/0ghK6zZFvqbQz/17b78iVEwk3aIeyGgPhMBJMYYix/42m
0cyae3EHicb8IUKwdjZnkBsz7YicXX4g3Hh3HuqCMrV373p+26MlTr4Eh5sbrKF4
6k7iwy8dQohIodMY02XkaWYY3/MYahzhHF6+ZQJKtg3hL13etfi35LkAVS3C76Jt
TLvBH9xaw1n+q2prQi/VvNEL2PuRV2xHzucA7Iy3TV1gLuUUciwRu0bOm8JAQieR
4bwiv4zrTEVKSctSJABJD1a62UHZSRlHTBEJLKaArRt1TkPGyJlJX8k+7hmUBcav
IUyGhUIhcZeHpCamUOdl2PxPq+FqWeh0eFSzqLq3uBIMIsNrbSoSHS9capG15kfw
e0c+ii1u5NsjuZvjg81777PAl1CmK3FhYdKfsVGuItSxjd+iniV9zP4r3pbVCTSF
CLAGb/5BP7+kGATzhPbadowN2F6hw4wATtHHWpWaltVljlmyOgzTA6dGXT+m4eSJ
kx5gA02sldmr1e0l+tvgf03lJK1wAtSPws6bFTAC0gZnx8wcFaac2wHb8EQ8VFYU
0ju5PQUyMpYEz0QGFPe2uo/lElBlLWN0F8tGsQ8y+0DbLb0pV9pFzYL6CDg5orod
zt03JI9Eq5CQjlXFsW8krJF6vPTXl41sH36es/FIohfF9YYdTT2lCMDWPQg7oVGg
nrZbKMGmsdcNejf60XYNhHF0Iqyjvvaz92zl2uVikCD2qZV3ERJ+0QuaUg+cjgmC
p+5r+BZ/5lXt2WrltsFUnbU9uYo2L/6oEvvtIbdb29gRn44Hu+oc0N+L9iegivaQ
9dkdRZXGF7/XZ/QLjondK0I0ejqUEYuF0DpQhdd6+WJZmPGlE62MimrS8rqjYMrZ
3rLShk2i77XXBz0FlabDEBRQFOIIJeC+SFnKzW62Y/Dj3t+iAQ7dMg4QbrGcdaIe
0j6NVJ/6bQk8IQDVkQwhTNvrCAnkcxq1oWH2Y9/yIc2iA2+ogTHNkJ5RX+aRWQSh
o4T79KGc7+oJMkftrwHhFE4w4pwTDqLePOWhHD6ayBWIqndM9DQpIF3GAI94mT7v
xuLhWyRNGEpsoFU6iXqE019prlPZhmTS4StMHJwqAp+/C/kcjI4KljZ1sLnEXkLp
T5KG3eOyKQi0AsDfC0f5sN6v7QIrqyZjt0rCyZ+RiCDy5+Waq0N41r2Hwj/nGef/
Mk/10XyZ8m+Ok5G+yPk4RGIpTIW2StnLeqzx8yUo8CnB4L8rRYmEe/74BDOQcd+P
Ow7gdYe+Ai0EzS0PRNltNzRGFiTb5bZ5EtnEIPOv+DdTQoVXc5P2WeXWNwU2rfTq
y37Ep5VYd2HHkjjfQgzooRQVxzT4N91vxO2x1lkHp39c4X/0OquLwb3abVx2dZQY
Rxyn+L7i3tbqrAOb7I/jYOlG7hw5YUhm11ubN0SEqXJ0GU52nX69TuQBu6sr1Ev0
07CDdqGEmgGhYe56CGZE6VaAJfiWb7z+vhyH/XKbchRXrYnJtbRjf/+5ERmSlOvd
GZL6/Z4xaDZUKuyHU/LnsW1KZ18EWiFehrAQ1dwmFVQk6VVZYFZc7mHsuMqrGTsx
rOwwYiIxihtxoQtROoop0Yio80gPRM2j7Bt0ISYhE4iv4ERepIq6QX/ivTk6xe+x
/IF0YGwlYcg4IV0rO9R/aLiK3wf0T0Uu80erlrs5fWI2RMIgOV8wwwooeTIV1a0n
suLdNejH9QL3N9W1LVMt2Nc6JN+DsNzJhsIzVlQQznLQFkN1Cn/N0rrbIlndhotO
vZnrKh/qQcLOgjSeEa7lZYNIvepEnykBt+fi6qa5fCOJ3670Y9Ozrc/xzZzL5T/r
IR3VQshxK4SSYde8WuW14s4G25m1NEIVF/x6gofOWdUNNPrB7Rg9P7VcnXx/Hx5Z
L+YuoCAbjsSHr+9mNUSklXSc7vJTwcWVHfhc+Sb5XGc63DsswOikWateaUauvfSi
gXPDrncexIj/tabOJELeaOYMocQWOmMnAAr9/Rz4Kk9ZkHsZtOSH9usUR2yh9y/f
+WTGMbghwej2eNMI5iYA3uTX3hNb6F7QMJ7vthYsulHENYXcRht15x1iaSo/mKLt
Re5DbazNtBjdCiVLltCVV9mpcj02sxOoPD9YQKl8WYQJ2bkZ8YOpQDhDmGEk+O7Z
/dG/F+oCD6p5fCv+NU5JdY7f3nQs3Kv4h4ulLwWVeIXJDu86T3iE2rf4eV4oaS3u
hArgH/vej6VxCM95rpDKRIiBx0kKJYhtFIrA3D7ahWI+JnmQXjwfh63PPXOGOHbS
xmdxv24jE3+u5tghiqqIYOuLtHX8Wwj6aC+exOXlqVOWO1zXZQHHe9NRfxK4H/lA
SZyaNti6m36tU4HmRlkpV3u0mvdh6nCDy1h8C8Z0Ua+vn4eKV7+AtWPBPQwoMOKa
mqbX6Dr69HXRj70fxB+hiIHiCVgKQo64j2mUzb4+5ZERlzDj2hyHhnNOo/DAdjCX
oHdeHa8WeuQvD2x4w6zGQM5fyIpiLcYFraWij0vizBhEj4lsQpK+T5OMluuwUv5o
g4nu2l/plL03QwVOfxbkh/ZKDHxYNKZi2aMDCaAtPI3Kwk027CnjpKi4qxO03Tsy
BmZJF2wP0vJlgFjnm05NtLuth+KzYkDn82DfxC8E88mhPtM98S5E1J4FSblvMi0/
LaFqdeF+ISU788t/31D6biqP4xO/868voL/HWTHrhXnM3JbOQhBsuZpsoo4SqbEf
ytIqtn+sJlvXM5sSuUts2xYblqvuzMapKYKPnacqiHhSDmr3l2+K+d2Plb8IMQ1F
wDcWxSdlQlxlR5DFedTRM7Mf0wrWPch6lXtblLNvp64ITeqY5vx/xX5agsiRrH40
hfFaQE304x91lqn0hqyL6sKS8Pc+MNfFZr8Ds8/+BstKmavpHYNckaaCAcUSBmUC
iVeKayCffBaw7LYd4o5s4jNXUJIk/DBZz3JelZz2MGunw+3p2kAk68BZ1S/TZWKG
YyhCVTtKAJD/5Kv60L4FO+491rw6mayZNC6M32/glwCiVorJo9ADXC8s1nSYc6Qf
mzy0tcZxkIbMACYFziITdd9P8dfyNuDa1jLApa+9uvdPiuw4338L3ceOvSYBI+ae
LXVbUULVW2KFDEXdc7uFDPp9Yw8K15ibfU3JOmYRVJ8KyoHFk7jLzL/WY4WErD5V
9TaAM3CWuBVSSkphBQH8E7WqFjV4JRXiVtCzD61lEDx0hdSf4kDfPXUQLhHzG1fj
clRcj+ajGWtHcZUqos2tVCgrjEyFpDFX7Wky4a5nSQLS9cuxDPauPNnSQOUzh092
5IOfODooy/HsdKIXj9jWxPfJpcj9tLi58ZWLrpXog9b1wAMapLVhfj4i0+zf38Ws
Nc/0A8cMfdrYcKD+PS1olTcGpWJuMm1khFTJWtp0TlG8e13MXdzAU7IUXxiGGi7D
hcQ7R9M0lc5OJ7ytRAr48iziIUC2r4ur8PmgDpxZpEcFpZwiSYzdeFWOOzax4qEG
Tv19ywN6LlXaO64ma3GmFOX5ouX/AXJWbuJBA2TysNE8IIAAOS46OFNPmFlHcgni
2ro5MoWKNsykziPKLRqDEyNBTrfqY7fCz5+8X7rE78jvxC2OIAFfwkvkYZW7rEAj
RkISmi+Gfwdjd1kfcZBDHiHhY254EiDs4pOeFD02HUG3eZ3Ct9/cKu7NX1jW0tuS
6nNAEEo5+aYJPjIzULjM7wE4aYCjCHGSUJvXziU5Pb0sYx7d8sYoNPll5oJKUoOt
3gb30olFYffIEZd9oxNvIM2bcsxNe34vMigUPJs5Bgm/U0lzTzfZxvu6JTIC5KXf
FVIEzJj/ZDKlS2mcqmEntWntGXq7gTLVKgvumxY9i44nj9T+ICo5zuNidxaJdJpf
G6C9JDPsQzRZveALo2Oe+MY4mTgkZeTxIrDDa4HCBr9flPP1sZQrbQmH2szzGELS
xE8x6+bn1t3iqfSLFflukg2gHzFj/dgocV/F6TSvF5EoerNGaSEGONAF87kg7l00
WhzQ2i9ntI+G2WPjbuML9NCw0DUeYZ0EUyneqpftZ7qGey4PXWdZ5BB3iUytq6bT
YFKWoYwWx0hDWyxESIBaUdiD/tgFafKbmYxlmpsCxM4/hRpwVf+atd784ROmu8+H
2/kQm4B1JfAA78IaINkoe29y9BN6xK4rzb60qLbu/EUNFGmoe9outfPqiiXetwCG
B/qOdHQqwLtipSDNcsZV6yXnHradImaFR5XKvrLmJsPrcyw5j5kSIv+zdTR0LbaH
RqSQmgLxvAvd5aco1lLeGVfyb0NhAJ7tJXXrFshdvMHrSQuxtiznf/zTG5mW2t4Y
R0j9DWIygs3huMCvu1vDmTmS1ZeN7D3OOHLkud6H2PajM/Ta5q9qx4YJFeFHDZDd
o97EKo8o8HhTvnmKXIKJAIOrR6hdsVWJQJwuUtcDWbyWlkLlExarvyZyba72M/NJ
g7jhSFI+ODZK9DoQ+Vq9mJos0fshyvDb1jjfPkEn/wdAYAYX0YN0ipuqoXi2ZwT8
WtrYMhHhkIDRASmRhbDh6TY38o+u9QBnt4H/PrD5jdcgItB+7gPKr7TDnY5W5CkY
+77gumjkbevtgcgD/G5qU2OilWTMgit4KmBY44sbQUkYN8Ih5trHTBzsSjCb8XjY
7ZB4QfR0X5BX/iQ+xjoa7Tg7udmB/amgMU6O/xiEqfFXsZ9zYo68hnrNpAw+puNt
jBE+EZUhbLQiop2O8kl6bg==
`pragma protect end_protected
