// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lB9y2nrB76PfFyxesEfjhSQzAtJVxQbe4NVvwTrpzpnMgopq6W2zD2LfL/+n+wNs
VTTU8HyPBp3H4bH4eLizcp6Lo/fEYLVyoIKSvheHCY3Oc5zpBPEJdV3lIKiTEEGh
spaRwkzZ3nb6NIHvFtGlKf/tt65NxldzV/n2EnN2YAc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 103472)
GF4pKRYCEfbDDGtgOslGjWOr4NXHKpABQ1zjxRaYAmohJXwkIaFnAM3NaoAzt70H
rZWjiwtqHwqQ5sZehUu7HW58rgz/Ru5eWtwWVmArNZLz2jKb3u1qrV6MmpQIA+hZ
jB/9T9DHfzipYN8gu9JrySBR1/LCWmSG6+eQZlEhqL5WcJHCfDNhpvqTxItqckv7
n6qkaPvN/DONuNqMZh0c9RPHA5Ow39nVvWBPZQynl3m158+NNhg2d+837IZhi2YL
OFGD0kuIFJfzyhml3VKLQqXcUiUO3keruLdS37GFcaZ5fG1igEqor+2WCrHg/vE8
9x0Ol13zBogBdpZeWR7S+awVTO02kNpb4TA6aYTefhFXQ2TvB59dWi54Xpi/SCpL
34Ci6vm7vPKOQVYwfN4u3EYZ0GqmqtwngA2e7f+LeSBKOsBOpAywTjyvsemwKBvl
7/2nUsDFW3i+gjp/YlpueirLdSNqW2mOrW+1zspHz40MMkPzvpjfii7LDW6DlI4q
icNNoc7ewO5DFvk5yfSgUuRDC91CX8QXAkILQCPiYr2mqUCT3XU+T3aehDN3G2uN
TfWiBYFnXj9sGgOMCQH+GDp0h3uCeWA/HahuydWsUoBNeh/DHfAbnuCMI1bC+LB5
v5SqugngKSZnPNHu8zUzGn6dy3NZ73ibDObhjdMGAVTW24j7ch3gkbZ8Jp5ii+M/
YTTLgbC81ud4kr0zFEhKihd5eDt6PS6tmzl+Hpnzbntit3/gg4ub4ktWpfbjWw1d
bF1Jdk/9jKyl9Z+x7pXYIjPS5nZIaLegrQOz+tekS4Hd5o5Q37wvyaBxEjZN432Q
xFcLDmrp7gYT0JZAjcAesbl8t+GlloY/as690LZKqk0I14A5gvi2qoOOrvbh+RQ/
xwNKfkqctquyo+a1ISTWNkbQH9PUahQgT6nb+GbFumGeimBimKtk9seHClXEBNQo
lJrIwaGc1IfRCmLh6P8w5UhUsCiZyoucLGKeLEXc6ezsShLQnTPyKyNnb5RCKNpx
zz/vali5lNAC9LNTOHgB7AqLpf4njf7a8pY3dpNRESumHykI71pwHFChu43kb8J9
XXZS0NWrckCxop5E1F6fDCWUtunbB8GCskc1DtDKuAHpKqW0kfRBxv8F7o8tCjO8
BMLAK58VQ3xRGZA5AM59f0CZvA4TFtyzHl6CU9y/V2+5pVgz1M0oGntZaAGPlKL1
TjYOH1/AKKNgnFdcsy1TEMF6iqgR+QEPtc6UoU+jcroVyL/FNFzc1ZJg7ODgIW8w
pe4W5h7VLpo7tVal7RyAFfqRxOR9w5wo2CwMk73iTfD4cRZro4o0W0IJXWQxV+zJ
S1gk8y5GG4IAHV5Irn7a52leA+DstcS/f21Wve3em5Y32LUkR7OZJ+7A+CihoJJ3
NrODgzKtZ+6feQZF3+j6Tp5KhpKv6rnfV5L+BYErm32EVdJ+j2s1b9UPuiM679/n
5uAzneZ6UwigxCp7RxO3wKK2Iutk7wtrBtKopk6FCt6BWVk9oF3VF4AkmW16KLBH
13fxKi8GM7qKlTtYIqcfzmVG6yDbp28DNmuacJhEO70W67ACZLDhEWN8RCvxOe9y
CLP/pku63P1ztZ/N+1NS9mt2uEeDV4kS7Vzp06z2xKRfeEsxeYgvApKh03xqHv1t
uJ193Q/PrUIXhhkle3i9o8VJiBxrHixT0frffSoV+T/tzIcFyS5qu91g/Q7bpI3D
o/fL+p7YeU3a4N44Cu/ygKmGvoGPfCnHzrEC3MO/dxPhSz5iDanVOED7wZutdMsM
O9+rCBb917plqD+8MV8G/Wi/F5zme4NpnVT6epQQo0/zx1dsgTlZnQqLlAYeVuWm
745N/WuzllmBZpfaVwYJbJ+iaW0S02+t4HW0Wksfn60emGBoUkCu+0Rzcqnu6MeD
NwMdyiuICmd0Ck5adPJnkXb/KerG2WMZ/aNN9PA83gXHlGUJ1MDLqVNrVN2tfXss
nP+e7nJly+g3C+xsZSlal+jNwdBiCTusfJ1sbplNyZ5gHc36ml+1OENwpXhKNP1o
KhXhaFnBMc6VUabnta3Pl/La7+G9fZys3q2PS5+eJPMi5o6+FNTJrA+OnmQz1gKI
+5crNx/DW3qPxU5qecVkhrB72cEhfelpKPIrarLqXILA5Puj5bJgDUwPga90gGB7
Jl0CpznE24KqhPNQUrdCBj10YTycTX/rHJYz7+4hL03Udqfvt/BKEz9qy+mxrfjL
ItL+2HKtsnMss9Z9/6MyOhZA6PpLwWUIkm16Jy3jRNhdWq1MaONr+PMbTh7Rnu+Y
E3WvmTfYnOYpaHSINEzvDBEdCQ/n0UorBwOQlZqPjPZP5PZ5gB+AkOYtjHh8QzNl
QGblO9t3XODdT1ComerdzLOYKBJy8LoXHlXODchHDIfK4Ip9l9MNiJ+1Q5ns8cjh
1TwPx0d/LkISfOum5GB7LyxHp1wDxk8wV3yrW9RAVYsUZPUH/Yi47/6LG4/AZgrg
6yDWTMwF9HYenXtDNFUhug5a1iZ4f3G/7MXtke5GqYW34k/Lbcvk5PEDLErfwosm
8xmLkFmTsVu+lID6d5qHb0F9Aq1B9epn1BoPbT9m28pnJ/L+mfC6OBeF3I5DRBv0
SbXzbStm7d9DeLTIwsYlw7pWif/FXD7IIssVhRlYtYeH1OqgWOItltctcO4ZvSfd
WWqRls2a2vRP3Lat1/Vliu3Lc0yNlAxAK7TVbFd0UInywlsP6xPyaDrXjZA4DE0D
J5fiDMLZ4/qeAeQS/wBTubVrTKJ+5ZAhPn72ayXX1a14Cr4BmwZDr/oqimtode2F
j7wsiqhr7PicrhpOdt6ZtR+dbdRHhLGHfO2PjP++DdbT5I1pFAs4xm3FPb37b9BO
bK4flxzgjbNfzZBwflQ1Ys0dhhLw8oUPglqjmAG18cg4OQi8rEGOJAHlyxRBhW9B
zOJK51MwvQp/ARX5nGVsdEap15te9tYT5akcl7jXbvZRA9bjvRcGUsHw4s0x0Ehi
aDl6FV27IbxmDkFF7SxO61JA6iWF3rdsCip7GgjFywmTCssuhFFxIob6Nk/Zy8r6
K+9niax7fqdqgtNz+U9VGVaC+xSAYspx0y1s/jduOz08/kCeLBgWYz/DOEHreC6T
qg3s+aj1JEL98ZD5D7/5XHV/ac7iKSUYEUtjrfqToidJMbHJ02BphVVe4YUO5V4T
FQAWlHzH88KyOW+ncvBI8HXrMt/0jhMyxqNpPbbEZDoGLkO9C5qu0RdNx937p2Oz
FU8mCAGsMQ5GeTbar32tV10XlTVgkdVAAETCouhmI6KESxCtx/vL1HF8eYJjouuI
afXk6Anc7sTQCilYPuiiWYqA4OkbrU9MEeLybUpxY2M1jXAmD9Be6pby1HToDU/w
Qsf0zBRok0TG0z9GRRkBtfkRdowxJwvZNa4qtTCUzoQ20p8DaVrt+NZvQjvInVsy
25uq4kvwcOMtEtM9Y0VrBvXrENOghDy37YrUwqKa4x6IBTVPkiH78xTXLX/c1s8E
UWJc2ZLOBPzOXXOjYEagnL2uJ/lnko2LeUb7RoxTRQz6yuKIPkt8w9EXxZBCxNnC
xztC6hAfD2rmeOlOu00YqLLHupD5tlQoCla41T62AX1jNlaRCPFG8Fxz1XN23O+1
TXoyr5dpzw8aTT02/wsUSO+5/a/TybJZEC1RjlXThj0+74tXyXlmN/S5dngPsMz/
GcCOYUED8fa1M/EiBhfm30QP9tbYDELDLe6OGLclEdk6j5IXcCX2vLwLgFw5FGmh
H5W4W6VOfN4GrI5PnF/fXXqxgTLl76QA6y5xViDiKewmLqKeGLy7GUaS7MSyDihr
lRZu0tZLa5Q5T+qRr1adBEzshYfG/zW3HPR4A5Kd2XWFnguub3za256uhSjLpt2p
DlfmKJjwVTnNdAqe9RIOwysTwoZI67XVIlELdsNNlnwUE1h0VDBGaW2rgrtkOoE1
sDkfD/nQj5P2GSQGIIj43fakylp92lKo1O85W/UtNCq1mxWSldw+gENddJB0HZ18
I8J3qSZOkig8kmkZQ/SbNHMiDngnYP+QNxjoGGG17JI6QyaiwsKkKv8l+34brSvD
zexCjEoL5AkZFWEfFTp4KyVDVzgu6LyvS/h6fsyTEXqSAsvC+EM5maXQ4/fzmhZ4
wiVt64m45mLhc3mS/ZRMqDTCZoWJ0+e014TU7GOS9a8jFdvNcVVwRQ3FgOuxuLO6
3/UcNXkQFQW8zQ8ibR2/GxTWbSuHs3sYRm0+E/1Vh0G/s8VqzQxYKUv6BhTFtWnu
XmSPuuZa5NxV33SoubXWB4fctJqjqVlZwIVas80N6XpdxODrKckweTN6Rk0wAcnb
1q0w4e0eS4Dy6xqeC925rNvXqtg3Qdzy25li/clpXooH4YJWyxB76VPbWrL/RLqh
3JwDiszkDaX5Csr7bBHeNq+cosmva/B3Rhaur2d1U427sHF8CkKpis1oy9RFqkwk
tfnw+vRXrCkO0lpes0RT/x2S1T4oXI1MjH4agFfgWXcGxVjioWG1z61u1obOQX6q
aWU6jE4C5awvBdTgXY19N/6Nddzm6oZ1kGm1/uje2AyGAYrScH4N6xP9pZE2PwME
uMxWz9CpfoaxAoNwJqdjjCZu4iGmJ5ocyvOUcXQgWB6Dbcdr2/j0HF6d0HeNM9Ga
N9kLSQ2iWpVT5YE7gZF9W9nAXXKKzFKVSlkIgMOuae9G8CABv8qXrN9LtLOVuTOk
EzNVps+0uzIx8HFhtJ8nQKj+oWbGQr7q0JGQn1bObK53fViWP66K39UMuWrLvtE8
ME8tq7p7ALaGxLnfQEzwvjlBv2whG1jW7xSKuNuvOjHjHGEbK/mvwtgqsQDVoZ50
evVgzkDj/3Q4R5Bd1ToQ8o3bVQpahra7fvbshHRlqbCQHRo/0GYwOLra23XHr9hb
mVLByZOLKn7V7ZpVIqS7JK/gkYhbeQFvb+MyAzNv9xvGhY7zbsrnijYzd13SD53J
kRycILOFmXMMFH4wbycblCtgP29sNmMYmGAtiFKgk++23lTwEi80g4+9jRHR9esw
v4r4v+cLhZUn4zjiFPwJFaTpHDdxjzGk6wGcc/lBZKyZxnKEXcrNieLcNUe/kOYl
kUmSthfNzk9VPkkiiAl/dt3Ks9qc4jmpzHUlP8Jma9J3vr+vvVIwC49+jmm4YH8i
A0uGJxOhGXySYx8QIhTmkTZ3/BtLE+fsIskhN9F1v1/sxRgdAaqyCPopJtrWML6P
MzNCOdsYngv8fgmdk7FIemEKlBOldCwR80lAuRIk0YN8lYtl3Q1CXEZWEFGcYYbj
Cma/ZHPV5zslF+B/VD1cjxoQZUpqiPKyoz+5RspDmcznK3S7vYAsa8XZBsfopmGx
/b5tpFmcDcQP07ZTqMKblpY3BSKkjLotTESzdImRVBEtNCEEAydfVqWZ1xj3wMP2
F1Qvu8feFNoJXQrZlnRf++ZxstKBGmf/VWl1vZGfxaD0xT2hMJL+Hon/HZ1+STcl
DXi2h4Hi1mPTSIRDYh0C3pdkgQtcDwOfvxbmTA6+tOC9E8nD1ysGyDAabVrH7Vv3
f3fNoeVTs3qVrsmEt2hTaDD8ptH7k7ChKsvZeRRsdkVoYFh/HvoCZxdFt7XvVjfU
PLgcyCJrh/4/JA4BljslmGiCijJeWxejzUmb4YK8Uh+ZyVqIGYonZoE2eSufVrhl
aTJsaEL7maqd4VusVNsVcmu8NcK0RuduHBqAJvHS2/zeYqOd6uuurLBuMboUGycS
CBp6O1TC4tn80Se2HEm4EwnnPFc8tg5dpfyA6YW7GQyLVJAWiOe8Df3mA2JwKlLT
P/yk6z51iDL3z2ZKWNLfNu0pDUO1egjTwqxgwuaRA1w0j5KdiTDIFHhCc/SqH008
y0lNOLTNdxEkZMi7NCaSN9sVnAWgV+6gij9AfMyl+NkXKtaay5xnRC1hRiYInIj5
6Z4Byg8w448VYGD5FLX0MSeFmsjFGOeB86d/Ynf1RGE9J4na3FCXrEVc75N3Jf+U
HvGLoNzv2i81NpALWsNWLn4skfxrYPxSiIKRJtOew1xd8FXZ+wo5bjLnccPCp5Cg
gBWKdYLU9W/97GXt7H0XsYSmZ504Q9fMcC3vwjA6pVLK16tDZ6/YDoQOiT8YEYof
0k22mQHoah7siY660GhuewtkHibRe6O+qtPKhtaqEKjn0+Zl5uxjx3mlvXLtN0XV
naMBDz9M8q2ykwUiFur8KfkB6yTjuksapCfTwBt+0YrtSwL8CMrzZSFGg4YGZVk1
n9kP+DQl7uyVSqgV1WPUdFH5McYd6dy0TrIqx01BFvLPmJW3BoXuRXC4UqHr17S/
zd/LilhMts1VVwlUtrjlxm9Wnw3S4k0uYDGQ/rwKMtn5YiPYsiLMxrZVDNZARjDy
+JXHE4ZYoXtch61x5aQz+yiFFKBRtBvUJTb0ZZEEr2Hseid7V3hMwSaJXxCP8cqL
hcu9Q+v+HAEzIntskiBvUGSv1LdoGkbEViLbvKmhtn1nVnb1PNsd6qZUNerTgHVm
F2dZSxUqynkHlxR7GU4/Z2lwlLAR0tqR5oj2EOhV1EekdovIXaWCuKe1GIzIWMLR
TUru8xmZ4Kv82JNkYyO8BH5G6UwFOLnRgwkyRGAfimC+enY6ebmIsb+TaYzaaqSg
OdQU/rdtGUo3vrUbl/NOCIjYLN/+ShvPaR+UwZtO8zBNIIQges0H3dV9dWanSujD
33kVrfiJD/YmNOi0QB9qrwXAt+xIILZwEvN6i/SYzQcZYIN/8draglnrJtM/eINn
SeedFBN2neo4aX8BJAdKSGKTqh1NOx/wBNU8eLaTIRUES0qep16Id7x1uYiOD4Ki
W8bmiSGwUmIbNRJYnObeQjVO11z8Bk9tXwNPdH/bF8I/jSjCTuErYypzFi0mPEgD
BMDx2rKk9mB8rApPi4kJGacd4pxwvi+xtprkIMPKBkD32eUdr3GLOXKIaTVGYuiG
3PROiuA1F4Ns0LKyh2OobHM/uXUOuwS0KgRn6ggluGnFI6MiP+DTxHLd8H0YPUxr
00BxDYyqQ26+RJVdzJZwLylyLs1egnSQiNrvQZsybXC6plIz5vewtX9uQ5lSHVyX
yPVDqsjWR3nr5sxttubAJpJ7rWWYN6NqmdgjiaX91vwhue5XgG2g3bs8ZEpcWMEl
LgdKeBr9kQi2BHIA1VWY19Mb8XMTDPh++09kHqq2Hqc8AK4vmPEyvOPcD0uZhFb1
BYp1E4ckASzo+Fmw8fK48ZRLRHQ6m+Py63S8ZM72hnJvTBOGv/qbbWH5sv6zaSex
aUmCvtHM0NpxeTje71UyqrtuPm6QV3h7q4kJxDGGuRzRZbRxFIiuV8Kxv9Kf/2T4
JPhJHhLEfc5K7hNPbf7JTuieFxPRTA1IgWuN4c83XL3qIJn/hgMtJrhDv+iU163I
tM0MMeEs/vCWNvD8bgRHAkdIFTWJOAzfUFFJsYBlRlPBDydJSYg3UYbTnZfRu79n
gU1xlVVv8ejtMg9h1XCEVcVPs4ob5W/T/MzUUfjSVK6katQ/kHhF3CY2yNmYX1sL
f3zdqVc++UHEhmxnvk2MB8Rv41YQi9kLOOs7QcEmhkmPeeue2FmFEw5wbGVLcv/o
5jWsFOBTuAWkN37Cu2SmJ2AEvSgL429KDfk/7kVl6t819ck2Q1f1WqxHmpqcNfOc
/ALxcbvQZ9Hhwm05kBhg3UvAio8maoDnh6YRnCGzskQXHfDXGAujs63TaCxqimmC
2VArqbP4A7iYpeA3X6bzxl2kJmyzLv8EP3JlX+r6LxPxx6H+F7bFXNCalrzW26Ss
q8uahccQBwtZZA0/2IO+xLYJkwwCWLU9c6de4afD0chpRqNo86waUysenNc5Cq2O
458V1vphmtj3FxEk7FMyIRIvY/FV8Nxkm7LM2xezfXnBFgfzW5HAC2V9jMAv0hK1
LqfYjz0/dVm1RO4aYvoiEhBtG9jtP3TqDX3XhyKv5YdFAVlt7h01o4TpX5g2w+94
0JzRxXrgsY7EoiE1qOWZ8mryH+YeSiEJk0/tDXlgaI5yAaBQwOphzDoIxHJKc8EN
DYWzfKWo4DPp55G6PzRw0TRiqyyYvLJ3Lw7XOQL2XPQFxXm/qMxPorcZp0jrXYK5
AzMdoElxZJ4AQQlWclGOvCRifuwTTc0PLZbxKz8oOwGqJlznvb+TKOJDr9Hrq+jh
1PfXCPpGe4LFr9LEtyyIY6ySApQWBJrNsjQuMydgqHkn8wyyyVAZRihb1iqQrAlY
rSReOzHXqyaoVObfUrfW9iBcXLwWwYPA1yLcXkgfYyIez0vQc+XfYHxGU5ltuOH/
JvjizAyypT8wIDmRh2e1FKxTWvEVuW/r1QgUphUcdkPMi2akQoKdDcuRpFJHas8C
R6rnhUZXcgSBtDp/qhPxe/1ytfvgSy7gUpGmYJ23VldthTQByLMZc1KuGXUw/rCr
d9TWkUbZljWSy4/7eR1H8YWfGaZ0Mp6+AP2Yj6hwlV13Yktzp0W2e3D9LgjtEUwM
0OeZ4wO1VE6GgGf/OX6q3EoAsnGFqPhc9vmiT4UdP+CYrbnVlM1gj+L9QxnHx6Pn
aAmOUOsiPrma7ZZO4hyqmy2JTPLhqWVkuZHIrDW3SpGt5uJC3p4FlGjhmk4k2Psn
VlsdyhJh/QiqwvtKIq+h4Q+6gzdH8tyTTep4jE+jtTfNh7yeuxCgnv3bkpbxUI0n
d2G2RaJYMfZ2aWRsQ2UuSwjZHSzGG1uzg1sX5TpA3QYNLPWi6/NSDPxNhA3AoZRY
lfXF4r8qdA8xkHwyr6r7zRGsYDB0LWp+SFcVUZKha39iY3hOltsesd/QUowX8aOa
TNbGdlWHK6Ldz63jOFk85bejjr9UvkafWttlyoZ/nzv9iB44JQzrGdXX965kDxYW
5odr10NOVi6DogTKMTjHV+Am5kPvO2yIXaYtbj2anFoN1qM2R9hecB+uyRdu+keh
NvvDn0QYesJIe+u8tXLfle8W8XydNFCwmACx+aE7e1+f+EJlZJqKWrqNbtGRpxzr
tngTgwiqUO9SDVeHFR8pOxzMfNkaxjHPYnEocdVj14oti4eyjpypO/TnRdRNfA+s
EHnNoFR2xEqevr3scJZcY6nmtaGe965pQQN3Xpye617olCYEIMZ1vdZ63OKhaOZC
4oxsi7+2R3RVSJb2AbLOzTm8bWyp1Yh66LAX752zvpm8ZHD2BPAzL9WUUxkVxaBd
nMNoqG8uk36wt4QTG1EIcoEuQVs3VEETJWpD/jvvhix63+hkHICVZCox42yds6wm
rMpcCejizU1Wdof4TofOgV5v+BwAMA7JsMzaJP0Tem1Kn9cxKnJD5OGn9ZVhChcM
xwLjX6ueWykZZAcygdkOsKDRXOdiEUTN+mWS6GHWTEkYfr6y3JQ3xcFL4ZrhzUyV
wXZXNIpw2C2HGw1Y2V3fU+mfK9kyeRiHJj2QS+eJdlMenHBwuJ9DJFZtqJfOBve/
yQ8ft1LKlmPuq33w2chpIfj5uOBHDLrV9MIdYuBB1Tj9EVPg8tD/xEQrjSduV5sO
86pmXRgKPqRbnBtC/ZehQsq2uwXlemusXrVQlfGn4AX0/FS+aNl3lpXI8pxJCdhu
jz4fAtULPNV2My3YkNY7NATW34pys5EVUwwk9NjnVtRgCnlL/nPXi7sAyAnJ/9+m
66qfySdxZjlxoKNOj6hMInAF0BsitCpMv5A6k9nhVxmt8w+9JxvGVSyANdaDZxSw
zsa+2Pmq7YS9E2g4+xpvfURA+wr5owFPIE7OVDsYu8VR2vPZCngyGA3YLKJmf/5d
6gNVaz7uewiZEFamVFSG+ZlDBBq7nrycyZhB64QI+s6/ek0/2YW8WrIfj9A4AGDH
7Kjei41XvNoCdNQLoabfI8ZVxbMFSde8k9VbTuA8d0msjmHvhgk/h35arlvg6Jgw
FHGDE/wuBjAWtMOhEQ9DxZeT5C2xtuoAmENGCCHNkkb/C6LE0J5E9QPBltKvbSxf
l93V5W1o8pA2LQZ6aAfFMriPK8ufyQ0SIVp5h8rwA0UpfARZYag415IX4I3t/kc+
2Dz1ZZ7eVybat/p0eOEGqOxdu8gIgd5gOUzpEpkPk7/0dgFIJObaiuZLVkqlV25P
zUudCVlHyh/jsnYoMx9BgEk+39nt7vBgFKAHuYeRkGthwZs1RcSC/4G8uVwwpA4T
/4rSmfxpgeWSQpQ2NXkjn91YxYek+JemiiFNixGYx8ggAUtdWBRZ2z1HDRUeiiSt
22b1sVZo8yFDC6FWlYI6fRwx19jLGWWFW0GFa9SIigksdQbT7PL5Dlm9E0Oj93zd
qEFQ9HmLY9D6QqPH/EmufREF8iwflqiC/4sgYadoQPJCGSauvRzWobV9awK+hYSr
+Ys9uFTujtqUWt80Ic56ntuEyWOZdkN5XoTIguyyya5C2pq97D/8rwZ8UqzaAC4b
CmlVw5gdbcM0Ns4HHe7e575Z4yrz1c2S/0WUeGExq0HVzxZXoynQYs7xvtLF9/UU
44tdE7AQ9//74yAmfGECy1jo4y+/bzAHmA0b23F3KkrIU3+HFAd2Qts2XMzp1XHJ
qm5P9wMEiSPsHJE3X9GUFIRn9Mqs6F47IYKrlxTiQIUrLSAA/ZXdfV/AzyMS7PwV
d6jt0JutA/VQD80pffBC3Opqm4TAHUzZ46AMH4al+gWF3explXYxyuxZ3FD9Pif8
3z2Y/0oyKngDzH2iEbOQ3KqqoeHpd7hkfoREXA4OAgimZI/4TFXKwysgaPFOUYQn
aA50VAASDYoQjTTlgRrJ5jSw1F4h8/27mJjLrMA3jLjnwQ9esoUyUiWnTEudzCyo
t4xFBaE32KjH3un+PUAhZf4M2E0AwochgoulzYUwQnD9hVRDPhONbuwtC86VLAQ7
aG0MM6PK1GU28oZGMK9LFTLYjJacLl9ZH/2m+J8RZV1xbLivMr0KOWMHroHrYgiP
0kYBVYsBVjPWH8QwE0ePrsrZS+eLggTgXnTVGmEA8Ue6UT1c7uryhqCEyUFCtnus
NptgGQ4/YE39yG9eTFLLVpJ94CpNTgyKH8ZODX059GI9bBuh1fSuYQYrTIaDOIfW
2Zle/eSlDeqvdpl4dceE1/xvaCZq/IN59bcwZ5BvM+vdFRDDKAldS2suUdD65AU2
1MqpHLWxztznoHT/dUUpK8rKxOIHL5hpVdIT5kkKcn4VoI82U2rc4HE3TqBBXB3C
gsCo5RAhk1+Wk1uMZjHSgszg90bUlBW3DPkPKqo3sNURIIa2tQemhktbGHsqyXey
WvskGaxNny2ggOrIHNCXq+quNp41V+xqCrnbYB/ei3iuGhl001f6wUjG2QVnO+s7
8qaHaxmVu2ygjp9hnc3QUuwkCf7wuPFDAq8PGoGGjy0BnkflXUDAGByX7UNqXVLk
U47ssslVecontIH7ExaelV3t7CucufNeRUguB8Ce1tV8hudfnR9X8vZ5XQcZeYEK
A8lrZZuqN6LhPYUMXn+tqvjhrcW7T558UL8GuHSboAxx8sKBypRcIV4UkgUezbrV
rhtr2/Pz/Ge61P3cT8QafOU7U4ZomF7eXlBWlTL49V6K3frQhHqlnP7wjtkOFna7
SNpzbUeD1yIHx0yE/s6sYx2Fcels1qIeYNSNK4XvQ88PqInGEO6Wq+zkfCGwtZrv
iF22+MbzDOPXJkViwCYB6ntd9vO+e7sAZJPpzKsDxCtrdNSVlNP5VjyeRP0wRg9v
VQFy1QjNI0suhgPA7GFYCfJ6ivmWHKshAHPJSHSqZjQwHynBoWvFfl7FDXS6bZm4
4EFi2JqS0DHg19rV69LjE0vX37UkrJdJtlC5bSqxOnjvZtPaoKyYK8JOLAfZxQt1
VHtG+kH9TVgp/bOcNSbpaPgEwMEhxM5GWenEziUDzf+FG2X0dTILGibpTE6V1NB+
QwiuExNjdlPl9WrtegTc+P/00/h60fttLbjp+fEb0SO4JD2+JgdnTDkov7RY9/Fj
A0kz/7e6R/RdfAx/wGQY69aWI6RFw02b1ebqRhRzWW5q2XD+7d1f9wwnPZDRokpD
nehrhMER9uZCK1idyNFgyPlPh0kUf5m24cTswH+g60f7fjBL/z+ZPNO15XKB3Nv7
La5RTLcx7ilmaKA+9hhSh3KhBJR8lRIhqdNilp9hNzMI8zB9HyXNnBMRUOxm7zuK
pZ0FWJ1WRPRUOuvpRTimk4NVQm/t1Vvde/a/EFwsBUfDdmtJCxLejCeLm2kxCV6N
mX5DCj4VaTxEx0de3/gYUrSmgfuDxYSDge76k2XmFHDFHiUbqs+NPegYkvgNIlGZ
Rvl6Jnd/V35FFySAH7SRDac/ciSU6tkxQ3l4m662zCcESCVXKHdfbFVmof9BBWqM
1EwiWwN07siR3d/f4K1zej/ZrjDIcAYFO3WcS6puvzM7qbtsMTL4XPGHGHsyyV2w
o9HT5XbwIXG/7iKvysVCu2DX9ceqZcdA3SkCcU6pT2Of86DW5oE1cvyxXnGlCqjb
TLyivy+Qs1/krdb3vXYHWvjECV86OMHEFeSKbvaeCteZ28XbKbk70HTlTlTeajwH
+hBUrvpSTVNRWyexGXNySzR3nFFUnw5TvFIU4I2LK4iny8SpP1MJTqrrbYbyn91n
6T9H+EDRpGq3a3MBd26jxU6/fAExLwj8Se0Fgfv3dqNM8+c2yWTbXljfjxaFH4HU
9hEH7iYczieo3n2wCquc+4DrBTwUhs6fstLCZlh+08PQYimFG0DTyofrt7Rn8f4T
QpMHLnAn9MfQyCKpiciBD5S8OMO5DHzu0LThVxMlFkUsiLlRy515qRQZWGTNvwiq
ZxvotN4jBDXprx6cJXKQj3gDAZevZ/fuC0DqHHvusCfyyBuBevYNlKRei6cKPTH4
t7hfOX1Bo8KtPnGU2+DSxq6Guf66m6pY/tXjFG8KgJ2Gj60JMvVkiXcZyn54hxkV
nKMptQpyYNlEOpDwqWdfGXTbZLheu6IxLC2neH1WQGI3mZ0DtRUNMfOIIF2vLlIU
lBZswfxZNZ4/MyoKRIPgp5kRzgcr+b1jeuRiYbw8yXa3rhAnm10hX/A1yXUTUVb2
CvIyPVsFWW5IjU1/DIK2aM4q/v8Z7suASC/4c+mxQEW3j2UQl49cU1iuW9f+cCFO
I2qFh4sDkKYa7Zi/2rRrY+GquU/UDUMD/TqjywH88NSaViTvum9DSSKwesfiuwiO
cF9CgBlNdQgp5P+/2ukKT1ktUFmqFCMdwi/CyKoOtLTU4OowOdRj5ITpesPqDc10
S4/TmmPCRScMkwWVXPAQxvzud217ocVkO8wE2i4mmIJSG7YycT3jZmwxHlqQ+4OV
EvpGL11K56RU5Lm1FPMfA4/0pzhcLOswWMi1XFJV1INBCiu2cMze+4zq+9JZPxeI
59dfd4dYouQghlfSU0lLhT6gv3HeqOut8FmtmaLRoh8iBQw4GqejXGOpFCgJB23O
yeHg6K9QjZu39q+IqtZhuHfYzEdwO97ko/211uwhbjpazNU0R8atx6314E5G0uoR
c3Lf7M4hQQqWGpgIg+oRIZ3H9ghgFrIVdup4z6dTv2h8bKhPDjL34l9pVqs6wlq6
FP+LOI74JM67wMXjVEpvtOpILh391oGkyZC/JVFgh0fMGQcOon9sKIKp+ZdPRxOz
WqtEBll2U8gN+Yiy1UI0/w+Yl28z2YqEGIUmotxafk/cnYv0uSDpipLSUHk39tEX
B4f9x3ODPCsRG7Af5seMXKxxKMPuz8+F9Fh52OoY/mrQPrt3BL6RP0/cbdF2B3w9
UiCSF6i5KYAq6R2Hx6EeXdOrnv/mhWBysFQUtg8TI+G6L9lWZbfpImmsZ4o8D1FM
b0QuyvidTosbLbOlFeNv7z6lx2mUEwpWvUvkhXPQLIveCIQHLQeOXZU7AO5Ic7ET
R0xrf8iDe4RWpqZHKKdrvZmrue1mSvnXHHGpKhY0iYdvu4QDUvkv/9uMdAcUejv6
kw4vK0myh8qmWHhe4BaV9okcMLbciGHUNUq3NGwsjFgF+bf4D1YRuVfZEKQrLsm6
fPy/X98glQctJO9Wf5Z4M1Dn+Jib1f8W+HnAkMJmsk0PKijCSnfu0RySG5WX3VoW
vwWOjcElIN21h+irKqYoe1RPifOcoqCJUFanYMMMs/wQs1Sl6oQsrpTyZLhctmFt
GiTvc4To+/rUQ/A0ZhWFLZo20hPTewOL08/KyjnEmgT/5SGo4OzJrLwpdyuNQRP+
jjN/0lOizcqy+ksDfbGoIAZprD1y0L5wDaYIfhpne5RVd9Zz3+W1+EyFZHCvfQ5A
6dPhDXR5uPr2I5QJQg4V819CA5sWj2x3uWo19uRzN91kIcFaG/dsgg9ncPyeIvAs
+ZSDHSScm9A/UlrJYNvUkEigmrQO2vGqIJVdNfTeDWiRjfOE70ZiVhxO0HNmH7pT
AamFQvgVL8xQa8vY4JbO3iRQzwa/T8MY7W8ZdBnouZ4HX8Rgm+1WhbPYVLGqs00M
YaNS6i0HVxPa9nE5a6488PrBA+aAFXLwXfviJWdtVegPFSZxajAaNrYD1cHkBLYR
S+MEfM08lloDyZzFtzc+/JHt2i8rgJf3b1u0IWpjwb/IX0M5fcYPZu55UjqjAbLq
0dcQ/Xb9AyMwUQe8heGdozZLrUicGrITThveBn95i0wLMQm3ICFWbG7e5wgOY8iI
YOLfd1CHHiEK5ILg3//iQGCTncdBVRNXnpSJmLVMUCLJNRqUxYVAr1W9UDtURBrY
cBLbttHTubwv7SIDWEO8UPfltofaEMOWhqI5AE1i0FIe+oEEI+qoPNMP+Umxbvc/
+8fwhtOPPQGNtQN7I32zKZuFBHdwCZSHsrVCEPNg9TLTl4hOTbgwpm0mhePkuaWA
hU3kuIJ26cRZZhK2FdWb05mUOsKHLQEc6AWdzXaM9R615tXwNEO1DasJ4cMty1Es
fHNQhGmyode6yCCqlQXaLtCoG1zIBc4fevETXBYS0+znsF7y6cmRnf+kvx5IkXNr
Xkfc00bgRg5U5dHgI48vDJkrQ/EZZc/FusEUDDM3L4KXwrf8Gl7DtvoMukAii72X
Gd2Gkla5LIHGT9iJ4jHHliPKhoFkLByyIC+WMazM4QmICHCNnzCOaB2vie3WPMzw
ZpH3kmq3rdqZytsBlcdBVTsJmY8C6fXbZ58nXgeyFDs4TD6D7SWkGvw9P/zyyBcC
CZA3910bWX1puY8JbFlKPQ0C1b1myF9VA4U/An6tX6xGG7/O8n5YJ7XuiXgfovYi
kU6frdqn5CemZ6KchgL8SSOmM7pbg5O4x6fRMn1ZXn4extMp6PPxZe7/0qaW2DZX
GWuSjomHTispYEaECmLYz7ZypbZh999yxTRfR5oslVTV/6X6QD6EHid9m8YUbNeq
sO4BfvcFJUeWOdOowKAzyz4jBPv1DRPDKwLROgot7hO6Df5k3lHhCmEpNS+TsXiX
R4rbo2ekHzc1DyWY8pMnzOUNJtgWNuxmE23cxV4Sj2pPh/oSIPRKPHGWUkD3QUmq
cKapIRCAGvAAexZ0m+xEEZcnSuC3FFhbnOnx8vZoN4qMDZe9uvBPKmemAZIt4bgG
11jrPvIsJnH5tg5xUirjA4FMiKM7vYsau9O0umoycvAhBQbWfXCApnYPcx/+7y9Z
ocxg5LqAyxocHy3p6AGLK8TPY+3DshE7OgTgXjawqEakGXgDRoiE3/QihFGnIh+x
l1Oup2IX0EKrHLdLpx+zraJd1WMuIox1Cq9iEXqGf+KDVJaosej2WbdWpgwtaOZN
Z6CaHcB9mxPczWdjLNuCDCMV1rRE/5KDoQbPRjxtl89jiKviVSxDvzAWbBkNDNWT
haIicNEficWn+Py17gnuhjTZEKCeBcg338KrQ8V0RbNvgPJZbge90+evj+bRDPC+
843IH8S5u9u8MfZutNsg+lvLQ+OIAasQeOOFTEFF6zuvPM0IaxSIq8dfk0pZHw+X
g1qmkeaEOWjdyD3BouBBOLeNa3G8+ejnftpkhjwzPM0p3O+ZPJ4K/2LBLx/D/BT9
FhObHRs4iv4nTT7leO2Lw06f42V7tMg6AnKdKzNZY0Fcvqg0Vs0JBUCvW73109Lc
2dsPmRrx5FANPl7BFmLggE5yO34FxdA/Vfys+DnXpVC9OTI9na4VvDcjEPT/JnCO
DryAshXE4FqmnXbrNIfdDJvMOxRT3hpQ7R5sB5bzCVfHWXCwmI10GisE701+JOp7
CMY9CxuF8pEEzRTUC3BKejY0gfNXEziaas26rv3Qwd5WcpYT7MGdx5QiOcVdx8SQ
D8lBSbUGGPhDzQU7DKQO4AEB8dselzeLyB/LNvtFnyLrsEQq03FoL//nqu6svwz/
nqYScZCT3MykSqy8bvkeHv+lAuxT6grMVqBPziuBn7mc8IZjaD9MYgoU1gS93xOn
pSpoEimv9EsCNGL7RVd//XvHvvxVagp2e2jRFrg7kXb/8EuQZtR8n0jIqeo77DIB
He2LeduRcaMIhsXu2nGbQyJ4P63GYYGmXYTYx3kyUpGzvgF9AhwOwQUVpcicpn4x
nkhuokmeas2rzYk7AQKt7kYgnT18I4PJ2+5/GaMEWIIN6bhHN4Jz+njHosp7cBhI
X35V9rC3nfDATDpWHLCYT2Irbp0GLUuaD1Z47hjb9BhowSBhAGQETh/T3TEjlLpC
YS3XqqLtOuDz8/jpqXca6Du3Iu5eksWNjnVt9LClYZqqrzT7FbW/pIPk3+vpRMkv
XMm05V//LmIJYLVh9CCJmqwlYAfoup+6BC/SAx77TY2kOgh5Ju81Un4M+HptggZL
zp5awpxFPzCKe4IWc6uoGYjq3Qo9jVzQ4hhVn0oE6Odeqx1qAeGi2UyDO7HYEmIv
jfwGNAJWkrjfQ3WnT/+HAKA0CDBhSOoyutrUB8kjuZbBtHtgqPKYHpBsqr3j9JS6
8OlOuj+y00+Y3mqiGj8Z7D+r3OtXSVniOe5Y+TT+u7DTTMsZJkw+TJoPklPTMyVU
ar7+b0zXj4sDlaIJL4PHz3iS0LOdbqSrjjj7O9AwLxcZr91chGmzrPOOTslYaADY
+3f/jS3JCDT9uaqTsmWS1rK21gBzwiuByHCWEc4WFyJ+UHLE3Nyu+dfn6ikJ9LGM
+VjRH8XxIdJL/lj/aMQCgjSeOOsCu/tNql5o4ZmAoKC3amzur3E6NzcaZi7caugr
GeY2w1p8LczCyqjAvPqSYEW/PuZo0Gk+YsIdpyuDG/UwWQ4YLpslFdn61Gn2talO
WYb58cuA+Fh9DBxpgxj2tYHRTvm+Lo0oUq7hYlnvaZqPyRpdtNbY3lU8W4ynEdG6
vyDekFN2JmIffyNw1quPSR04N0QLShDavietHKeAYWVIbSy9kuvUeV0ARF6NCM6N
8Bks8/smZSH/LYN4ZnTvgXyrA6xM8GhKKdk960E62qGUK1Ru7KVvLtH/zL0mZfMT
lgDqmr20B+D+cACfeNnEY57WZIV825H0DEbfqEq9ptlr0Z7G3agjSp7CQq0EPHW5
0aMm1kWekZ+sRCb1GfQ1Q7/6FpFW9Sp3hq4qOeaV78Fwar+piXEaZ6aREU1K9Zjv
UovB80IkO9SkQTVFOtnusu8wRjDMuzYD9wzJb4NUJww/vAzyxQYOLqZkNvzKB/VX
mBsuaxiWL1a8WQfaJ5g3HQUgcYZXjJiSC2sUkA1xRwF86SfEogn4MfympfTsHU2u
eylHfC6A5OqQ0wMY74+rYPquy/8niWK7Kx8m565nkrNFrE/YBAy3vNDwHJkO9c4Z
9uCin4lyE3znDTqphuSYKX4TfAFkKumUuB6fbuWr8Zs/jGyZmh8AETz8Bc5lLZXx
syoe2GXwasG/SwirjerHXa4oJf7GQCtEp4qloH/nbpqMr1s88Wgruvu1b//spTYg
Fjj6TvpFBURYZ7DnFN+TuD5uS1zftAEcCa/8ENRSEZdq+wOXcHuPnlizd2X0ZvhX
0mqj4yr2D/UGhMvX1C8XMUPluh+JdQu6xtg6lPia3eqo3lOo52yorFDxdYNsxx9c
+VHAK9i3ucV8JeGDzbGWL2vJy2w+JKFuYMOBpx7/rXloYYrh6xj/q46AgNq4fn2/
qd7XQlHZCpP1iF0IWIM4F3o3NtxH1pqFqsQffbaUxRTIZONqvCblT4D8cstENecM
7hHhkbxa/+qBOY2WnX81wN1BnLsoq/Fh351ksyYeBfHEbYCXEmzGPa6/sOyd79Cf
And/AaIp9bjEiPsNXJvjFzGpMiDvK+iIrZ6Ea9bYJDKrwzi6v99r2EalmvmSjDue
bBIsDw9KoCl1vmX4TvrKVredN2yFg1CENkaMSW/dl5ZEjSC4mA6DJRm4tDFkQbMD
CidY8kmjvUIfsGS5xQ5KUym2eG79eC4RITdH/4WksZsAIaems6SJ5S5FNyBGG/X4
J6rVmzAFgUY9ghXRN3XQ3nIfX+sXF/CYB9mO1Y33lBE0vpxa4n8x+d/QsP3lm+v0
2y8atTcc5JPnfxvS8RKxFr/ZPwzlIQVaSuvgOPWtd1yLQ/2A/djDS10wz//vgxds
9d8HVcmclgU1rGrcVqxDYtIyUvb6hfgEaOy8OWg3m0Tkd8Gl1GW12Ow+nERyo9hf
rfzVExAU6qHn8ckbTFKfQ3u36Laz4ZxZHyTI9cek4GL0dhvZ+PDAv8Us2fsRYOEL
hU7gLOFBKGrnajZAhcf/oJesfiddCUag3+cg625bCn116rm6ghTkzp3TKfpYryYn
njbK53k7f7uz+xrlSNgc2Eq/oZ6QEdI5Er5iGV8keeE8feptKgFEbUr/knv4A7v1
XrNCVL3krb9swi7mL0lIXa7tbgywTnGcznpNCcJ+kdrlvHDrL6hdnwysHaotFsEO
hmgtrh5Gclp74hU7iYQdUemf/Y+i9Zh3pUMcY2dsM0/5Yw0etCM3QZRnO2Nq7UH9
vtZzAN1QmhcinPteazUJB8APrCVOLkN15JEzJP1sw6zbOpmwgONJUSPtjD3LAdUb
u86N1x5Ay3qPOm49vAOmPKzWA3jCP7kiSQB8l4w/v0nWPbj6qfCBywcXRnNCEoIj
Ce0fRZT4J4ks6AAUF8Ren/USfQnuIP0dqAKW0K6QcZYzW2cHgX48EcJs67z413eS
htoOi5uE/r7ECkIx0Kq9EVrz/G1bWmdhe9FAFLabf3Oj6jI5gR+07W67d3L9mXTY
Wu3y4jychhxknnb90zqDpFv/ITBlg4SaWpQlNRTcOngvQ5ee7+zUdVZbZBgvTGlK
0PhCo5Bw40iUuE+BlUIACxdAUf6j5DsPx/APuxc0wZBrnA+1lhP6o1KSnd44Tp3o
in5hGTunithy6rDATsM9RmGmUH3s8l2ma+0FLYNeQHihrgYgP7Lb4XeC+9vPzePt
PEldY8/j21PBEq51E/zDzIDclrigUWwDfNrynlCYr0+ZlGf7tj78qMOvHgXrfQjb
X/bVXyCzVygaNyW+bu5XqFO61xjOEAfBih3BaABkmn9KjKl1mcV/X24kaHWJffvE
dftAL6wpu/g4pEJauiXaQNZIkLYkytxpm3jRSV9Ze4lntVVj/Q0w6KJFD47qONjT
Pg36gzf4ohToP8VFDjx40szMCOLYHHEdDzt6t8C5i0bi0h33h0ehnszaZWJg1qRP
AXoB2v4ciKj3y2/p6oFTQV3qAREsp3jPIF7B1i+Bu1AVY13uBxUBUvAMABMWzqTf
+iLhAP5ZIqk+Az/NF9BFknQ3S+Ld5YiYtyveEZn5mq5ulfdvMStHH0VP8ClWD8Ra
j0BY0HajnlqrsxFYCZJ7IBxEg3ekR9uuaQgY5rDhYByEL2MSbGHy0N6jPlAny+k1
GB08VrCjQWPMpivMUD/badCce/vm2tuoDJeaukmHfNYFz7RFRVllnnrMrWJrqlGQ
jdoObc8THi1xCY0RUYTun49/oHfkehU973G7dcCUxNBQXPmAX3BFTHTwR08HUUNi
vYpWPv2o5UXkb8A53as10DAm+M79lcurPrMgthSihnA2WimEZFIgSW0rxDz2NnVp
SMujoi2QAofdPAe98pzXL0mR8+tETRfF7eiYeFP9BySuMYQFWu+yo6Z+rL057/Az
FXEgVRHSlVEcTGYP96+08p3X11z/JyukyhiCh0jVA5NMkgJXPbNnm0M71xzojZ5B
HoGYaHVKURY1jEfaJ7RB3k/n9t54nAjzhdg+fpEl5sFBD7GzLTCK9B3UYxHMmtSo
dKJFRtt70MbSCmxOwpW10giSLY9o35nYKZK05B+tUMv1RGYb+i+dlFF4hyFK7FNK
1sbBpv6KYcxQleU8KbEOwmEHjP6tRxXpgNJew9cI4P6nyYH8TO3QcSDOUQ5A68XZ
QgyN/cWHi2MVsUEHVhATz+1exmNILALinUuUAnF1QIz3EvLzhW/8k2jFLa0sd64b
0oheyKaUdtQl1m69iLfgm3gafoewNVgC2TpEOv7WUJhs0Veai0BOzuJt7dB9Ly1V
PEsLDJXo29K8yfD+GCqMLTA314BH1SOyQnClYMhGpxvoQETQHubCDGOYgLakKX5M
YZ41fXDLRNUw1cGbpcZgHlpjm0oGzntKu4ixzt2NcJjPz4qKSxOG9drBZkUG21tY
EaxA2cNl/6pGdT7HIq0L+GcysG91MKfYWQPTxTx/3Daj+e5odvxcTmwmZtFsUeeP
6MROmPDA2Z9PK+6WMnX0kEXYU0CyKOsexTqM+RkAcTLEtcSkFkt+71xILiHBF/zZ
ZC4uck2zYuM/p/CPQ+SE/qltg2mkNeTqLb9UPRsRi9SZ13KRKwnO1ewwKowdYaik
S8PgIWoS+jXYuxYxmra4ABoad7x2bCBw2DGLvxTJXAZqzs/1Adj97Y6brfN7vJkk
meEIMtn++lau1IiEZVGqZTtyPdE8VMVS1t9He6g/4l/cJLD280Vud+Qs+Mxlvqf2
VONjjFCX5et/Tx7Bglcfw8bL80JWbY7DmygPTAiJudf7xS3b4FWWNhS3cRGkIiJa
eBKpGC+TNiaySgZBaLbG+CpGJbkN+0pIKJjlfgQyq66GosuvVvl2bwrs1iAQuGzh
mx9Aqm+xWvyjRPOPsl6vd/TvzDFw98lMukup2Vq0a3lgByZkfbeCBcgD1h1Os5CO
5vUKW1385e1Gnt5us2D9n53YoskMVPtc2Cq2fYkXUW0pKZ8rFYVz1s/eDOcHlhF8
c5grF19dLh+cbkPBXoHBQZnIIGeB+FXX1OMGEFslsCR/Lsz4sa0nak7NX0gpLgZl
7TA1DqjXnHkr69H3Fo4z4Tgy+ZRys9FDQKXPSxmI1yFXCXM3tEH5cfUIvjPvhvfW
eHjIrtAlZqkpTttQ3V5ni3IUaqhUsnPscbFdQMkuNXZt3tban8rCsCuJKFaYQ4SZ
p1oO+XJoePb6qWWi3GzwxNKBxKxCdtqNpX52DFAqV8dPH+eujdTuNOuT1pw++Kqq
9h5024ZCik6AlRy1epucJW9uQabgKbCoPBqDRW2tTpde5qoN7ZSPXF7QbO9jhDSD
XPKvlgfMB5w7b7c9/M1l8RIn93PnvoBUZfyjulAu/HP1yKf0ZccvrOVcs7D0m77s
sVHpjjjDcomuzjHpg5MQKN43Lwcvlf/C11glEX1wwBtrTeF5YCwOglY2I7zt8D1v
jkCKC7RijLMyty0+zJdkOvGcvVVxz3/Uo+EpBhrCsvsHDstd3Bz9Xph9kpNbywvS
tM0Xe7FT7aIuAKvHQjknjBDNxZ0z554r3ElIFN6rlun4qe+b+TEG8sL5dzRp8/nS
KElpFWLPgOxRaXIxUmO7o6i/DDYMMpmKrjTFPaY9tQ/vtrW7i9QOvW5eI9qKgsTV
2NcQMrQDiEWqpZrgNBc63vHzgfxWQe76wjl/Vbatiy7C/jg6o2hg37DfO88iL4Gw
9D3ssLVfHfut3ZTvrCrFQ+rA2iO3lrP4Q1eTMM2zdiSyad539VV2dFzyY5xNRvq0
1p+KR/jn/1KBuPEwOpGFkXL91iW8bDL8aytXXy/guJefINZ7SiOT56j7gWi9dUZq
UEdNy27wYCMqlTBNfNbkTXUrI383oNg6Cx806d0WsE7SWcj4wLE84YBu2SKZ3MUy
VA3PDyeFfvdvTuG162wDMLZi4v4CcLeeExeFh8HmiZu6QYE8Ek1lh5U+uD24GFEf
1QEUNj+sQYGIeX7Pwo2sFr1yKGr9fOxnVN2lfy1YsnJfNbjWO3Qv9llEP2nhYsNU
TSjOhx//wUDYIDcD26sqPuyU4X8dWp5Uh11t4/+EnMXFnXRaEgj1/3+q113zQLkp
K8dwd9WxFFyTpKXy+BFCZ3dQvVQGb20qS1rfpUTjT8F+MFk4/BYwY4C3fBOmh9Tf
5sI3io+2JpLNqk41vpm7Hr9WrLoVPKOPHPSw7++zWqll6QpJEP2fSxzb7CEPTtiY
50HYD2n0CinDaZ4sc2Tq4h3GcvPbOlOm9mGPxMQPgt6Ysf/4/YC+7DoB3O7gMNd0
1bl6lMcrUXg9aX69PIGVlezCGyzoyZl5jM5gtPxwJvV67unXiFth5Df4OOVXE8HE
6fBTbbWAYEf2ZwAgfXdOctxUuNzubCFTspqVk4Fgoz/dfR6obu/aNVOppYtFrN5i
rdn+hL3teMdlwRt8TvoZdDveUKqbyjmLrrWdRDy8vNbccZRdFyURbMGK4YbSzOgN
weEXcU6NNqvbC5rsUWuP09G43ygd0QpBDnzZhGyfMqdCeEBTqxyqxwiOI7yyD1/r
p8I2UVr7mC97iz8UYdVcSTowEwwHvQTQGEYM1KjNg7OFfxW9TLA+IY6JDh1gdn9J
BktqtpCxEs2xCrcdBsvOxSJftUqgEkZWiHkLFUT4BAZ55/uftnN/kqVq1ywoB2ke
T6pqxmwW9YMjIGcUHhS6UxRwgV9DFpM58J/L+M3YYJuteOuUlGsCPpkt5xfx1MXi
Bu0YflEBjJPfrP6f69gN83PmB/wBRKITslzxr/7PCGP9C+I4V1ccF8CD414jSUuL
pRfOuNaa2njCFax+AHG9SQxKlEkVVWdC+c054y9BKVka5Uw84JGoeaqsSS9g5P/9
Rn8yTYvhVJXvd7IMGHGXR0+8TEnA2Havlyc6mt2AxLO0xhrii6NIdsFFoT2nSC1/
ZPdadics5jnOpdwM/IvflmJsI3W4Z2lUJesnvoyRwyrttsqM1AwaEjaaZqkdwc9i
84860YhKrwszDBlCKjlMJ12oB9a7IcN0S0NpBPekRG++isOdRpfOVU8EcMBiFHUs
/rfonsDQwqzfhg3Dw96H9msVDcXa7LngH89cHWJT5CcNzV1M4niiZSKSchjHd4l9
qoKqIp1rTP5H4aYMriVQWukTIoqCHHoAG41BmdKJDJJYfBHKYwjfUWun5/cdHtTl
eAQFY2jtLkBCGukIaFzCdEjYQrWet2Nh3VG8r7gwJb1E3qpTyVUesOQU9Z9PmMJs
0ytAyiX5yhRIZD102xzGA34WJ7pWG+BGSGo5YkxzJtdriAq/WDpSyDz6NEgU0qVk
dZYXys6elHoDr/JYbUCRdWmx/shSZFYwJ4P+U115+VPyc48DsWVgnwrtLXz+Tc5d
7q5DZgaReMeHjsbduDUlyLS8aKN0R3VK9601sOB2rFIysW7Gx+Ys1VXnMqnv7G4m
sAf7L7SgoFHkGOy1wmL6xQx3zi4xMwMtEBELFL87dbJgJQ4Vo848iRyvge3yAZn5
c+Vp8Je2borXRUzl0vEgdR/RXTnUtDcPCHY6SmtWTU9P75nsfLTGU9Vn4/ZeMLfR
opHhuggauCELN8Bl/CWXjErEcFDkTm/AFSI8zOC1aYEq5hHBAPoDDrZD3FXKv4LR
bQ4/FjEZQXH4szh4BuEhRz4UWmZeHGW0eOv4f0B+ZZQnn08JBy56SfX+VhjqyWno
eoKHH/Mvgnx2IHKaqGaVtGy8bv8AfRNoLZ/mBSyCbxNxV5TvB2fUdSwmXXetiWhf
Q5HsTg43iVq+p2a9+Y8dQ5gR1DaIsuCoFBbWCdpOEPjhpAPmJ7GJ21irgcjtHW8n
Cux9tTrAszjg+sbvoY74rNyFMgWBgHc11XsblZFueeOvN64t8qb5zj58PLJVoErO
6yeyBg0Y/L0if97mfNFQFoDAGT0/SfmGm/taDQDp8p8NdQtd43P7lkGbVmP4C+Kd
s1/kKUGV5ZfvOp3tSCDIgpDSO68v1D8HZrxUCaC2Df86Siv/ycj/RtVOrBJPQRSd
yw/be/MYeaxpCdTl81eaYvabxNtXcw5aWasVn3bw5UH2yKUb3Tb/6yVCzZHxwmSa
8JkQkfSA51+KkDG8/B0OSDsUopOJpzcviGkhzHfHxz6Mwjk7Z72YvSY7iX3ry0xB
WOG3408qikFr/lfbS6teMdfQXHbnyRPMwhZk6iGD1GWekjGJyTrfGAdXGhzzTqDy
CXjJb1blsXrGVa7JLxmbtszRBM9ArD2TytxtySFZW91Si3b4Cm4w3qdMF+8ZQOoh
22Q5ZW36/QWCzEfiwv/VjdC00AOCyaN7yfWR4+ix0RS36BKw3M2cyQlUsllk/4Tv
HuJ3PepfA6ludYKB2oeTvRxTkXQodwbZsHetczKNqEmOATkuLbaHZO9GD7k581VM
BLxeLr+KCkpF9kcL/YiSsI7b5FctFO0Z3Roy8TTLx4elWGOAfBdWOccw09yAmC21
j8ubduqA7VU/k9mS4OoKPZ5kKfz40zFE1Kn0ocz+GokZXJfwIzRI54XRzm7rHUpH
c952PQRMl9DF0/kos5tJtmKG5stmBhk2Rl1wLVQby0thKRhQO5SPS5vJyGG4lLqN
Gf+Z9sMHJMDd1xhFK0LCxXDehl2TB3QlI1eFTQs8Nsl5X8No6jnuNAiUjN4nPnTH
X7tA+BSpEVVRyv/yqPq+vaDoxXAo+F6NbXbwbn2qnIevIOqwRE4boUh4z5/hQm28
FOTO+gyQzN506CWdtP3YR6bYrDGjKZwzH9byYeFxR+T03t4JA6wIhO1elxxSm+Q1
SnyZs3Zf06rpu92LGyY5ACdaWIOLijVTgHCe3byXZ9e7go+qcjMQcBczOh1EJ382
vg0iHvrh4GPPdhE5+SVgtwhftDly6DaChSdhHTQDE6Xx6ig4POJ44Qu+QpCJ5ySM
sH2FV9SVjl5+vMuGXXQCTPjbbYi514nzekRFqqWPvk0xtR1N1XJitUU7l3hgLO1X
0AvUmmHBxrgtQU/Xun1GyK5IvAnGB1o8/8MLw/Jm0oVZHgjciTZ56eG72zDFvZu2
pf4CR0s/DmCtGgsV28SuPr6a6onK9Ef8jbyc5zEz6Tbb5KCaOhJyU8Y+1bqPmPcm
YREsLZHn5OyEDqiIZ2RfK9E7Ec/bNdRF+AUeuYdL+nVmGGnaEK7VVqdXTc2RbPO6
gy/kBeS4AcbLJlVP5vQBhZ/VOjbJfXenwEhXqSt6yLlAZtIMYesbZNYJeeGHcyoW
UdafRpdQoZnrGxekOHmklcAWmeCj9IVd3kHUhqmH6zZgtbwpViAVyuvk5ci5P7tr
NnF7GAScoYxSlKgaIke6TigqLcYpibXGhLmYvrP1xT4DRQg9CvQucS1MQ+HspgXp
qhcNVd+o1gHIsQrGiSHHnaNL2ArChVeGy9wXypbpqatTmwcokFACRtlfL5i4krQF
Tm+wAP+zhioWA+9FLvcmoTe9qNX5L06RNeDYv0WPkVR6PAX1MB7XFUxIKa0BcYZ7
UFK7tRi9tc76zhjNBf3ZqyosxCdpXKD5Pyey6Eg6Kf3vYkk3RM3pjtKxSW1xzaNT
wOCDTkmAxB5kirVo9H4MkQm1vgiegPbUudmfELKVvtzqt7nCO65sbbCmtqDbxagj
+3/dCRdvxHs9QlAb4MUdLVp4+TMVdluxp90twIYFVgEva+t3sS/g3S42XEb/SoUl
hnpSpXdW1HFmQG3J22HKkWoFSIgazLsv5okUJvS9DPSc96T62c59eK0FssbMoGO7
eeBh08M5/WAD+BVPxW2bNdL6bYTIPmPvT2CAZ8X1ETKnjgeO5X4bTORZ3YBZ2i4p
liB2YnUq8ku/O1EiMKkUr6lZJ220KWhZZXQrh9qbpK8+mgIDveIIH7eCh805SAGL
+oHw3er4WD8QN7jTtZRdnWms1mnlHbKb7+k4QN9z7UjAFLj8CyZJBDcn6S62yR2J
zCy9uZlyPwj5MeOHTXIQWbszJ7OkCptN8VqQSvMMtatYilBJSwyFJzbXEWKXlXwE
o6kpYsdPN6ZWXn9EooMa0PlVrc/utxesX8XtmWooNY+5XW4S7JrZyWHruOiR1emN
4CtU15kJQlQi0S9rbC5xGGhNXGBfqpKbfp30kjEgtslCxVwo5E6RyACF8Wc3JqEX
bDxF6ocv+e0d8XMkU1v88JdIBTX89JM9rmK6VF1kd7ODrPStrHBmRG7hDk6SnB4X
h7U8D4vqycPqcSZSKFCF7LZsDkugBcklvHMFdcwmCu/2mAUxViEXW7+Hut123SVr
HTLh4ra3ywFZ4yOGfW2mOdjOGU1DGhk8oCgpAghMRt67ZMn2tO/TQDd/Us4BpIo1
z8SNuUSgRqqs72ndk+u+CrpgmRu4vp8vyghta8LlgiGrMfs/vjTvynENpPJMyJkk
sxnvOYxNpBnD85mJr1M27xBEniYZj9W3p+roJurJogWEPHI33JmkwXSbCXpg0JbP
r49E1EgJ/ozfypAwpMc/ZB089gF1XgsBogke4ObuqeKXKLE2WGyrVlCJrWcr6BhI
eyWppiA8+6sATlBBbZDBA0I/HM2VwWtr0iHWti/cLEbSknSCwWOLG7m44lFQdOBz
COBx3DaNMbZibVxFzmWYsD5CQ1hy+KUAiHjxK/xnD0OaFMlQZAcoPZmKe2NxqqmU
i/T5zyzSOowGjL9RhdhRE2SvdI1LVxFxJCswtgAJmu247ipfNh/2pHjMCiN40fLw
Alan7fduLoHLdMZ5zLRFyF2EGn+D0Z4Opb7L3EJRC7y3Nb4FkSdse3ajffY8LOA6
5zDIT8sWbnaXHhEbVlqu62NXnMlyc2U3k9W2SeGLz+nQVbdkgWDgPoBb+6yO/YwZ
FL9AEbknsjNAYZH4tcJ6ywz1MuFM1MnWII6T1y691Bg2BuV6UiQKzwdvt3zOH1h/
wmusLPoVg2vVRw9QLyvFu5keVHcH0sJXOR5bSOYITM7EbkKW7NqOELdUhMUATmoQ
bJI5jloHrL4PZ6k2yiG/L3kPy7z1a9J8gpVVs5Md6fqFXVnZ59jjAe9r8BytUJAY
CE0eG+oIMaNVlyXddM5cFc37OMasM3Bd8PLTDJX521Xml0n5/PnPFc0Z7Jw1e/lW
D+a8I2UvxBJJ666dFo/D+eDVENW2A7L3lI48xtiUmNQVRS1NxSsMsRHYU+d5vD/p
cbIFLuaHv33XGTOlTKKkL9TpLdJpt4LIF0ijUdkvC3WFUQeNrdZvEd2E/t4WXAkn
RQivGp2TKA5omjWh3Fm6T5luLYill84kMQsiuFbTOYle2j9XcZ5Iux2GHpGlBDZO
WY9kQj5fSs0UmLICYigylMUnnjelsvozSgdLijr93HFn7gU5XjSfszyN3S1pFMlU
QlKyvV19xDSmyg6I7an9n5dqNEHF1BXLBU6ojQc83G66bqkjNbJ3xVCtbinGxS82
ezReBKi9QP0X9wfbK8iMeMRKUI0qaYOVjdZfQrranq6UeeN2hjzsJCwk+ZWrBaVK
8YnmVwC5KMWrpYGIWmZu9Lpe0Cd62kyU0jfuUSktdLavzVSY4zBuxBG0ALMwttMw
bMM7yGQ92H5NGIKBrcot5hBPlgc7RQeZ92adCDX+lVkL7lrNuNrthsOgAe4FqKJj
s7BXtLV52ngl1H6bz6Jd8gJ6FhHKcPUH9i8GpmYcX7k2UySrhusL0HJZW+cGcxhh
uV0Wa7JnonLMw354IGi0+MZv7BHxqtYz8jqdgj8Vtl74UOeS7OFPgbwS+fHr50V5
Ktr66hJnOCrLyFObxQqzzIkwea1yOR4marURlOGCwNq7Mn9Qi+oLm0y4AVmCC38U
R8AUEwbCoWVO2+lmjdTxXvABa5CxLiUnNEGzth16VVYodWlztKaD7Kx0I4UQ2iif
oTAP/dAuA3oOtlpcEl5DgqbP9g2b6DvQY9GTinlHvoWxfqG3LyisKeQ3nv0H/MQS
z9aFa477ZFuHwjQlhxhojJ4vSnm+tz9StxCGsjLN+s9/T+26JctqMbPuhpLVYZ3X
jbR+vYn1ojO/Gf7LPWX4TWIiRxkwHvdlhFkNJTwgLqQ26FlO0EjCeG0HbOt19yz+
pETZ2qECWpkg9yDGHeixC60/moFlbe0tLd6RKMa5OmURRfryK2BWRW6M1962pIxT
sjuylA+it7o9zZlzeUoTJSYh5PvWJ3FJ+i2XIdm+5ZukOdx7i8/xEO93pbUVZlFO
w/hpq26zSlOH3F+lIYU36U+q6sKkDvwRwgjaeXyqP14+7MaHY8IHgot3YSuOZQ2B
ZM1+sT66KHOWJeJx1W6iYfZbBhiE3B5MLyXbLWKRibxOXp4Vr0okJ3VMcSqnvXYW
QFhYiJE2keVU5KVCJRLLnQ7w63kShAO1h/Hh3SxS+0ghSgsg+fGDPst/VWqMtl7f
icSpWZ5XPglap8CdEh8/3Z58J5+a57oAQ0RWr1BNN2ANYDHPoAIRmXmA1PbjM9Q6
Ye5fJR/w3mAkExyAO03db1fQlYxT0vpXE5+O/OczJp+ywD5wM/Q6Gmyzqk+KcNXn
XZwoP+OMxEYa3DKO0kZrG4BdlT/vbRn1WyuQm1JyDbABq+sB849SEm3ZD36mKQDF
pfsTu5wUVM5FFyFwTmFuiQiStkBR659h2j3YP/LgPG2y4SCog9GUVLUZKo/SIG0J
KQLMsKjaml0vN3+di5Uwor6nrBXBPFtuUI0/CJJ39BgCeMdAt8X64dlZTox9/2Ai
EZFKrdgadkiVvVKlcSBaSM8HOJKRnwOYB8i1ZcSTA0ZZImBdcBl2nZbu8bhuvr7y
mfMku1JeomhyScyIygtLVbczZl7+9NrxbKW7rh2dqLQXcifHhrLwjSb64PUyXEM9
Rx1IxapeCJyKZfgTH9Wctbq61DhKZsdXZx0qNubSJw2Mp+JhbqgamnEu75g/ZTmg
CYDLbR65s1O3ViJ86AtsDNkHrc6h4YtWNdzTbjYkLQSenpNKnsbA0Kk2YrUOcOLI
28P7518e3zs7xaN96nOocaP/aaL4F9GhYLdL8WrsQHNpS/lFGTHXQFunKEMwthFM
xt/4uqhA7zU2UuIoiTzLRiCExf1LjyHPicU6IISMd+PGcQaF8+o5aUqe8HBhFDW+
XRLFi7wGyArjFgBsergKJTOVqrdsV5rInFcWdvfSvodJdTaAqZIn06zjbiAPpvVk
SGCffBCEwWjF4Brczur5QMnjmowiLZ9Hy1I0PD74G+jbmeI3UgU/NFug5Av+Dcmz
kO56XcnsG3cW0toI8JscOd4xW5tG/yJV53F6yqTbz0obVOkCOSqguAT5Xe84iRgr
scr9Dq/z5Y6LqnySiItnZ5nZ2/IiNMf8ArWQpFfYYiczDRWeNpabawZrE8goxwtW
YBJqRveYbiTa/A1EjmkhDr0+oX7nArN47ahZxLNlSUGZLwmmGWegYK57e0Cw+dj0
yZcpNzNCeEuP27EAxwpY/eoykiOaMQANntorQ3fNhZAV7/+DVjY6Pv5UqhSUyotv
E85UzDsqxwSuFFGTf+c0hS3eiyQusqoVmWkRDyjnDMnqiGlo03l/ugOjDm0+3Xe2
xZ3YW7VDDhs3VWceTnPAkx+2XaJQVaa7xfHvLp83IR321cVGgBEpi9evtcCwzdzM
VcdyBFrc5XucU5A9VHXUi2zPwBhQMmPy0t/n/huYGD4GdQXJjLcgKSpNgQzLwrbA
8UbKkG3wzIS1MZyYQWgS4Mh5U2JNn3Kq0nLIweCtIgXXUZS3KG32Cq6iir6XtQJ6
ne/FBcWxPXz5vKmWm5yshxcQUvrKZBwVYFu9E1UkusJOL6PwDiQ9t76aNjOPDNHN
Urk0BgJW+/XvPGxv47xg0aooKyrKnLES74eDT3p6/B7WrG9/3UYiOJwldHdjQfcn
lHPQUIuBWrk3cfiI8WnsjW2t1p3Zsd07E5OtF+AlONDfNyVFtyImL+GKiF6qHkl/
eSsXDgQjBcIkj10wkmbBdrLs+RWnxYubYGE1fYjSz8iOkncyA3zsjdNMPXDa9IZU
/zb+7VrusdDCsXxp104mwMZHjR8T5V76gR95GxiCoQCEGK+JKdd8r0ZbBxLNakbf
QmoaOXiVMZbfpY/Wc4CkgVMQ1nwfE56P04VmlZhOuxwwDODnBl60GwQkrnC9ufba
r+DiL1vtl755ljdmuFFleY/Dg4TdxMKy/TjjcB7ACSTIjKEwhbOlkTy9HGc7Iapk
1IVxv5h8VllY1TE0KVaniVgMFTRYP2DEjY0up6tyj5YYZPGCQwylreXxMm9EpLTF
wlE5qq+FVLFtXQDaSTX8WVvt9gjbnCu9/WcPKQiiaQBlAGRJX6ZhOBe/x822Ys/Q
4m5Jwtmbqeo0J9Tb512AKt10UePtm5yIm53DSzrYGaR3tIVEKYOjPTs8jijS96tt
MgfAdNiKxSbmNQ9JKN0z7Xi9DONwpmx4WIuEF7655ObelUoM1LgLrNXzCpkd0J+u
NBEn4ZPD0erXu7tkAQkslejSBnTlbtfpoqtXUnVWmmEdexV/vq5EDq3EHIFQ3TaO
Guqfor7tDRfNk4kcLnwQGKEfbR96IHeVXE2hbijaJMyWdrWGlNG9GY7P6VTQZD1X
/DEiVCWUzTCw+hXge16ZYOW8HZerljGrLTJ/dD9eGm4SMyvLPFaRg8VyeZBU8M9l
vFBY4NqNPeyjrjudgWA5HmJc9nUs/oOmLY/dlm6Stda0/T3SMjWnALAlhW3RkT2W
SItUVxcDdHXuYWxEAOCvTBFYBHOdy+ptagF6OkxNdZf/MVuZBtkvI8UcG12uwssE
Kp9XoVlcQo7vAUJ20OsCI/w+sIFO+U0Ylu8Ny9O19WBMgS47VIzoGjv983R5dEl0
FnqLQcDbu8fnnnjN5jvjNfbfL6+SDqGUlUzx/aun7p3lDXlan5qBRCExHS0o9PX4
IROHcPOgKHKf8IimuOkP67N0pq+B+TxmMR8TtCateqPDosBmvjarlnXio9hmKsTz
0gsgThnYXbbvnh6JZ+K7ddqX+C8iNb254H6QR/e9mnrBboS2m2Uk2QOFcFeHzk5X
CKLbNHUHNykvRbRXO6FQxL0wdbKPLEKIziqCB7v9f1rriVwq3FzUtN79bdU2cWw+
tqgBiUg1hEMo+OVqvmX0iNZnw4pFkvwwPcqYFg2bmbhwumszwWVvpSHCge7izBkb
xjTgHhKpB4Or+ZqCD0zFvmTwq/hyoUJOQKl+aeAyFZvEDfm+fZZR72GLu1GUIMo3
R5rye4bz3B6kUGbXRTg8EjrKr/BuJIPWdQ6KZP0YGCYrWKFTGYhhvbBhLmA7gfbo
Drf3re6YM7HyxCwYojVMF6oYg4fWsG2oWTbxXL7FJUi1kQZMS5q+qqzCtMA8vFeS
Yt1kBkWr+K4j40VlParZmGsMQHBYOpqxJBPjF0YYXOfH025+aFaTaS+UvSnjIVoZ
d+BM8PjKy5ftTZs2vwUwRilGZMD8D7Rn+Styb5lge4M0tu7JOPB+usEHtNKRg2H9
1QoUo8SDdc+dYPj7LIozjw+fqIlRzUllV+3qJtW1Feemp82mO/ylrcDfcBMgwqnp
Q780HRntvpH5NaIAfo0qym0VrZ5b7wB8lkY7yvtVQHjZze0xH9qSkYXfyMMJPXY5
qJGmmiLXnP8YkYq8gSzNEh+FQLlO7wfq65hm+AX1TFpbF/p0GktBYbn57l+fZ91p
mIkACOypy1GgU0SKCmhsFifOs72at0CL73kAHlVG9gORzbr66wt2KBkCqR0ZCIRi
JfhX4IQSn1Db4d2pD5cGytY9WdiDFgcrN6bMt+4LPNAaC5LRLVKG1Mqq95t6lUgv
H8+thlx4+2LsvhvDyHj3wHr8ZPRYrn8H/Ww3gcKEx6YQ3QeugDx7/s44d0lhbnU3
PdXuJywCDuS39R1tijl8Jz8ajyJ538zJA1WwgeFTF3PhoH5RXWG0DK0aqstNxJ/U
4PefjM0SbqO8Sgq0ACN/nBJhdR5Y3CORm2REdKzC0l/dGWjl+4Gg0/OC1v4LW42t
qjBtG1JLOADf0hwXVOtfPEtIKcD6LlGoYx7f6yoN/okefseRhvviDi4E0v0eqzwa
zb5FCFQ0mEO2iYny3e3EIXASaJbcHmvfS58/PHyRX4P62yZvgkJEYtIQJpM8s0vT
R9d8/OTayEqR9oqNIphAmCx4B6A7xswOUxvXuXxppPdqHPFrKPne0RYyL3P6TXQ2
fNDGAPvMenHuscemfQwPKrN/uYvouO/LxQ32jJIiMFdXQBFGrL+8B6vPyWvKtug5
GzN6wgrgzn+yad+FQJqea9eQCl27RmOuUSTPhHsikssbZBdwdOKFRrTn3vzZRilX
o+ixPTc2Tt//5oTKoBIGaU9DNGjCPUSodTeycnagVdyhy64ou5Rcq4nx82DrSuGU
CAB3xtQ7WQdeJCe/+Hj82ElCta8+XrPp1ZxTGiO4SELlcdRbzahhkwF2Sna9YIc3
knLt4O+jA09zXMZTEV9sGGBDgaq7fQ/pOZ7UYaTQWdoABgHXizBEgm4jxOvmPKso
eNhkx7nRCjg1JgvqcEzKxUvPm9AbS0W/tRASOMD7bEZhSA9bTia0GyrNux7BlRE0
sLQ92cmq2Yl5iKlEiSqMEspfVvKWKuFo08ERnBFlQcRlKLPqzuEWmgJSlQg38I3s
oGn24cy9HabgresSUTcGGksGVHrrTROiUgGSI7d7gPNPv0PN9VN9t961AHqTlDEe
yg1P6ebi94/WDVzvKZVEnJW2XL+91CfIY7oR2KtGkyj9EibBWKQHRtf06F0NIYcN
/xk8FwVMeWFNshMq4V3V9RccekSvQjAHXFb5Vs6rpbtNeIkZdwwD5oWMxIE6Sak3
uGxG4MOk8SJXDEdE0HzmE69e6rzWHjx036Nc5aNVk8hMP5hc7EgRbaA4ztbVAHgT
R/55hZP7+RQxl4+DDODK3TMt0w+IoOZgeDA5XQlq2TBG7HFftxzZKGLnr1TKnV5U
HbVpN695y8pWAjJFRuX3e456H7ReDR2z6pEApab0/YfqNOtCEh+iQ5lCHoVl4PxW
Jm8VpRef59svjocv/0CP5BNPSvxMzzNYtYjfaHBoNf6MlAA0TGTBsUSM/x/2Tg8o
6kCgpxWpQ6AZzhRwtkP4HS1qOr66aRc0k6J1L+vpgnxdwuGafHzc2VbjIB41xyzN
JjH5fcTH7WaSWyggF4xfvXvuf3rDisan2J71vFZnOitOd0rc+qEmUACbZoiMBob6
gYkK2vAnLz0PYwoi2ZF7/KuUmVueahzm5VPuUkbhdHL01u6kRkGkFPOaUoZkPRZs
7syOFUW/SDzTATXkKainHSeY1rfTMV343RkpSulwY6vcnMW3BMVRjnoY5g2jHwbA
xkav9gmAsWQcSxPnJDeVIJaWozVTWBcj6/AisIZw3l5ddE2HoMwqjpkLzehwmAn+
aXrvIGXT2SKPnr802Gp3ozuSysHxxxV+dAV5THrq+x2ED73FLX74O/pAn/3vlaFy
Q3qF0dBKkdZtABaUoaj3ylbASPT7K7OLDIERB5SDd/OyCfwFclk+KWynYFleN8Qm
VuM3B1A4iSS7k95BrcyJNzPZnx3lAAx2lA5FfriBsyF3emgEB87/i7xuIqN8mei0
bhQxFL4OVnTAua9+HL0ruP1pUGJ3ZK34OL6xRU0HIlHsueU54w8/mNA3AqP9P1/M
bZ4zcLenIjRbPQ5DsfNksqDVFRbfQ1Emw+vznLd8jYYbT6KvYgcd9dW4kUugCRtj
TcBkdoyMOF0SSFSoySyVE6RWEBkq0P2KWBOW7GJULNLxnyTlICTn/oU5tcwD98B5
om3HEjZt3thQVnTteJMcbAINS1UVV0wsKpLdiu93+0wTT2PwCwtoo6tT8XvVtI8d
dVyEBwzdXtwv1ERNkcZManWknseI/Z1gPbHm7KJzu+3xOSjfYxK/m+eCGAWbtmgR
0SAEtFFQx+74YsYosfEhS5m2X2yTSgZX/TmTb8xPmsNlpdejrUUdiaXAwKzkkHBx
aD8O5hp2wFCRKd+LxlXMWuWdB2IhlAWrZBggtunReLy8fLedoHmV+siEsp52S8L6
FkEPjiQ9ZSHRPuImXY+2iClT5mc0MTCFgJ1pnw7CJwbgnzGCuVJQeVg1rZL45Vqk
BN5KMG9T58aPmXTGpBppZaLEDvNxUb+UFgICUl9z+AG+JfLU2gvB1emCLiKabMLA
zSEW/L30j9QAC/3cKNs3u/NCezqGv8dCwcxqqYaRAX6A2VxcV8QFeEWh7zf9MVaH
rmDW3qzmrWQbu6h5peR3T5+gBiATheFK+owhD4tAIFoH/UJLm1+UkOeqB34Mq1tO
QoCQI0ujE4FaKhnlk+YpexzpIHuGG1HUJjoKm7ky7pn0HQxdvDt0a4PgpDl/LXWO
OHtH40JNAMoFJUJiKh+8Nei7JA4t78OpZWpvvWZSGZATJjXPX4gTxTdBYsLLO4yG
NBr53TmDfGXuk7mRzuegMFyQpYeALAsTkSW7uowjHjQhP5NolsRQhTZSFDNVFWVN
ioUw4QDpElFaOc+75LE3rywf2nh/HPBNWnGRRzeEIl9n61P4K10PPJmZAhooK6Qh
5lh8qalpvWul+dO9PGjTSX4Qb3NsrdnL0ex06CiinuaDqLrOtzykR7OgdRLZVnWB
ymFpa4IqOFew8C4/KDiY6Cpq/urhybHYXmIdCRJhRYeTKaC+/XeJZWiruSyXImJq
WTTmtkToZxuxrvPp46mbirG720NLdZY/AiXtczFu1QkJdFPRB8Ikm97WyV8hnn6H
uiuUBgJiLSROFqmH44VwFwD2tRJR4WiO5QoirFYyd7gmr6xtpqn3vWEoa+++O3Bi
qV8jAE9IvjNwANk2kH53NqIp1cC/UIDszJMScJh1Q4/8U0rEfHCrTHpEQfOUlBoS
T0lzmyRN6TzXocWMA8jj9hC+XaeKGcL/CRZRssUw/MQj8elTb5AyihmajOrAV+lU
/51dqPelGnbNGgfq62s5hnHqLNIM7+49KXB6DsFetrR2fPSzMisjjNdpmNFb3rtA
Ff1sdCKcq+F1w42IQPxPEY2UIMD/1o6sECZ7woiKwKh2SKr41hLmrhP6NWeIt02L
l36wY+hcldehecBEc4VepDn1rrTRl0imrOSz+7OWJQoBrNREXCx3DIVxFyWELZ9Z
Joj72Y/IRV7uig60jzTk9RF3cSUJhFXr1mGtuWc1uz0Qn3Aj/Hr3i+DAEdpaQzrZ
Cm1KaPG2i+jhS4rvppIiRFVYiwXcU0O9yyEGPMUbavsghWz671t4QIJWjvV9bwoO
7pcIigtUYpYBi9x3m3JPbgCKIhhg500kh/g9B4lO8tud9WFPIB8Ka3BLMfokC9Z8
xW0G1E4+nWNfJuUqfrkV1Qvlb9LAA5SiNDQEsBvctm2C9mlP37dsj/imOF+R8ww4
1/15iptOs/JmTXzb77PIU0C41/o7gcjux60zex2kxOt0YQzemquARXSFvjFOuGnL
FsSonmQjWJ4IJrVjiIvck3huDi7qp9XzTeqZZaydM3p57eRmdMHqk2KEDj9xMTIH
Tmm38KRruzogrDoheYDBkjiFigp8INhsIBm7+2Q1Y6m2jGWTpjXnTTTgoQZnaXz+
WewNaXEw2/tTvezanF0ktesK3xm6BDHRCsYebxULJJuovx6e0BfApX9ejB6WqjXU
ULNpJRpeQgBud+ivfw0ICVWKKR/wmh3BAes56VNtOvWStvj0WDVqmwtlAgWfIdMz
w1YOPWzk13Lbnn6IbERJOERrwBm/rv8NmF6pxsBWCvpjB4zJyTLBmX32UgeexQAj
+k57bVfI9SItBBPCOyFWTPNnGhG9ruYqhrZd3YQDtXHHGH2L9Cwl6gp5cWVGYPlI
wYT3hrXcnTgYcNx+N11UPr6uz74gnx9hYkRRPrqoqgx3zZUpmg3gpJeg7kNA11WK
HCKQS1pm/vQCbGaFQ1tHjWjsWSA+d+IZO4cLTv2v6GsRsrvgdImeyyHVRXMHbzW3
8rZOVgLLnjQcuML1WEAHKSvNVE6VNbkyN61mym92P1yhsTza+XBsc29ufKUZdOUD
mDqkTtjTPteGq7U/D1isu/Xu4j3NpONmpIxkej34OBMBysgXEhfYCBXee2eyzc3b
pCIof3FRFUA3hH9tdTRLj2KkrCCfzPQio2Mjg9I8/8cm/imZ5cK/ApP0yc0B7/OY
ft4GrZKWFPIK/0jLFHHlLBLeRdLSAUBztAw3lAfJl+PGkWNQj/XGAj9OPjMDxWcZ
s2+7wGdTqEA3kBvknyHikvv7DTXW1pIVA0jVE1TqbzwaTRK3fNcrF9gxJLNd0qCr
hd1/8F+OPOLmo5UNvgvUjbZfru030QauHq/xO8bi3ajvr4LHhBpFzT3GQGePD5ZE
MgYothoHBM3RnnHJpnxJCOWAXDMR79nOIW+tuM2OKoNLqd9RNBPDy91kvoKHXE9J
Xi4hjqJSOh36DAIghXEDw7NvGrHR/Rdq350gds8h+zlwuWbaowD8p0capyV/j4lC
fBmOGxgS7+oa/vGDp31vCL+6DPTQn0j2OiOMbk6D/dWPASjmF9D7M37klRVzuK4e
2AIUIY30+muUuDTZi+cd1hp1ILANvp7wrQxPV9l8k/AjeV8o+OYUwNeQx6xKgBFs
hOSoRT1ty7dQM9IzrCKwAQ+DKBOUEcGL2gQZTWyonBzzKj0IXnH4EJ1HKgJdLn20
lxejR058c4Z8mRK51J+HKfWy+ScvrXIKU7Ha/BtJJnG5bhpishp1YpHbYiOoMjBc
uWyV1gDrjewrnrX0A39wseQtAgB9l9e12CrHYhmrQdZ2PNZsRlBbLD+XBJBlqZCM
vLAWO9LhxV+FweY354sPZCU6e0BdME4D8TejWxYUX1JGslHGT04GWQTD58re+BMC
RdrgvOIbQB6UyFShQNqsdRIursM+gqPwKBq2UzcETYJzh9kQbMW/N8fzjMzeO62h
mXIKkc6gj9xIa4Hhkae6U28DE6MDF0BZEj+I58h9ylDMwvjKHlsug9zRI0i2sffG
/ooi4+vfTuEuHdq4nsR0aQu0si+8tEbRcd5aK7mnpNe+aLxzBHHKb70VjRSFA0sq
nY0284+6i1QSNb+sbn0HFWIpGGtstRhq3v9SPt9JnPEkXNH5vn7FyyPhnAzJmpFs
87kHumof7kJehbhsN6tf/jKxZ1yOrsakqJ23+CuGTvoYjlfs8ocii84HP6t1XJwN
Tg+HFyssXOywI7Zq3OMKVjnaBYTKP7c1Ma+TDKDWNkG5zacPedpd5Q6y7WIqkeCn
vlL/6XME5G3CRKw9KYZRGyatrRgTtzqzSNdalffEjPVuPpCho7tGSZeZYiZV/NPf
92AmPcCq7G5uPsK9Ph/fF9KmLIXeyxbAzi3D9Icqw2kuWf8JxQphUKoyCUH7ItlC
MAWsW6VZw0YWgiyvyBK5ysNjOFkA+6KOpxlLgf+fzrx2YwaSOMxfTiahOFzNa50f
Mu5IW5KqDmst7ZvDSgB/1qLQWlsToSUl1WFGf7a2pH91eoQ07auNbW51k6LNQa6R
ESB6aVlI0JVuCbXBUKMvGxM/wccBSYcQhAnrxfqlmegxjiXa1W4FCEq9ITacoFWr
Q4eGVBhySlYGcEgPxnXM71f3/MwDMSlJJ+lnwwIvnea45SpOXmMofk0m/laowgjn
7gPIG7/kKuWqmt0RzQo9RWAu3qMfuZVVw+kIuJsRDohJvbKzT5MV8WCMz/CqRSuD
FebbVGZgn84GDNI3iHKCa7wG26tRi/uYdU4SqgYFFnv+y4nDp8ej94GJPtAiKvho
N7q9eTC/REyzX7yxPmKeU06t8QoCYkVrXc19bTqYK1LNypjrKdit3d/8j0FX897c
++ev6DeSKBYuea7BQDusLZp/9tozIfZ/eCI6OoEIuX8pjhmPXBR+DbanSpELG74o
PD5mr7oYCI75hwZP1JqSMxPKIESRichl75e/WvHp897pdW1QhrSPGJe1NYgUHA29
QVz3OqUTHpP0Uzg736L0mqkBWOjJW3hm1hk5lhCw6YZWbLDwvXTTqyX4FcVIlMNf
ip2jv2IofL/rcyGGF/SYWcMq2Q/Yrg62GfpoGBO/gWx/5IB5M3MivM197w0LjrKh
q4OgGL5mrCaGAmQQkK2r+0KNnWgL1ZQY8xBoQgqUowsnbsC7AIDSzYbbZ53hbs45
78LSpBpvSIBQd0etilJgrb3Ehb2Y2wVDA0FkLtF0iE4usFo4e+rkXMmtw4aDBGLV
BXp9dk3sCymdTqINbpeeTOOqYy54DNPt2oUqvtH7upqRNjTwPQtqA433ueVDAlaO
vWNOMQK+/D9ZE4TPvLmVN2nPuX4SPWlLbYVrUpNftA6C3KJvtfpq3FH/XgDSunqu
dnOXkvUeQ2S4SfIp5fbQBehl0v3VRcGaI2GP1Mgo/JRbBOTnycfgntpEyX49lWBp
SwDc8wtWu4k5oJ+KS3R/Q+krtvBmU9NFmi3fGcHrQLH+1OeLv2RsVUNrGDN9GbRC
/HG2F9EEjpG3NHixREciOQ5VZQmLVOUYUdOZYWL0tgyEkY/yYN7KLi+wFPkVqTmG
S/8TKlNF5UvSZ469eznXuKXJfzSy9Iqh5pW8rYi/Twq1NqBzuJc8I49V6cPSZdO4
26ZI9iKYazLVH++k1sI2taGEsXkOAsOmEdo/e46koOxssRHNY8GXj9S6VqKR407s
jQIEQOL1/g9hNjKfQkpFDBy2figl4SAg+gZiPISnysbv6+89O8bVGF1W+iEDStOg
rXe4HjT4+n+L/CfqAeZsccFtrjKByNJmqjj/T49xfRFP/33EvrNIcnXylqmk2rXX
sOJS60qlrLj5LxRccRqFB+XVlD/IxRoucPmzAIxHy1g9L8ERi0robQfYI9T6nSQq
UAheQUh2HZM9B4BQ7ktFxgq9HEgbJcAzN/oIHHYMOLi9/vhKmw/SL0ASgBToVs2P
AMzsXZk3TjqcwMoenVMXqzP3n+a7gThWtYx4bkDaaGj8kh7R/GkuPEjuQntohNWS
1ZwC6PJu20BZIeXqOxY+NSNkqTEeKd4l5sIkqX/VVfNyeVF5xPIQwTb5/Z65W7BP
6eLZv2JVnkzHLkUJbYm6j8XtvjrXYlDYA4Ubsnxyl0HXWcs2O/JGK9z5YXxITA7e
uAF9mS6iNn+dkizLDeRSVEq6/pHFFsVHGVlE6cMVltgmguPicL5S1337RY1+I+VP
pvMZYFpsKJZ/IfA6hnaklXrCDTjQqwDSMjCnukLv5BH+bTUwdJiBP/eLTiLcxooA
M0zeMoDguee1OlXOpqrOlRLj7+OsMSIFdk7JFqALwXD0Zpl2aIKxciTZJLGC/cjZ
6hNcTW1ZYyGUfiNd/ZA9O5TmC3cr0ksjGWtamjGGk/wAPH5vxlddZminwjY074MK
E3tXwgdWbJEMhXbnRKfGUmq51xhluE/ZRBxAESNXrGTGTSbiF4qH7uSm/N/xo99/
432kWicb4fLlvlXGOBI1hZquLddkBp/ahpuzi39QR9WuLm7oNozMN3f0AWUDX6NZ
L1ByQzyZYVQE4Vptb+BNspjQ9N1P6pA5jatOws52aqbtboRYGTqtaLwJuXzN+k8v
jxcjm1cupzDuQnBmMbPQmZgjDHNwia663ObTU7s+2Ll5gUg9nvBfYnMS0YhGREpO
ke2Q9xvOLyoJIwFUZtpCdGS9N6fCjoV1xtrY5YjTSCYnj33reZsRDb7aqZL26nNF
VXKYAdpb/XMArVrW0G5N0G0SKtFAVn7qy7oSfRt/FBUWiXRaJLHgZh2B65r2Cd8o
5auWYVSaxXhxKNUU5vpPsDy6PA2xzgVO9ATthFRkQg0l5c1oRQvtg4TVAH1/pdeJ
Pgr5UD0glWF3R9NHnBBOMz/SZfhkEXXA16ekK+hmxW80s/Hk3hRsRLjDXGVkNrXY
5R40saVu0GIsXiHw9Z2vkjOjPsCqM3ojWQ9Kf4wICApu3H+x6Q+lK4en/mdn0S43
nT64nqIdIcEwRMpMESw/TPRITaXFgsWdl8yxLzvhkvHrehjhD1+5AUJV7AyufCmy
oiQlMBgJAZOi1HbE9I//8htu9C7XXKstsoMP/LpHptLtaPat+WAEvD9Km4P7iwTU
2lcleDNbjgt/Jzst0uKMW2TXNH8LnQXI3w16JpQoNUL27Cgn+5IQUUj1iyRjc+Ye
ToR+uYyAkI+kvAJ2UksQKbLv3H4InKB6W6GgYq49fQxGv3BOxACDJAYwuIpiPnuv
OhXu8TQTYJJFrIohn/sVYyYjREQprBRND9u7WLA4WsVmfTDtFyiJPEWBWv3yl7CJ
bqIew7IyI1IvL2BuYd6aMg6EzW5dtGPvU1M6eBq/S6FoOqC0VrkNuJFjYAZenoj3
fDZfgKhPzKF0Bf136nwDAOp2cgSr3Rc9sSvbkq8/QAm9DHTzhVshsSVPjpdnty1Z
rBfQCumnJzJZS7sn6J9jYAwpe58gCVH00gIcJ6ivaqdGbPBiHJguCR+qtcmYZGYP
jmiv6kZtq+iqbrs6ysTBLCfjLsn+CMgmpelImmgSr+JuM0GNsOagenQ+co/wAgPj
Pv5nobLrp6pOEAhDMYT4mZYFj9IDtmqFxO5dnphMEkUM0EO+Ivqmc+WYMUO/1tqB
iLmSklMMatE/bSai1TkxmrZvPH/kMcQariHJY7P+iPOJInc9qeJAi3PTx4vC/gLJ
FIwbfWTNTlCw4/Ps07kvRezHU/5FFVeHDvx66zMGfnkGEqttTFdAtNcDYHsKFpQ9
TCiAV9Ww/J5ArMEcTc01O2qmUI/1QKV1LgnzCV/M3X/a6XHAVsznQpLMSjr5UdHk
i2dl8iB3dV931uYuhHaAbuTlgY/9eXYGulU+PXr0ja+73RdeuS9WFyWBqZ5aVOfb
0XSxaBmOWld8OtdgJHnF568YLdHmAFqfC7/AF6V+N+n+6Ep0Cyv8kEnaTsRsH9Zb
QV7LFkA5uS8CZ29bxynt+uS286JkBdnK7LSVBRxbd43pJO7XZYQDkAk/89xZH6Ff
5TItC/XwnrYrYaVXZunRkYGOLikqKQEZjtD7Fou3NvGW2v5W+nRaMKPyavANZ1LI
4fRR4yZcBVpRw3d2nTsMZLK47QpVTnx8KpT3z8Q5T8eAPZ+zlODJQuDO+JWENFfj
jri3lf7oom/LRvpto006uVgb/WJcN+LnGjh2/23ljDSr32ejhqee5UtPDasaa3pW
EfwggvrreWEeDu1rBuyqgEw19btWJfzKQQDb7OJgGAZzgcYq20AXOH78KerHT8bs
y2+EUzu+KlkkgPrHmPssd0RIMnZCm3R4LyB4LHWdDzFwV8s7Qv6DgyfkOS+PTarm
v7hWxL3TA0pdDHNTUkB09Dh/KNEKwunpcLPs8SuWX2LzVKIoODoCO/+aCuWmZA1/
AmKexkKX6ZWSzxFEfKpfHD7ueV89UmqQ6dzPkwa1I9ooLO5LLMcel5zFakqhGIyO
NVuJFuy3dewL27KvyoevOslxFGjfq3SgtZobbaCst2qU+g39BVaQGhj4aqsADBDa
yc92mW4wjUtd81za9jTQZoLibN+rVcxO52yUCR2ur8+oF4DAi8C9Gun5r2Mff0TP
Vkzmh53b8WyJmOssd6F+MX9i0A+Y0x026sYOs2KWRkSkI9glFYRL3CqlMXY9OP8O
cyg+6NLQSZnycyVIl82yP6ZbVnetFLeE9ey05tdlVcRw9z3OP+mEyhYxiRjzOgjH
Ww1e/X4hBfSuqpYiA2qc6t/CK9k3dBm7TI9EM1uMn7sIntjt+Sw/FQDtUUzUo2y1
SEvEQOxexj7IjXz7gpjfFh46PhmuOyBM0GbnJZFpNUP/6bNGmJWXbXNpV4dz6rA3
FmZSW6k+hyD0D/vffQh9GXzTFUdFmS7DjXZd+jvkfFPqePIAJCNcnIdsUpYOy3kx
VmM8YOeRD8JAWweuazs6O2QpsDd6oVEXbAYLH8WY/evYpH2eXYBwFw3w7MoXtXA2
wT397lDWgKrj276UYQmWRHxQxiakZCuN8DlIR43nA/fBk7zD6NsgoMcA/Sy/GJ9z
vmRK3d6YcLJ9yRCffW/qp+6g0X+OE7GqQNjpd3UhJLEdf3vUiQZEc8/opF4fNAlP
z64slYqLFFAnPxYE1wzHn8GnHS4V+MoVQaAqwGeJfDVxCW++BO+O7sa7C/UUk2xx
XJlYd2hfNm3xxviXxE5lVB9EOqui2LTlWGcfVL6ewaVuVnDRjoPhAKN/KEGhTsUM
8i3cKuyByz2XbMCBCaIh7MvjR5RY4KxatyKeOiGZteX20tdkCKRnB3v19mqzdntD
kYC3t/T16QEvzcVY5RDr0wJl0XdafJW2mZy3l5TuLW5KC1wxqyQXsUxkPyDWsSNR
M3ziBg4JuTqosR+WKbaTPXSIF+aiq7uMd5W2iTB2GAVriJVNMNcizmoSVABSfFYI
JE6bEPKILH9Rn7/uJT1mWn0Qk5t4oLnnplfF1v7sItQ3y1otE1qP+9THz/eWyTDM
Xc8MjLX9IiLrm38v9Xy4ahCGiKdGMuDi8BikqhAlRx0WYawuHyS8o7U+FRtRxToR
UL6hD53o/3PbC41LDmoMp31d6LmDLMvxrw2dVqNE7UYGpR+rE8xhY42V4Fia8mpz
qmezfPfCdWTopy6s/Aa8HYpx9lEQjG6gurO6vM53UtkjFkZpqNFOOvgY9uPEwaBK
rZ8N78CZj+MXVPYXi16CDjHQX1FVnbHGjV/kPQ4dpMwZb+dwy++W5FtXGE5d9aoa
ZuFwoSGAnPl9DhSupZJpA5bf2svfse0aHbJWvAoP33KmnQtj0+7FP+y6ERSbQF1m
aQHrNe/Rnae0TyEDX4AyxtDdlhx+NVjE+mqae4UlgEFnlyv3OXQZ6n+XsrAr6kaR
bfFq2rZwZAnzDTUDB4mVdc9PaDYG1vQSt+XNI5ubMkFLp9Ztct8uLnsaVrNSp86E
gAs0sQyIOV51LG5uQvvq8kRjP1wJfSk8MaqAm+Uj3UXOdK8lrHiNoxZ4F1s1ZXh4
ftIjAMMoiiuNNegZw44j82lZeEafRW/hDWRQeC/LADvBU12jlorzRTCSUbwVEvAa
YL1pfaR2QM8G3ioKrn4PFd0+kgc2iwyg/6zatZsqUissZeWRTvx9h8ZSLZMiUy5h
QOt7PDb1wBP63WOecVpC3SKoceskO9yAx+YinTf8XF6/3+9OvIsOKq77r6NYawpe
y/FOZFg8yJeE/9F46P1ARhcBfBIBFWVYeef6poYM+4QbZtyBQg34G84hvzdaQVWF
T48ogrfnpOnGbAdnIG0UyTf9wTql6yf9SOdpFTfiB4auvmGsMTj7pHskIWaAM1Oj
h65IP7qQM6dlzlPnquprBDOb3Bsn2NxIZKtXQ8Yn/OJqnTPQNDfABlQ5WCm6B54V
oyUv9lokia4l/FNVyaPhhvAnRbvFlMq+Z31jLZMgY+94RXnq3MLntoZtvVJZ9LTR
pbCyhDsQnFZbhQ0DRy6W6rwtiEWxIpHsQTF5yxrjQRNiwPCvrQ4OcvVmmJVUKqAH
XLjU/7Uj+u0eLYDnPF0V5t4PBl8750F9ITOitVBcgUspZTWdPj7iaqA8GKcYcD8j
yMVN+Ef4p1IL6VxfhTTk2hxL9kL+5moXpDnY7rHt++S3ynlWAA4xlFE9AJA3KH3U
8mZJDBp4ObRKrKKZtuHZYLJNVRCSzlq4MnKlW4VdGYewHPLLsVE56E9RN4ey6Ha/
H/Xg4avfY+63nI7uMoFDZs9eN57J7cNOzyJmK2urzlPY92oVLASYAzuKIh3HQv2r
Wx5pmbs2KaZwpBMb+N28ft/bgY34R5qIXLzG0TsC//C7tU3DKCZe7o8b28fZjPqL
A/aW60+TGPjLhuGghqoTPvTO3WYlEOYIk/NDRcr5XgVdyzX+FctDLZL5p0uMRZ1P
oL6IPwGbYAL/2gMZX609BUH4+8eVHhRfj/t2bfAMkNZT6QwGQFW4p33mhXL3/KVr
b3PsSCKNSjh0MK0r9HRXcVCPRt8fUfCzZqWSgZ8dvDuiI2Aq0EPtnp+Gn2zl581X
6G7U/U1Czx3yQOuXTM5/BcmqQDZv3i3DP6uTQKGZvMMG6e7Yr5doRnmBEYvs1RQs
q6EZvuzW1689OJXprXOLo+RCL7yjf5QmTJOZfwAJAtaI0K8VlFrD1kYWSVV6G3aH
ffYGWCbctPR5JorXeL7fRX4fzUDsb7QCnYUBrNCpVMsD9HOkeeVkN4KZAqGcz9xf
JGhDH+bQ3tjOAackkyv64wN8rhbFx1s50TOUjE6X3QhMaMZZBdEQh403WpdmOXeX
x1AlQRcjdUZHH6Iu5EJD/ZA611oxpgYIEibrtduE5jmZxiq9tdjZQjy1b6uynsWU
WXpDjPzQjSUkZMbkmdeDYNAsgDKJI/ailp2Gs2WZA6JSPp0FRDEKl4ZZqdrZoxpH
eizkyR/e4eJSTxFQJn86fWhrW41cvbOfsprsdmau7Ms6hyystQ7ocaBCsnc0qBD5
g5c6w/yVFpvSlKABG0mmtDqMPTQYwBMvi3CwM/TjbmqpfyKLR7ztUFM4GFFbgCEc
p3J3mVgt5Fhz59X2GMinKZUnBGRjeyjnhQcGeow4YFOMG5W3P4LIX6i2AepZ+WqY
lCqIzW9mj0NRERUFJcofnAxMFXU+4CepoAOUMPptJLVHomjKj0j9NVodMtK4Xl4c
55iuUlAutNNBSn7VbEFSIfcuCwMzuJGX+2annWt/0InA+Gg6BoThy1Z+m8Qusz8D
B3XGekUfUDV4qYYDYiFVN8NwYmxdyur+tfeEIoILIgvsmcsm+WS5UOsHA8ER1VEb
FwklgGLaXLGRUKmr2SvUmXV2m0lGfToHM9SKfJ5IUWqD/3p6tz5pubcTUwV/k3+v
7N9pp1eTTvKt5xLLvga44S4SSBD4EmDBumK5LT+w6cTSf73gMZ0LAq6Ra5f3pIIT
5xphlqhOWVFlP7pTGXj5+B5a3uiFd1PGDXCo8pT5HBWDc+NDqK1Wsm2/Nuem5A7o
WdJs1Dpu6MVyDPeD6/gyBTUX5Smw6aA/NIX2FiqQ4HgNKbwEaade+sIfGS2ki+gX
htkRojy3rV05DbAdoHTaS43+0XwS/m1Z2aWA4xVmClDjB3ZGWNIEWxCKdeJ5rx3Q
MXvxdsAgFUz/WiiblzOfxs482daTDSBNvHrA040FTkv8Gzr/JFsGzqxShhLWRx32
KnHTtS8oCAFYN/UXXYGxd/ZmAuVZlOowt/QuINj23uP0oOA5QtQyiFm8Pc4/iJq3
ml/TKk8YDZ9I5Cpi8AE03tePoq/Wv8vtC020Mvs09lTnbzQqDYMiMYya/pDILdZh
u2cZXuAyOko3GOQRgime7I0tIgG4RlAQPGmkw7EGepoxr6mzfZ11awgPzwGyp19N
gs1wg6BbnfHlOfsauXeCL3tuqTr0v3KlLz7OnDETjYdnGIjyrjoS+yuDxpN3eIg7
9usPDh05S8FI5wpQYuwq1pZb9UUyMyTXkPIaskysfUW3K4YCkn6ofss7X/kX2RJZ
8M4nqPN7WPdOYOpT7y3qoTWVRVrbZS//YVZ1JLmZRqorWf+gMFmfMT52LJkD0+h6
u6DVR/+Sg+k38zjYBDDbooUIJ9QV+RoT3dH6VU1NkMPnn3DNWVR+2jGhUMTyBzom
n+5m+5bGgJIi39oD/zdjD1wPjI26CpABC5UVhkyVW99bw7ZkRnmu7gdRkRU7TOCK
lZGR8B5KPz29SV2NsD86HUxGCYrflydtIlKBZXZs8kSamBEsASH8YMznP2ghL6q7
IB8tfPgAAtdGClE4pkM29GYFUKTCn4J7hAwyQc5d1MTjrB5JIlkVvTSd6Bz9hcdk
UFbs/D99imR6EdJgEDk6DKWRMi/MP0VW0RK149dM4pbdrZBJGZOB2IU/Jgn0xeTZ
RNodAJ1sV9oKO6aGGI7eJZxjYHVermB3NyTFA2abiVf+pDxpKtiRgZ/Bd0zRU2rd
gYGxxVwV0HrUnAd0vowNIj2KIq8sx9nT4Hsrs0K/UqsMgg6tFGGUh58QywslYLGV
exlKdsvxVQuWzOqrlLrA35Q6Oaizi+Q1tL38nM+DsvQ/5loNsF3ST857EXJAz4sF
YU1nqlnmptKvSiiG3HSKtFnPQpzNFvCt0v/d2jFUDsx9QIPzkKwRbXDle7hTSzyD
HcJdpsiMqBUJ6w1jrW77sC+GCrZaE9043u63dl3SXVJpOCMJ+H+FMa+nAipb2uuf
mbUhSGYkJjB+l3NVcV7WBpiCNo4VJL3mYEi6oRXrlRgCsnm8vo+bus/KD43Rc4cS
l1cNYLS0y2W5cHRtitFkK2+ebr2Num02CgPkhbisik4Ae4846Sfmos9voxEcTZ0G
PIuRqauPuZV5XdanwnwXgB4ykMf9d1vzvq2tYYrPaUxQcz75UKiTRCsCHIi0O+hw
hSRzNYgf/ObvO+U65nRotN6UCbinLd88Zujo/iSQma4GRcZa1x1OGwaNuQVOdQju
vd03RB4eoBRcnAoE0ojhWLchW3v5pXUNWNB2su9N2pKnqpF+zCH37y2Zh77ww6+F
am6u17wxQxHFDZRiPvrxjB4oWfrQiskmkmZCcA9gRIZXdSewLoHLmiY2dG1zxoNN
whT5mvYwmUq/EVub3WnKf/BMyWFUAeTNUJ7OzfeaeV7qKTunLXBNFLn2mz8cOwAt
5ks2dozdyh5jrj6ykHhdZuWCdKFg4d9zwp0Ijf3MEikhcZsiBdJ5fzeVTXB43H8e
OtZC5nHJ9N3gC4H2Kq7VRXnuhuG8t2e5GemdLIuKkmnsaAEbBxSc92hjhHFPBR7o
hcDTmriQHyGUu0U3nxVxXgeD6YQCw5XuzAAvWJ/oc/CvBWPN/8OYZXnnEjTRzu+w
AXP+4Foawz2mgLEVAklcILRAzYCHwNGy9TdfbvqCxqwGp6c4Gya2gnt6w6GUE6lc
DiL23uKjlhxr9yFvqwcc3bAHs8CHtnAOHqF+u7duO5i6RlUsMTUPqjUWMlwX4uMC
xa8qGafiuCEZzY3Y64ed8BXuxGLLjxQN37I1FALR70ivvVPVPNEY4vr1/RdQjuCG
QDFaRdwam9ELwU1hpC3+fiV6Eu7LXfIgCh2b0uC7OGlnrsv3QNSE9P9BzjKwi3LN
5WJRuvALybQc6OAV66YxELvAXD4ljX5LGJDaMHNxbAk2ihNDga9o6IjahQmDZOKa
tYuw7c1FIyWZpOgI1y96PgBoJy2O3/6+Gdz6ti8PFJbxBvis2Vk+X0wkSshRvbMJ
Pkc4dpXu9KB457dYOoAtkSLgHl+cj7usXRAfMqOktuSmqPfl3MC1B3+7I8kUQwqn
KImiGQOS4zE4/GNaS/bzyRo9ZvhMwXfzPdExekp89huAQS8Vexz5dkRH9ksuzOq1
Py9TK0YfqaGokoTUk9Kl639kb8BxgmAtr3pi/ASqgsCxFGQvDRT71+lkBBSUjp6o
njf3HIvEZdaFecsPYq2IbxWNtVlFz0YeSd4l2QJh4Hd25HFIFotcK8DtIV4W+fvJ
c9vNWSUyNZqt6BURVyJx35uB+d3DDz0A/0zy2uWbSMi9pALNNsCMMR5QdtIDiVMc
B5RFEUFo35K0PMk7gx7Yb3F+pXFUIHUKuljt8FAWyehG0Xl7zdPoYvugozDHu732
SeINmhpu6hdVY07wIXDLRBbo+MxN/ClHkAEI1BvkMZUf+NfJPa31PCGx/jRY57Nz
uWCXIMyZAqsYv8hcvtCdip7PWx8wSiZSIaS3pIoAWVp8Xf/YyZrDqFimo1m+FQEA
4DuK62GLMsg9p9QcipIOjw2fMaMCK4PB8P+bj04brkq6cD/meX9huOC7BItCURSS
ZUojhLEarNHeobHnMFTYJkLQx0kLWTjK0ltI2uv8TExlf9DSAxxrnHAqMkqDmfQO
ODTNK/LAmp9Ip1boXIcFgGu/5H+dGTq2o4BkGVqy0URZxrxTW3/SJuBKiaW0sZhw
6m6gyUjit9Y9qENS+9jSpYjNHsmpHTipnXV28mAbjTGzbkFb469EPYEgD+62c5Lb
2iUTQdkSTtFs8/25umVcGUrCrQCe+kJpt9hsBdwhj7RvRkwNkQF0QorRS6tV8hk+
Yc408NWYPmM34yzm5h25+6XsRLgtYsa8bYSiZ2lCv4tHvojU0LX7g5U92Y1fwmXK
vpEsB0Xfvy2UpMuQqTrIbxaBMC141urokAawJ9rStg4KjNXDkzUI8641Kle5em8/
6Qu9lhfvcKWQxUNO8HFF9YvbHnGTWspQWMZ7AwZGjrykRPi1KMiWWYgod21vRH+R
m2hEp9gduDFIET+tcyKaA93TYAKjLGD7ibPtweXR8EpqUfhP/p7bQPV46KWxWdpy
xLRA+gpjZ6yn0ijs/yiG9g5H1be7tRcchmfQkAPEuGJ2IAn0oql2J4kMGMnVza8+
fF8KJO/LExZNk6CCyh6T5HAmsyIVIu8y2T91jVI+QAydyd4B2ex7Oj9P36vSMMhe
ewMT8ADumC3XAnXYOZjvhUOoW1KIqkZkwFzWFkUFkJm2CDoEyq27bffrIPhvVp7H
eqFane4c8GkwUabgC3QmgFaO57sF7bZixRg9iQIIu55QfjfXfX5YSb92yDG2ZHnB
Q5KRWCN/sr7zdUiThB6kpYjvxLN2wFuK/VCQPqQ0XkoHCziEkH6eiO9Sa1aAa2hj
/tnTCuD3En38hrest3eZPSW4MOxH6nX/0idcanhrYqLHUne+dZB3XXUizs3OoEJa
zEi1zGaG+uNDhBQNyleSJ9KpaD8Vv78gL8oHzVHF3pEOSGgAdHESyBfxm4PIawqg
ooNjoCpFbh0KwjvVP5lmVh+JtHa6JMUycyjFHAMEwLiX0LT580flcE3FEQ9y+dKf
dqeuup0qbkZDGDUfMNtjx3GtNVAPO3PhCIwbLr7BkgDKeTKjfGGtI4K92oAXNgaI
MrKG7/UUk9OC/EVwBvR6gQesTkDS2kG2UItixRg7mwajHBFIROamM3DNPG7ckBn3
ugxWc7w9V7HEDcI+L6q59/UcyfiDxqjHHIu+Ijrr7zB00YOTTSiVGtAzjkoZYFpr
v2dptPkN9iKSY6Lwf2U8suuSxQiEc20uySZ8os5dFE9sF+3+Tr0wJEPm3kiwzrMv
uKNfus1wIsIWPczcP0yuPCSA7eH6RdXQuBnNJWTHwOzEBnhTOqQL8cpPwDmVFUUm
hW19ZYVKHEhu1TqnBGYyhGaHA9N1O6G4clZ9WE1Rh7ujfDLTEMaLFSps4qJxh4ZR
DVboPWuUS9T8mE4L/31t7IkdLigxCX0Vu2lwVTjHNoum0FAFbXk90YnOC+DZ7Gwn
44VRAS7nCDTqzpiubnL37ijNPEYJyKqhSb4nQPPF9oQE+ubXkkNXbhjPzQWlirza
SoZEV4eJ/wJEGpfcnIbrzXrfkhzh5ZdTU+RjWLe9H5yG+kLkSB6wBAHsYGkgkjFo
IabZkz6FSlq2l30tmAnNbNzJFvesBXYOx/YhSv6F0IO2T9XqAY9OWDSWOn9PI0iU
KjZoSfdRipP0jnFUzn1vmOHElUAEOXcWvlAyOEY6KO1v5rerzfjdg3U4T56tvG3A
n5ysoR0e4HlrSzgPwsMO95s7iq8mSMcB1VEz7cpkWG1ikF6RkHgnkPCfxL7dWPag
Qlpi20bpgI9t1bbe4/nqZwKIyiIuzQiecqrYnOYjh/lmutiVls5ZeVjhu9t42qSE
ti2Ulw8pVudfxSTU7Pa14JjmWiiuMKA2175nhn/MCp5arE6x+rH4yLAEyY9a/szH
WDAuT0bAe9ME4GJPFlONxmrGOavyn4ZPm2IeOiXQEGBg1HPfBySipcC5xS5bSBau
PC2gcqBdjSkxYSs3j+wBOQ+a2F4HJS9ImMh4Ei1Nj5RoL9avb7NtI3MIA3cOAftC
vRd96fkEhweu0TDk1SahH4PEBEzAnvq4AE00SFvkyfq6JoD2tzgr/9bumo0Xwk3l
3hR9Zjeiya9u7f9U/4w8Cjt5uXCd+pSE0Sgg87qyMXO2N+4NaSqRiXu8CfYJXqtb
zko/PlbK82lEA424thqni8QxyYWoa1+gn57PCi/wUgXD9PcHX9ZGHutaTt4wOv5C
FO8ONUPrTDwsOANLQqJpVVLsJ0qzIPDGDsJzsFbj+2uBPaAhGnCApA+r6JQRg3y3
j/mj3Uf7hHR3b1mstSZLcuKfkVqzfDSWmdS/66BRmG6Wzn/jvnthxiXGmTt9diaK
mtx8X3nQNq/amLd+GdyQCO4GnqVtDTc/+A368QQUHevPcku1/VBm9sf8DbD5gtEE
WEC3QMS00Sb8QHFlzcUviBOd4ipRVkXuqjFLvZxiAQAE5qd96598/JUIrkqaRf0a
hBzt665uQAeznmmXuHfaKRqpfgNqBkI8UOlFWUQt6K97CbhWn+ehfbuP9kOt7F3y
twWrvC6H46chpFhQkWN9uQhSHgLtGnefSdBJh1igvzcE33VPwyTT8M4+DOiwo8kj
XhcgyIveOM9BCPW1yrwdz/9nFErpEy98kUi/Jmudt+KdykHbCqaUScPl+C3PRYiz
Mj/BvPruWEQuYaXsUlQtFKOB4NKMYaQKP8gEwRsnFUytOk6N3gkPZvOv1USTS0q0
tsnLgImfhiXx916AZeD2HMywonXBxjsl1xCssmQH5I0FIvvtM2KVVEjZb0ECidjm
uGt/DdDjg8DdcvYEw/OmZlbud4MF/m7iYJoX9KY5nakf5M1YHgdJIOCrBltHAmJI
RuHZQRznemA2GPhL4mqvVyhuCuLcuE3oj1JHItZQQTyCWwnqd9v2I1KtReb9N3V+
Yih6dyvJnDj77nIMdYwHiKvxToNtiHDgG1c2DAKLdx1FHN+9rL08CQKiA2cPOP2d
m1AquNS+uXCHd7MfpHo6/KyG22BCDyXTxNU2NgmbAFjxrQQxiXP67vDfHImtZDNR
82LmsyjOtnfmN8sUesjyBpE1pGNP2o9tAKtR2BdvzNJCehs19lSh5eg6OOMnmpk7
r00lInJbxLMrrqoY51Ivjpdxe9vtYeQFbso5Ql7zkql82hkbBGTfenrXq1azDqJf
s+Av32NQxdK4aBXv/3gocFn8Ikqqeg/QGK5rWwr/uvAyJe7bt6XEThh4h7I+5Rjb
NktqQk0UyDvMtvnUQsfJLW8aVVZXOs2LREk8WJ43VrQt07my8vOT62fzt5r+ZASp
DNCGvaMc1DVnG2hXbVHVO2+uYuR8s8b1HcNqlcyfeLYvrxE9e/fsV2gc0PK+XK9y
oypCYTAWDycQHlYAbYiJrQSTOs4glyO0q4G7SmKKssFLIuZbQgmQE/ORb4IT07C2
EB0BYpUVwOSVeO2jPfYf9QDJNgq4rmyuRMmyT1AOEbke7Fm/9kArGugbdBw1cL92
ezOvkAz21aY2v72RZhWfrs+bZjqDrZUVRbVmr1KuXdrCDmS/hGmCFaqTQGIpbKh5
oJkqWA29JNfXQaK1bagt6nAZtQ6ojAgFTeAuHuV3rl5zsDlEMM5niT2CYi7ao6HE
wH3x8jAnd/tCrdcLLqcuUNxnndV2ccghBuIwoxKNPxWmKFDyYlnHZtaX2xg6M3Ka
oADEh319ync7wiFmjWwBBX6cK5Poo4XWYqtkQZVO8fCh6U8Fb4txiX+xOR5WnJDL
D9bZVRzv558lUpnFRTYCx2T0OuHMBrz8Ch2Yx0SNofnCRweKvNPvUYXKZx0A9ko8
dHFDt79IJdsqnTsOCcC9DTzjBBcre8qePipkVkotZ/K6mqmp26DN0XEFUvBLf5pS
8SijGCjfuh96T/sJLzDZdpb8I2sfQDXLUK0oX4+zO89Cspr9x+1u412dLX88Zz8H
/C/2oq57V+TBUPkhjp+0qlyi/0T/1W4JxJjNNadSsK42h4dVLIBpiBdodo0H9rru
OA2NmPsyWSLAdaxWpOJPRHRAQ3o4cQAtRBlWifbDqMeBY8pBfpCbrFcpY6P56df+
eR5S4ws3wHnZqqaVv7XdWeZHxvikp0yE1nZe8tSaLTJ3BJg54j47bUiuGFYeb0Xq
A5Y7xEcsv/Xbnrv/8zCisCO5ku8YNcIgz3E5RJnW2T1YN7knORPA/Yf5757rLM9Z
lwyw8rIm+Et6K3XpNPXjOZS8sbrIUu+sSu8bVLZOEsMstgCCTtuPDqofl3vvJKUG
43fWhWJoTWc/ldmnNL1+gyOOmslmRntIft4cnzfm4UaPgjC5BxDFH3vLmRcCUoaw
vOSVl/UtquqtOpLMFvMZ5O76QAnjF0zytIqGbPSt8lA0jeK027/7kHCusi8qk2hr
EzrIdTB/BFDmcMpt3Zla/+nXwkMulaJ/Iw/Mt2NOu93gv+ypQhNqRTP5NEd/Xmgr
mT4QkaZ8qOjBBiETvArjdjcVq+McLLElV78DQgA2NCzdEZtz9EwX9f72b9OSVVK7
3lUqVKiNcJpmyCFCW8iE589t41/ZSu1e6EpvyYKHXHNxXymb09/M/bsz0ruqEOwn
UlWdxcwyudEghgX86g1n+e5tMxJ3fGARvv9bzsWY4fX2T7ro7qun31xa/P86RWRx
rtS8BeUGq0EI0KB2EwtQ+9xzCxH14wVlMvUV2ySEuWOummfZYXriixxQLFvFWtMu
sgi8Y52Nv0OpwsVoH+FxwR9JiX43MDo6TSo+cUkZFHgQgxlCWX0MmBwOy8EPzLzX
9N0tefZXC2uwyD2l8C9NzvF3eCYn0jfRJQ+pMcN0qtYuhLUmBItDBrOb5uPeEPJX
Z6qanVFT1CGCkj2woBxSuhm2OETHkjrbZDro+IE1or5PHM/IoBUHKAoG4Tvqfh5T
3wNTjxgFjSLy2NbKIj6cSS4AfKSIY1T3Xp9XCeAZPoM1EVdbgYNL2076QcFEfHGL
hKV5eHqOLM4OtnhOsSJvsnyjzsG/v0/fNc5lQD19S+rS0VRmzqgoxA0jdO9we92J
7vVCcjYuTBexfhBuSmXlPH7sfvkNZ2dDnmqdeDe6IuzW2xQO/veTCuFzvctQmJ+l
sOIdzYOOIZTlxpYIwtmbN0w0ntcvISkOA0Cn6XeEJlOsDDlQlw5hE1Gckxk+h/8H
tkABkyWMuqt8x618gnCrCwipb/D5dpLVNVzHfXBChMIThTvi12Z/PGTrEurgk/i0
LlwpBRNG67t/toKFoQ08+W3H48TPlsA1nDz6U+5MwTeN+5OKmehvZ9KebqY8oF8S
b+6rY6p8z7uwmu/jUUVx4Jsyf2yisMaAsc0gne8Oe4wJw/Wx+8tciJX2quiU1+yH
4+Pjw/9+esO+qFAC3MiQwzNh/f3/uCjjQhB0gwLshhGf3uQK8Kkmm+N05WDR7ATT
d32PYPG/Lhx8QsKWZHP9fDqQS7i/JNyxGuzT10FbGpkCkVu4Zr8esQ47gbiny7u1
7/8ZkUg04NVLmT/0QANBKrvWcyj6O77Wa6kINC9cUn60gaS4zzkyhw2RPmGKevX8
CNB1YOna51hxpv53nQorb6zAXYn3ORQ2l+OR2xEhz8gkTnZnkx4BA5FNKx0RYnrL
Lsp5mA5GIFdNwQQc5LvwWyMyWuNB2tiEYQZzAywe+77npL+aD7XCw2MB1l6NlDT1
H5+ph5kT5MIeTGVbaNmtwIp9b8xGIrAqHsXOJnLQhMiJQRlUbXQGxMzAXUC+Xcs5
Lvd0CuDV75Fi723RkEBtHNCMxCuUT7HEAE1D1ustr6XB5RjUySVJZ8xVAPOLV388
yVvFSHNWt+MEbruTSWF+Owan7/JkIBYsb08fVMYW0HlJ8W3zhd05twzNl0yRXisO
ju7aeywokdYvNQiZ7Nm6IVfQelaQom29r2BIOz/hE7YKHF5Z1bHNmuTVq8DyYlEH
dTUanpgjUPJzbKFLZQBTQ7vPXWaU2rVn15B6tpL4Yitntw8ZohOY/7n+jvXpfZQe
ctfd9PTII6b68eGOj+41jgnGXI2K8RKsOBOEhBAYKnRxyD6McuJGMjZu2VwgIw6J
yDrL+BkBAXJ4syOhw61wgXy6BdnP8LbF3r8DFX8dYWA8hRctnJQLLRhOPFzJj2ld
QytCKAVjdEiLcR4jjqhna8dn8GXxQe3KTePu3BkG8LoxxHnqItBXKmALO8+ELJaA
nSwNhm3P0hdhG+5D4UQstTcn42YOMVNIIkQvI1f++AIJ8UVAOEKXUM0EGSArF8Go
K1TjqCzNna94tiQrHR9TNT/XOHkzbGzKJAyRx7xMMGe9G9TUYTLi3GjGrbmCGpUH
gqavCZD9ffldBtpV+NY6G23DdROT1LnNQ6mWTLN9ZTwvSKTw9lPv3d+z9JBq0uDH
2NP7ObUke7ByYq5QfHYLe0QA4vnh3DYp3nQNx9dmzhk5lyjCPiazzgKd3cY2lf1V
kfbRMQvc1V4izOuBZNY7vC7YMZYy2BfKAmj101F0NDehlJYWoMIimtThLsf6QNev
VZA+p0ywh77y99Ie2guZMN/XvPX22Db9eRan3qI+jtLfGO68PbddbTerQ8e3H3aL
qEEPkgPgz4rauX6uuN0t9nhjfZS+cd3rlPBqbMu8jy5qtCQjUDF98R9EJXtHVRxc
TSSZQsindsU4HsEvTzDHiQROcZOmgZxMJk8MRsdYCjYXqMZzrEHK6ShDvTPn5Woh
Wv5MmlnSrcKAYlq5YUb6oFs06zFDVbJBgGxj8NCA7lIh19EMdqG46ZuIOo1W+WJT
JP5zVa+UF37tf0U1/Cu6e01+fgIkCP0GycQgjS47ejN+f1VSuJ6kNNNoAjvZlcPM
YnZjitjT7LM2vEkF8br9KIcJVG6tffCLD3TTjMz6uTFuQGwi4CCkvcsDARYb2nqV
6mkIMDJmIC3vB2D/sGfcgDyL8GjbipbcvbvolNL8kcn2XOAIZYtm5db+el+XlF79
CDe5X94fZAxwworFJBa+G+XlzH1OAzRbWxNodHPU+TEZvW2PuuaN+4JXSoCv6HPw
102ViLswfe8nnzOcCqEMz7GpRRQMo8nwHbZWwSThwkMmFUHeOd5nvDIABpHnUI6B
isqYHN4vSZV1Smam4q6MbdQ4RDdP/Dj8i4lTiXGraj6J5845eT+INCdKmYqBKZsV
jqTEp2RWmyt4JFRmnrRmy6NTUgkbhvq/SlXbSszDyL08b+KR/TDa/b2LeJpGOHwx
fZj3jg7GBF74qI3q13TJKG7I/wwVgYlteZ+FAD8/rUkfMascps3Qfh7aoj0wkZOr
9jOUOSli5AgUybt7Lh8k6PtqE8wgBGIX+zFLnfkf2FSTNkB5EgpArDSCETNYq3ft
ObsHhgwsrJJli3jJueRsBMnEvapRUrrUSE8+GQb0tryC14VQvgpMF2LFbc/YXuqX
Eqk/YcLdBbiWJ0VrFlqL49res4JC+erdhsjolYi7lKYxARBn0QZJhIzFeRWVQr3W
bVAvUrJbWZBgUL7ujuZZq89MYETfr820SA5ar886/wEgnqqqBiV5/bYn0yGG+JVm
Vj7uDtO++iIbAVt/IGJHEp5dMbUjpK1zr0rkStK76/KuH7c9GXmXdoDLRoTY5XmW
kOP5TnB5eCTcGgxajo6+hYq8PIpi+WjVqkNsBUlCVv0OnFZHdTl75ps+u/XQ3dH0
2qW0y+Vn98liOgIk6VoLhO/3RYZJTVHlF2arP7QkJu0D2G1WUH7wPxhDupm9oors
wvP4KrXyQsu1/+kV/SrFHCVwVdbeXEIQsngFzBu1rCgLot5dS8GHPJWbyXirw2gb
B/1/3zxvcjybcobNeGpJoE5pj+NVfMnLCjQdPA/2lp3eo4o2givM7xVTlpRnoZK6
KjnXYdfX5QVGGioo0p+EnEydE3riq6+QnMbo6nF2EvZVxwBfjkgbyqJSs3I3hyyb
B9aWmAmw33/+4yM/Sf6F9rVPoRwDVU/6k/U80+d+VGZ8lRvFi/uMxNHF6q0XNVOV
vEuQIYnqnT1kNGOj/UwVJXcay+VAxTia8ZoxloCD+xcfvuaBHmEv+gWUpmoFI6rX
vLyRGW3UtGVUVDMHad6jcYYtfSiJ0/kj0lg6PcT6sQc1FiOfUfFxHd3L40AVhqpX
/8ab646a654eu/llgrq0JBa1c8ffVodKO9VIozwOTcA6TBEfjPLnRLhZy8boFKil
cBwW8Sm3RPmE0aSAsQ+cYITW9FBTdVjL+1rw6WxRQeHqWj80fNzqcaIyrhz2DeUq
Zefriu/OMr/x4Fmhd5Nng4/nwJoMEhIohTp78+DruaAH9lOPNbetXmzOqrnY2Oo9
fkZjKC7xtaLnhBY3WXGo/1svo6Jw31p4gWNOaTyDEmj+YUf67VBHBXjv+JoWy5/m
vHK5JIkPekZRpPfwRMYsfJCcQSd8kvkGQd0k9ADePIct7UIYqw4dKBZgebY4175/
SDXz2xN22lkxDpk0yYZQuTLsTWnEfsewiYYzKiYtDMCEt86bbF+ZOP+hoI78HT/6
bo6jM6bHwdKWywU1tmKxba+KQ8pq7LEx+2TUgMySo3ncp/R9cECzCWFDG8PNJdCJ
GwoeEXoMLd6RtB6xj8kKZQwl64UsY3nujzfzVkiigOidIk7A+AzDlhg0FXFMGMLP
3WdSPIcGAwudTv2CgIsJKWsNW+Os6VG50hwvA+mqgPwu3vhxK8FrYOkypeoDb6TN
PIbGgAKSBn6CPgwHArhhux5FhupTxXg9+c6JlwRD5+jpkUlxQhFZMYF5BCMAx0et
eUi0RKYsC3cYIreiSDOEtdxrNPwop/wakrbzWTym7I4/6xpsHzoR74kQUSo/itPI
2azM8+FkTIDLAh1BkO2jyV7NA3Yvc+1wzZnvlRANjPUgMx1xXKxALXgG2S23B3Is
LBQVM8mV/9QQKLmbHEwhTvNKTRLlI6efoSdQKwfN1i/MG5UmtCDlMlleUj/6O4w8
NiJH4745klC02UPAw7gInrVTUYRqVLrR2iMF5/jNXTBxdvbF9uVqwFTPiIj9wDxR
DwIb9zItika6MT804YHIsFwi0Thf8Z02gD5SZFcxzoNuzodMR//gkHphFnBVUIjm
8XbABNNWjYEjGFQkpfkWu9meySFw2jIMzG7R4K6LHtx0B/vpKQ4+HioCDUGT+Mw2
xhjyMcjZJpe1zfO4PyaIqipbV994lykoB6uQAyPtlGW0JEPbRnS5eGIcWzSpjDs1
NTm8HZsEgmoGQ4g00jd32hOWo87gcTZuA1ekrOs186XnSxRD0nBN4OQIKFFLYaet
wks6alLVMrFDtS0L+LS9dnnoRwWjxEuef6KTCPuQxXMAJRVFVE7NghKiEUahFoGd
eHBBBi0Mmo/gycjlLpDDTrc1Ir2FBuTJ0vwjHhefJMTmKhIlo4ksKIJBDUVzCoqH
i8zjIsKl7ehZyzcsXDdyNuDICaewJ90X/b5MgGThZRrpxeqLXJJWx78DS+FR51SH
a+KryuzLNzAGl2oKCxm8Pv/8rsCfVIGWNqwJ1ZmMITUyzYblIhXQQvaX6sHnel4+
e/tZ10tzzVKSwfXpjijvmzubld5sfJik4AgXu2AqIY+IDxGaEa5FJQCBm/XW9Xp7
5PL+noCoSpycrqXbTIfHoUnydkGVS6aw3+Z+sErx6snO9jeMdBTHEjPQXl6qmN+Z
79zn4YTyqngUxreaBKcZ4m36omEX0lujzZ2Qk+hZ+FGWf1lxmaWmmw7nIJhNAt2m
bsCNJn1KC76ziZnscG8/ya+k2P1FVbNYs/tFjAOeRn7MBW4yBhCuYcIi7bSMjWai
2Cpls2cjqHzYfSXPrXSzRB8qNfJAJis0ugjmhd/mRVDYYfJXN+n0nyKQ2HpG+bHk
h9I+PYKLNdlZVTsQhzx1M1n5to+WcXUMfltt8bFmEpfXzxxN7g748iW0IKFXJsyk
ztQmU/6/Hide0HcoWOrHE/AGaPkLzVu+hcfXemR4IK3uUjJgqegtvdbbQ2slySde
rueVLkD7H8rPKxyDN70cVbf0jz6TI7sm9G98+6wQF1qr/VhkR4xltz9jRWnS7BWs
it+6eBVpbvGLK96ZnZe4Mx9s67GoM/bnEnpyoBCYZGAQAPLJlrnzSMdzbJ4lG0Lm
Cboma6445AZKTVyE4QjpJwfXgv7r5V59MbbsU4l2cth+WjNc5R3dG28Cmu7J8JRr
8+rID+X8sXZcDjJuYrAtIvcixBww572kaP2zVo8IV+uzEJhwVf6m/bGLa0l1CWgW
h8H2XHyEBcoJUtGTkNkqOURlpIDLPpijnl8kJiE7roZaNZF8UWgCtomGvwlOR4Lz
UIW40zBrnJXIA9Ej7MevWi0p/M4ygH9EFu8+9iDhVemjxTBaAVNPxw2ZKHv3nOQV
lkblsXE3cz3dX93cwEBq793zGqNEpSk6jk/eU1ZwTuVBLHe7WECOOw9UsyZkeRGZ
U3yc0JoOkye0lfPc4KRc6y91MNwX6EJVALUJ3Ut3/HXMbEIBVOqMuQS3xgcgG/MF
qXgD5WN5VYiueOd1fG9cu8k33S/PSHyWKsDPqY5LlT5tY6CN5JCbebkWh+v4Y8Qb
E3MOqTA+bqD2MLVc+TxNQuqoV63BYBeXkVDpm29ccfhCR3H/gMM3b4tV+OETmDr0
cy0FXvHhdtSa/c7gJ4ntI47UFQrOYuBAI+AwMsyJ0Zv64baeLopZcCD6Ue8fIF3z
FHVuE/wBCXCgV0g7nnOOLlZ93nk7CSrSIxd88HSkld7SBj+ptRCPqoThkyrsKKYu
cQi6ti6HlzSKtudyPwcYO6mQrHqaXYgq/W7tcnsg/32QXUENio4crIPWa1hGS/jz
pf5rg9WiARD28wpehGZHVlQBWZEgV1gHGkeV2rxdEJ/xQARpHcXRyUxAhNkQuAAh
8eoDvQWgqANODgxSqkc6YqnX1o6lZwwVZkQ28UgB4qsf9Oy+b3z1nXVVUB+PhGc4
4gK9emb/mETvQG8D9GX4bERjRBA3FPgxmZKNhfS76l4F8y5oSSkCHJuRivUVDVru
xHoRwXUL+zk+0ADw42YAjdVSb+jGvUYfYXVg4fqSMjtBD8m8vebcmfL1ynIjIv8w
qt0jv2CGnw8pG1aaAGwJ7HDs+ts5keXOWT7Qljpf8GCK2OFRMTvmj/4RI2xPLzR9
OHEedmXaj4lT+k2qlaEeo2XbHAwmX0CiR0Uw/35ccB4/FIqGgkETClnYFXqZUwgh
Touyx2twhLqY5vlpjR2p3TCRz+/jxHcghbpDaoXunu6+hDWNh4FSawLZi6YSR/gt
xJohSvw2OUtFJAopPqL8PRA6RyXJ2y/E2W0tY3QZjl9a+lEy73uT/NzCMIXegoez
/M/8YE80f/SqH1b6ygnQa/2gSym+w7igM55NJJ0GgThOwfppmmlLaEmg46MKYDS0
HKQ/kbOCOHGEtNb55pHL1cmcT3ll+xM0W+oULOB/pzurKkdwFNmGeN93O86BfnQz
5KZfNtEBam/SKSGUkuAi5MqJWkAS17fQZxQvtGfXKbk6BpD61gNcExROurqGGY/Z
Xa0xENQ4WiPIK/dMZb1z4nEfp5zUItYTygukhAbXauyPp6W2uWwBHllPte/dGjai
GRz7bFkfq6a8gKoKjNEZTHm64b8qRLqZM/HTS6eWLO1tbUPZhbS/f/cVp0DOx3br
jYZkUjuxfzbU2P87Val0AnWYJDs76VNeSjvm0BCgaeYqRn2wCcHIFOWvLg/FwOLO
AyItkoSvd8bKpgmA9OK4zLLFfBa4ToOWl5cge2gigH+UBUtTGrJYDyHcxEDDVCLv
QxZqNNdJ6Yq9dVCx+Gq6Imgol/6p+VXTdOMPaNhJOWb5YgOKg7aeLYUBRug9U9Fw
kAS7pfCvED+rPaO6HfbYrYFMqv32gtz5L7SxzD8i/V9rLKNFhwv9g0Zpyanpj65T
g1U0UwodcdNvg1XCadSwldjAkef/loO9W8AApImgtMeuv6SC4qXTmI1uAYl4iB6c
it1ObWLL2VghDs/5LAf5hSpvc3/g968Ky1zJPNec9UyBfEsrZTpschsYFiRQr44e
hGewtUUjihc9MOM3HW1LqJfxZixsIDsdBJ74YVmf+VJl5YD4V7B4t8DIE0OvLbiV
ZDL7BhWonJWX0MEIvp+xONgjvD8ZmhGKbnTnaXQgF3Tpy3x4WQunwTc2FsWeS78A
ZAQzifKZJUahrh8nrclI6Pqx8QX6gS2B48Q3XunNqDAdHrpil9btSEFgOdOTPXzz
DMZ3z4WhrCp9+gjf+EDSXGfqtIUPGqkY8xJj5Q5yAvHOrkFHhOlcV8dqeCVCG9XN
dsP1CzQWj/Hg0jV9B+5S5JUhtvJs6hLB3Bh1YhTHAP9UivK6AgBpNv1awfg48Tt8
BoRA7Gpd8C6IeMIAMihRIJXwQNhS5go6ry08YiFTcdbjg8vcpm6RP4wCryOtPScM
Zd5kQH72P5YUFIrnt97681EPeiVg6cOA6WJIjnt7ezQK4OQVKuU7YH3Q9X40JtYS
5Dm3mt2ff1iQjppEOxZqbkK/f3fzc7DXu/3kEyAehR89DxOp4g3g5J8nHGj0Hhov
SjfyMGA0ex4+KcxI3vg78N6y6gls7DrcEE1eGvUpUxw8wfGlrw//+GDJcg5y0RQT
Hfhq2SZAurDNGG2GBf+0vgn32XofIGuYOmllCqHmSSsXPzPtNeXnuXBsKeXXm2nE
W6TIKw0qkracq8yDlXHylin11QMPeiMbppplkTuTg0m1h5Y2/dI7WYrkOxntWt5h
i7eUxdCQfFzUwHC4hu3e0IuQtw8xcS8B+Me8MkCfcyudhTolb8+zNdMmEannIFVM
KKFNAL9NRETy+BD5wRJ4wqvmIpcJxNTpAsFr8NVYZZn7rskUYXQTjdn+EUrIN4uW
bQAzXV8QYQOJqknluWz9vXOhB2gVCDrJfp123hF7wbq9ote/yByuJiNa8po2F9zV
qH4zMsAxUBwTGoDMr+5HBglNIgdKuzEbKCf+1OFHpn8DSpvhgZ6PKzAakd5kmDUt
FiUfec47Qj6DjVypv4sFriH4rds3L/GfZHwz5ZXRSu+JhTUI/wAJtShfCBhEX+3B
rHn5n3FOyFQ6lcLFpcO4RXWjEgRiC+PIEXhX/GOdf4VrJmSJ2ij0ei46PXNir0I5
MWeIfg6ZcuRC3lTdwRr0a1faVDJ8QKuQcV/IbfKmcTI3ZZ+JFJGFte+owW0Pai38
uqY91FYr5vL1JEEPUdZvLhWPVqSLXe75yM2FoStG0GYEzN3oRCXXi6zLqhZ9N/h8
XUFfb81Sfff2asOoeiPVRPV90adiS/FX7bKgPWMZUeLtqRlcnJsu6iX50qmQF11x
G8Zwha7DQYpcN1nKbBJAtzN/jQ+Yj4cI3c/5Vo62idB0p5LofqV/f9qXODYGI8v3
+2hgPjLyhN7D+o9alNZqZJP67cExaLF1/Lop1Xs6onNww+bNcCaIrZfXGvLvv63r
WNj48ZS3gfyD4a4vdGSD+675YWfW4frB+QuNDzlVER0vGlW2Az9x6U6/yj6IhqEg
6R19VKQxNiLrgrDnQW//dHlY90VKcH6gWB8aoTCIZmlYb74OnNbSpo4+g9XWkcqV
9oUl3TWHIbNrauSJ5WELoNi4K1+BhKWMNO0hMGsBY/CoSwr7AqWWfqMmigBihFK4
ZgTNzAAgRuIUK1Ibcp9LV8wqZ68Qgr1OavN7VNqJNh4KciZHe/PQYr49Q0aOHrrd
eFdNFmUJOOi0q6m07PfSF9H+hqSvKQIz2yc4m778YzAzns42hE2GCGN/attNtnHX
ia/BnYIown6pywyD4x6s4p3cmDRgmFoPXR9Ns/92QN9NdZuK/uKPV6t/osAYlQat
F/YyM+2W//Thy1zjm2y6ybVWycsbD0YNJpafzdqBTGKFIeaB0VMFSJ2xM3wQAM/D
PCU1uKkcO83Axm6rUor5LhvwVsVbNF6beCJps/n5OaplVmlJ8/oVSTnlL/o/DhqL
Hk0I0MciEjE3W/UjYr4/IgBJOFfz6fLUpHfGrJb+Uq32LIt4u6gfMehZJX708PTo
pSujue5veFGHYugu/j7c2X6zqH9Y8MuhLvP1PPojdY0nh0mpDaWTKKZ2Oa9vr3pD
si4g38vI/vIsoa4qMbXpOJ3c+FwNyx3Z2c1YMUmfNzIWsRFn5NWuswAtxp+Pva5X
B7ehRQf63N67dZrGzsMBEWnkUZ1jPB+PzjYi9pbXg0xTwgq+bdh+VvlzlOefH4yW
hoH3+2SJdNatV9sVC0pcw9niOLhrEjAcyVZZ1xcgQ72XRuoGJDnYkJehF24Chocb
dod7rZEH8KmRiL4PfMnbB9oYEzAsUR5mEErbTDCFZ2ApOPx+SnEDceeWBbo4ds4S
tsq+uRT+rIvUd4PEcpmTeg3qNpYT51OjDDvCgBWtjZkUJbq1SQ8CNXh9F7++gzkT
zSZHma6aTl6HDjs5gl6G7VXOEF4ryi35FTEpN0XK3CmVTo/GnwBEmcsxCUw4d55A
3QEBpYV1DOTjxzaV/0ZNeVGztNNg7q6E1qoG6EqK1mkfPn4jcbabLShboxtL09mY
Q/cKeXi4hP4rgg9MJT4pHh1K9CAoi2QFxxsmf7TmltGhB3SrjtRmqo46n1jcIVw7
ZVlgpTTzGoAH2yDTMaabidRCAde4QZsefM5gt0Tcy0koos8betELDC+Aj6GVSlLp
mG3DlO67v1RM7E++V/AhNlzy0D1bIPYk9GYj75+o2skuy3GI5ljMOVH0stAEozwY
bVivn+ASUjd0XXlstS52RrVVFGe1/cogDIjQnLwyH6PUZ3kC3o4zOZh6I/mKyBvo
+FdEsliFErVaH0tLhevG38RjAv+i4a31W/XscAifrqDp2nqF3jzVhC4CufbZnnGt
WSwEvfG4Rud4eCtgiSacsDyzViJlumrBNmAJzbl4KUOZfBJyb4L++RRLItZwSd/t
UJifPmjItSzmheJVskMRYnKhYsS5cqlhXwLTg77oHk1oXFUHTEqPjLW7y1MiSy9m
rkaaUQuMWcxOvbDyldvg5ZHoDI8JuYM3nBo8R7mmwGf70KGBm9FoWguf+dHFRpFY
3a2ixr6rWS6tES+l9cypm/tTUo1hLN207+z9cGNlqAglRMG3A/RizmfDWPr2gnnn
gWgMJBKdDQ9KYnVJ8IcGD8AyWjldmz4AEO2DIk0k08WqTrnCMLeyPAkEERp3s4MU
gY0GX8jTlh8DULDtoKxm3MhC2AxO5yjAFfOa+X0Sb+3tUEPQnx7sAy3837w5XwJg
FSf2p/qABUlo+pOkoU+pJhLbFrunEbaJcqGgabR5k3DczHvfTsgTB792qnzTmts0
lOPDPEjurAqaTPx/IcgGxs5Oh1F3o0W5XvikdtaUoUUBhOu0CJprgLIwyIqDnaG2
6m4ARLgjGuUjSBOFKEK1db6jcwfO7yoWQmxKu3HOHEdhItKxX8BE1qxCn7tRHbBz
weWcfztDZnL0sYab+HPV8YLFAvcT3/HvVAM4AnUgB/WmiLPYsEkkOZV2ke7k+syD
64YrUhLiolSTEJKAn5a71BwWtso1+6DAfi9Xe1qOuF7Lc+KD+ttlS0PHY1KFmNH2
L9sAqAdIPTlWD+44+Q26/Bpe0bM8wlzRAB2jA3Kq4ZX3WvG2WrSInhkD0nvTWpCE
rlmqLNB6+yea7t7SkSu5d1MuMtZUz9Z4B4Oc1I3k1WCtpaapn/fjLO0BXFYcz/8W
zVdo7jvoZSTs81nLZGGEt+VL4ocy6tUngjK5MwGwDeSkP7VQMnVv8p4gioa1qzjn
CaRm4Uqu+XCHLkMCFUgZBDKNTfqgMJwXqqxkL3G/r/5GME9p/BLRrJQrcsrcLL+S
5KJZRc1rzuMMFIjHB/W5Yl0WlHveOMJQzqTgF5Ac/viqphYbqkOtb4CDNl+6omDt
Z6kQqZCzDAUUW4FaOsCzvWPCuQmXqGH/qicdAJe0NWTbX/go4a0TZIikZ8uzsoEw
gi2HfVpJOwHceH86v/0ARx2cmwFwQ9ilg9Kb5V7d7mdXS0v8Jx9TR9AKZm0lnF6n
A26R8S5vQ7zmdcJBvvVK9LsKFCrJ9sSlJf9AyDSW6J+30HMO/IhXJ3fJjorFHcdo
yjn80PM1xdxt0qTiTQt0kJG89uGGjpnFR3E42NPdxADzmaCmQzIg4b8pw3iUJSZi
H0SM//AQCXXHXkTtUz5NStmSnDW6dKR5qG8lAKIWjW3A6OKYUTAma0AowT7Z+/7j
qxVFIGDSN0fPKy7lh3q6RQ8NW8DwGv4FQVnY1h8MVFE7gXmlEjSM8TkAolRqn+yc
G0GVcmDSkr1FFtasHtwvaz6Zbg7rmN/YGokiPM665V1/nXLy1xjlYTGwWIasRyie
DNbD3UPYMAt/PrG3YOhaROBb8CXwHmrKxBmluBGpzHr83m92U44Alhb8N0/oZBal
QP7iwyAUyYgpJPNc/J1RT4lcxtvFKEnDMyjMsfNkL259O3UlGhRv+l+izBXjNVDI
CRwZFz7tlYzH7pSjTwT2AXs1huDR7iXcnbZWdd8te6tJlaAvXgBTnMqxaum+vrZ/
DQSbajyQoc+hdbxCzhcfGA2Tj3B0pqzIGNReCJ/rCZG/KJa/1ERsKFdudIiVvozW
XsNuu817H1Bszy6X5DxhfhTn+d/prOtCVIN75L8FcZKsKhbyymadSzbmmB6NlLA6
s3em/zFXc3TdVWrGnktD9d2Y2mHF8oXnwZKXW+gyqcSAX8DWkZYHUYhXzz4v9gcD
GsJs+JOtEksauMS+J+9yiIcA1vczA4oqNWjHAn/4gAhI/LDAPUEltfOCSxlLGDqV
V/vdfiUN9FGdtuWzcXdIYgJkwdIhYttT/9rEtVYetEF12Nb5xC6ZjWrDnF13eptj
irQjneCf1d3MhztEyAY7uTeI+xe9lpvGGOOqq2enY4YirKyvKjay8qoGFqYSNudV
wQco1uh+QJrdaKH1oefhK16Fy/COvitQ6UPjvB+yWeTGF1bbCZJuBHmK2KAcWj0Y
sElVznAdY/q4fdK8NFUNU301itHr8aPlFmeE6AZE2pNUuCkj7Y8UqBz8fD5ijfV+
xz4HfoDLMGagbHv2yeZLo7+071Hr2zOMdY9CEGEDhb4jJdG+0Or1jcnCaqCEUyDI
V/fODKxNoW9srkEfOkxFCafe0rz9JpRIDyuZBvIaytPmoUGALNVcXk48FWaJALNt
K+uugvx3pIBfM2T/S+kkox6zp3GaYt1xHdq6DHtXc4ZKJaV89vzxlwm2KuHcWTDa
V+RzE66ILt5oHmmZa0EdIuK2UXbl2XeMegXX0gKKw4AhwhPqTDihILbHTp6ypOb3
KgUo8XLZLWZANdVIKGtF70zQ5o98lQBNol0oy4JzPNLFfDMPO3jeyqjO4X0Iq/Vz
7fcXu+k3A1Ji5uzqRcw5iwWyvkYVQ1tf8u+VW5rqlf7T7g58Ug82xWyRJO9jm3GQ
pEKUoatyGar99eBhOTG5qBpYhnqfaOG6E66SCVKkkuz3katLOQ4ygn1JvxhxWgSL
pZ5Z88dXPTocT1qgULrIMHx7K2ToPsZW4ea8Z2fjhoYHg+h1nazm3C0LeuY004Xy
E6hplDtJzhled9EPMh0qJjuZN7fj3+dqvjAN9Lm8CT3iYlKSocQsDG8xnfg8X5nQ
VorT9iDf04zQJyHM9fFTo/2lGfdMmL1GtmvnZzx8/stHdaq6XK5aOpbOaxwXKIqi
G5dMTtlSgt5mk5n3tqMtzsSaZoKLLDMf6LuNyBT63F0m+4jOmyWGdX0jJ7VYiK83
N4BlLaq5lI1isA77wzrP4nrwjGcAfICGAff5tC2F3IqKBcMQAfxNK1jo+K9dH/be
SfWaOcWn8qIvx75qlYHeZER7bazqQXrj8d5Z+N52QoXFDbMqS9XGuS3v1Qs4bgQa
YUP0Mo8VcyGDAYluGMf5hSnX6CIlq87KdnFyA5oHehbx8XgJnC2ElUh/x+yEexrE
c1qE74u/qhZUKucUiuG5sAtGjOJj3yHrS34gNfrbylIR1OW5cFFxjvf/Iz7mNe4X
I2jtN3a8SDXb8hDyEeOIKT/DQtj6U73a1Xv/+bIvXd19u8+F0X45X2HZc9mfBDGG
Rj4BKioaqdLxzUW8Kg6q/QtyaXsSlArgPbnVOCpCXm1csYXGwmaaRb7sHB9JZx7Q
lQEGXKxE/9UDHUP+juTDTKjB6vbU7Ieqq1VxUowmG7GwRnqy0n6BNUn0tXKNxdo1
7jDSHI2blQoVsm4K59uUNV9Ai/Jnk58lINXSi3tQTVb9zLzz3qRvUHHMoyXkRo7e
c8RMUs5zWG7h7ILq9WgeZ7qCAv9p24dfMXmCp3K12Zr3o5iKta85NUqI6+qlg2Ss
qp3evdNrtkptKDQyMaxnFOn06Z02X8+or+V2JT7eFEDtvAIb3WQrm9Tnp9y4yjO2
US5IypgpluQYAEdBUM6L9FcKEDAV+1Wbjl9X/bLtygNAQZzaS1VmHzm+FSsj4B1e
chOdJOPPVnYt/coQs0rTDokJ7U70Yc+JI+Ytv41Opx3D20DRD8flzZJnAhVjHGKC
lc07FTb0SRy3UUKF69/cBnV9+ZnJ/yKKeQbrrEuvWIMU4/IxUnMGWVhgSu1xvI/A
iXjut3SpuiBGYk7pFzMQDR7gTPz5XhhgrjqdF0TF98F+wu0qpn+I5GVds6Z/IAKl
tXQQHjtHIUfophbde+b4kkA7dU5Vl+Oa/WkbtvooIpIMDvBNBJ6OmC1wZVijONpk
6uB3At/W2tAqVpDvpaMPxp3ESxExY++wyeEUGDHVX6DZrGgE18H1UHEbGEijo/hs
hXX4s8pUbeT+Rr7yVOyaCk+k94C/aEeZnJHQnTl/zkmA0CvvoRCAY59a5R0mAylI
yxaAze5XHEItHKJ2clQVaTPGO6nOfkLLHieFJaGBt62XoWp9PbfaZF0sRYRTg5WA
1l7lBchgk1V+cVIlcj6t8auJ6c0eMkB2rTy4fhPjH33tSlJbCtO6uz2plm9Ov4oz
vFvff3IkAt14Cm2OFenvdh4Jw4ZJJ7qcdNbpGwb4jel7P668MIULzIHqr19iu8Yq
Hr+V84D/C1vcdGKnUpHxfaP2gw4dkqleTFarnMZkhiqM34fBfLPwffgrDSVbz1DW
Q7Uago5354KPnJbMjR3eMmueJO42j2fGrYoBpr/ZPyZm50tw7EyxXVha2jkps99e
sEmXwV6+1Y/NgXBTfESOTp6Hg309lFTlbUVmWdei+gxpwAcQ0SUlfDos4JMOvfBN
+JhFNw/T+i+lpGnTonA4234FIlnVKdGFZruBnScNzIRYzyUOVDJ0S4l2jszz4RLR
s0rsbkXFgxA2H9vb1DQi0dkhuQVcFacgwkyZKMXk6mdQ61YWJj05ibs16PGb0Ujp
dGRVqfvhskJrQfPLectFT3pO5rpeDZPX1GWexRUT8DXeAj30kYQwBf9sVZQBN/Lk
7nYOuw4WWVc+DTWOfBumwqvItkKSMEH0Z42GE9kJ5NQ4IPLNWZP9JvANhLbmL0O4
Aexkm0Pt08ggEqywrmvLimjahISXz8AP94363u+RUuMsGk9v2XtF9T+UHkFAPBsT
gp9IIIs8zLcd3pZ+419g9lxpr6xq/mjmPUNj+8RujoT10uFqgA14cKxazVMPQWxz
3hq3JWhWikA8WSiVcgdKN5RG8jZo10u3xZtj+CZhL3Jn66GfIIERvEddwZzVATqb
QVOZiCw5EuVeVRiPV/unKzVky5DC5HVHAejPgbNv7FtkbVReDMrl+u42i+QzYjzZ
BR4Fkagmy/Ua5FnycD968lO6poYwW0mUsTa2GXkzQPrIcZOrY/D0G2m7bdBTeMT2
l9TWjhWxQLtiI9ZqrnfaXHWlRrwKSIXG4qTr17n+UXjsQ5POsH+Y7uOhfnmD1ZIu
6ju1Lp7L+4vAxLpYb2zoIPL7Fd71FMBbKsFMW0gIWCFed2Z34s0ucS/dTGgASIf4
CRCs7+opWAM0L3CXsHpoR6PbW3shNUVb0krHBIy/07qc1mUOruh0eSkZn1YSMvU1
viH5AeviDFs5OhfHnr5qHD++stPhO8263tvI+qdcisEzIFhRsdightRF03S21DuS
aQsl25inu9XnAhhmSr50eFjfBgw1iBK5dwiX/NzUV1PvN3EG/sLo8X3zdBZeq57X
8hsqSh/E0o5E7WijpUSR8D7bJw5HD4ZfXaYvo3MuIVj47j6oLZUILFEg0vLVC7lt
BuwjXYiqH5QiLSnLOawwqX6QkVSGH4fhTA+OwVflu72/ggW/RN4vtWFxWml/bKmC
4JfC20Xaasc8/FmtjoR2pF1P6qMHppN2aEmfjPNQZ8UgeaWPrJ6Tsb2O99WE//9y
mk8/m/I5nFQC1GgT8ngQytD/TWYMr9f4XOqq5fz/5ygvAznH6a2T1n6XU1s6+ZQq
hk+s1b8Ng09iAJeJAYG8tU3LMXvvrn+RkRbcWpe31v0q8rZ/AF2XhrUgNjOv6Z2u
P0kpo2SstHhK+LNhDsMYHJZqonI3AcPQkZpB7QFTbzEMINUE0i2jDZ8yAv0vuTS6
OKyObehzcqhEI2r0vwNM1bRRSpo8hWbdUqWhfaZQrLLaQirNWcCwT9LOsTWh0Pp4
wp/0vs4IUpMlsle7OjcwQCk72cTcr6djOSDZHLbsPrP9suxEGeYlEnuIeU+ExZoZ
k9W6B2Qy06F5yaNJfFs74bXUzkm+kFrsD13yB/WRYRj8l7XkuuU7D3rfvfJs+fkB
LmpKHhu2w0SRBHHs1voQfqDuz1CQdVdl5kenzsanmtqvTlkJ5rmrynlOPFVXl5zb
69IYsmHM47i7ZPmI8fOw22fzZjqBElyX7meXCVrPVCPKUZ9t8K/R+IPCSdqqAIAv
dBt+jzWOMNREB2dMwFlGDc5dag8/kOjU+QHtv2CMnci7uah3q52bMP86mGqZ7mQ3
bsBADdMUtr2RS+HtbBeNxYDYXk+gO+rCZm+SX/j72kBEO4uYoSo83l4rNasbv+YG
YZw4WzPVoh/q/J7KEfO3kDKq64BpOuV8UllEeH9dQ82aygkH1WFfq1pJnLce5O7f
Jk4cFpWlAriVUqd+nizL8Vtz/ZMfGMnM8xTy7UFMiLmLD6jBig7f4KN0hm9xyoOn
sjwvhTTEi5qHBowrg27u6JQpvCI8y4e0qCk/xr1zdvuU8e7Sywl3L0H3mDDsRmEV
BozCZYaJbmkDVmIacatcekNCcsI4CHQOfAsKY2yZwBuAMFnG8wEZ+euXDDBBI6MC
wDXfso86ICN0EYFSVM14R/xCJK6HvVwR0VQs2b4I1Z+fvB3MqORAY/6Sz/Nu9b9K
URM1qgzBDG43a0ro1U/tle+zg5aAaonDChy7kjAal2KuEpH5Fe7T+oyKxQTsV7It
Fp8rmz9HMU888jLPeXcTcl6dUSYEOkue/+I6gkP0bJmK92sOlzp4sOX8QAt3R5P/
lysez9+yQTFsFfAI5JTA7dmU4k1gveTNAYh5j6nuwFsnZXpWZ4zSFVZjCN2Gc4PC
T8nfrGd/Ckmj+Gr0wAr+pIqTbS8ZFiCi3MDj4DCrZm5i/FbeAWuQ+NYJVsfuZW4O
ubaTDBA69DDa9yie9iBGqFKcP1Q85IzGrKh2RBcqVhQpxQ4U+dRhhjJxLkUi9DHN
ohW3VLfCHtMOJrMXlRIE19B+6LQk+d8Tj/LVjbaZhmm4B72orbNe2FqivVtgA6/z
zbi6ocKNpOzYuhhKdQsgoj1C4rNWRl32yRm4Gb9e5EF2bj15Vd3Q4jc8i+RcGpny
SYffQiBsJjSpV1ZATquRdsUuNJYOhZ15BVYD+Hpi0WD0waQDcHDlq2PCTI0K/aPr
Ax8N8/+f3RaRvuHCGc0m3LQJWzgtzQFACoxn0HC4rSB7Os2ALlaWbAzqaSQxQolO
2U5GGNCKqdNb1X5GE9G94mDvDg2J4QWwYarQmZ7tEzuuAnp2Dc1KfXJd5q3s9lql
XFbx4zmWQL/+z9PjHw8gFe2/Bk0KM4I6DIDpGVGpYYs1XQJbBbiIA/GHF1GNaczY
OrHfN3Hl9CQ7wkp/h823o6UMRsttS1OGDQSKTm0/IEStGCaTYOwGPSpD3ejsu2XC
RGtDMaLBzNAy7I1zB2TugqsVaA2AcOhZFvQg8GxGUggrlmc98yjNMrtN06ppCsp/
ksVGbijuVlNoH5hhBXjZcp9swXSbJXKPYgoUMwXTQrjFyMs4+t0+bwM4LfuknGMe
2aynjSC++fPB8xqxVGNxJJq82Q0ITO0gU00Y8KNDEVeAd2Rk4k77tPMnT6Y0kK5z
FlaIX8k2TGFmjuGQLNCtk9w0xmGjCHI+orBiuUcTjTl+EczXz/mENzVdL8JhilC7
O6KsKj4bxDmYy3Y1Cien2udjpVG51JEkxZ1eCQVOSqGbb3RlaIMCnI20EGU6UUXl
KTWQNI+82yeKMZOUGkQvQiEPhVsKSizCRNRfvZfPtDh3pJZ0W3TMsZYamAKytwTb
KeacKv8MXlIQSrYvfAO6uTcIJ9+Q1pmS2byx6DofD9NFvpUX6KL44XB1WGjos6nB
d3/IH0P9j4CPcJoZPztzU9wdbsE0EHP6j9kqMbczU+dkF9mv58CTEegeMBBt7naA
yAnDMNTOLergVE0wrvAXG4SHBBFMUx/dA7AZyG+IYeo+QvcDjGJVOmL7ElPszyG2
MiJVwb7l6svifktexi9GAABNQvVJ3c0b2D1X0hAh6BYw3HZ4w7GYY1zBCuconrMx
+BmWPDov6ckwR+fMh0HGXBE9en+LdpibnZxvKUoJoOfe+xxZD9pMR5eFvK6glHdz
Sv5JMIi7MTeyX6LwqXB7+OjqW3KnW3LcN6uxVCQrCyg3xAs0GBlVDg32be8FTqg/
xU/oLrA5LJAYkDM8VDzS10IUdj/AsFgEqnXx0aXWt/+Vi0VNJV9gYrIdu7rgTjkx
Vw0aYkU9rNPvujSMHvxXRPgnxK8iMQkFYolB8bA/QgOlpoQ1jir3xiXqDBU5Bi07
08KNI9IYSQMGx6TD3ptG//FrC8bJ16X0OSZ2Nl4JE/8MDSry+bCCADGwatK7t3ae
Cu58h1WVcLCHbH09Eq7EnJY2zp2XEG9isXXtjHKZT5q9s/GyUUM6wI2cF4Jm9cRJ
yLSc2k4P1aaAdpmGCU2ubzyMXe8jTedTNLpZWEk+eOwQx8QTPH2Y1BCfi8NSupTM
xxNfUN5nI9MEyWmvlEmd0W/S22Sx12AEhnI8xma6770Vv5vl+IZ01ks6d+ssOmTy
aNlQE6wuG00u4Z90EsGZvZun20g1Edj4K2dro/P/8pMtwRpwQfWgEcV4lPF5ajk5
KbjFRbM1gU9eyeGLCc6mFiD1Pl68fBK5BIi2pqixrQdYeHOEXR3ECCfObURav/OP
8YyF3rfudvRbwAW9v/xRVASI3UdpPwJr3Iw2qqIc11MonZTIYr/opJnoWlhS3MGX
OLKZMMQMFM2FBnLNhRAz4RAlZqhXaYloE+TCu9cR74hih+Hug79r3vFCP23Z7qMq
uxb5SgpegsxE9hDUmjQeONzh+rofbTjXhc4n20pbnnnHpB1GLzikay4Wr7RXSxjP
469D1nv7ynFL17Tt0aPlTZkggYtqv1uHEr7crI6N95J6qNGjlKmsiV6c/Qh7GNeI
8abNn6NK7oF9OdYwxW4S8Lw2Oo4uaK3CXFW48vAPDQBdIz41b7XA6+5YyCDw4Pt1
GJw10IbYwOJhT4+Q2hSBWlQv3dGqE9O/qY5/U9j5t+pVhz4Kb4RphANOKUReqSgC
0Nh+JzWpGCwy/XCz0q6lvCuXWkZkfrwStdkw2M8kF1XIaBgwQsIaSjIi/0vUnaHK
6hSX00Z/H5dODtqISlAk5DBJkB9s488P19a5LMZQanRr0m1Zpv6dSBqIDp2cvMqG
gICzGUgM9ETbcqRsmzL1JKeWG0Y7ph4zHoJjCfcuRME6fjY0uDD8R39rouItLdo1
aLXVBy4mBZaPIEo/Kn7LvVpFzqQ7CV8VjXlnboqF/vTBTzlJxBwXpGlRu4dhVQYE
rlabCI/LW168V1zI5epATuMYifFtpunFMsOCUwa4+GRIQKfyGs9lXKbThVgvukZz
j8QsCvzhkHGgV4cu5jFen56QId2ZJjidxHeU32MQOOgisuY+16lmGUwtxSKgxbWi
NHYwDU3O3zl9IzCtqguvBmAZjVQiP++rPYJLPADv4MT4UtfKGX5q3QhbNsV6Q9IZ
g1dvUWuIVDmDDG6PF8cNmGOzN8VB4IXHF/i9rCcJbKNd+/9L8twfwJH7FMqdAq5j
G9XQZx7wr2ZNNHGY0IwRzw2eIZQCV9WsA2GcG2PQIjuRyajxxhWgXDh+OPtsYAx9
OFqTmqSOjIgLIkMQrpSVkJEwvVazM2CcSVV68Qgf1tEd2hKcUCRn+ePCr8IP+HHS
ZTzOgqSe1nqeVFrWzTU5QgkI4C1r63+zkd2APbZUq/w03d/F7yrd4dfnLhcl7o+u
VpGGsLjW53pR6/9sreV1iDUSxfIIeqAgbADcgtAffhB8gRcA/BQwBHB6eAky7vX9
9WrnTsydBkrYPy4eFzu8iesCkCXDnfKmR1bzLZ/Vn6w+FuXjPIMFH1QXjCh5jn/i
TBsRoNZ9ks7OnjAvf58yhqD+t2YNAip1lVymSyaLj/CU6rZ9ghn8JpSfaqsoL3h0
ZyXFJZW3Lc/0ksOA0752rF2WBaTDwmyV3ayLeIjdzj+2jwGFPwe0q5H8zvN5dyL+
LL73k099HG1TUnTczLcjZX2N8gDiQYXzSYSDd1qDZlBeuQJvVeU4nEYH+cFi4/vK
/1Z/3Wjawn5nRphNd1ojAPxq8sUrMJReFPsnPCxVCNj2bdFUUFqGbVvzeZMPp4HP
k0+Y9EhQKaH6pQKtzuqzJseXoWg/Vc8qxCb2w81x0/3sC1bb+d2H4DFFQy2TznBE
OlvmBx4hTr5HXJXy3+Qk1eV0p2++TCqFiez6d/IhWD8NEI68hkWfJ9tXRznb2RgA
GLMeWgtDEcq5wjjcQpWi0zipCwENVRRybL3CysICePjnfjoc0/uL2W5srSQlKfM7
35uqE7Q/42OJMXC8rRntFOnFqdrMQLnmzYo+pqJZbYLyPbu0ZCoPLbpRt0gf5Y16
4XgicZbdxjA1jNgKDc7phJ0FiYvInj15fOOw+3SiRAPjotaODtiKL0GBJ7isOhkg
Nl9ULbBL3TA3iW9CIPd8C3d2MKUqoUFyyP1bbEO+ELXkPVIdScCaWXeSSV0GHj92
AW/nWytHUKkwKUzulgyzNZuqnhG78djhfk/BOtVTTZRylUjkR4RGh/gl25LSIG+2
CtgkJPFi85CINgpCSt2rk4gvWRQ6EATAQxqkPaOHPIPfhRWyb/p9/d501TwoVeE+
SWqX17drOnYb1F3Be+DVWcKEKW9x5pG19DCMNJ0PPAqjBe4JOrPpkGTYuyys2BNf
fMGN0ul0sUNtzcnYz4bkIbBpSc48YRok0lh33fdGz2667HloH0Pvkv2HMtQDmO7M
NqM5tkwuZc/BAUibNT4IwtUAtKabMZhSFM+2KQwkcyvI3/pu4fQ88BbFHcrmFEc0
rg74BMstOVh8BNciu3qlQLs01JkG1pJA9OsaY/8vWAh5udXzcXcvccseE5zgkCSy
7Du3tk2TlIe6okrWpraOwMaVZSoQWXnKoW9S84tXY/LALssYZj1t8zLGsRk36sZX
Q3oaAtcJZ1tTNEUOb/awZaxc1rG3XehYqPApLy83Tl1LPlI5yLiIb5/sKIUcnCZk
6c62O8CTv2M1EbCeBl2njj1tcTE7gAJ6X5JXp/jp9vo4+WyjcdWQjLNRt7TabVfc
MoUoWnfSNNjwzAb8KoxqwTV0ZqCAhbiUrrLbbAIMX/2akh6L+TEt4fQ4adY87vZh
dQsW7AgrBNrJmYFAyb/DxeVE2Xlbz85zCE4wvmqNEIBd19GVZQmFNDdVmkd5xApp
4anXIzL8yOCB/+y/seHMNOdSJ7vPwBYOU/KDgcJwZk7jigXZ9B0ZJZGiD6iGxNYw
TMGqpzpgnYG2qL81X+k4EBq9UDekmx3lUQQASgSeQ0Vfpn3b4tk5fO3e1XV6k9/n
heUtfQ0qJEzlz7ylifRUVqylhZkJBhJqztrzAQCEI/1bHdiww8peQpleVBTYxfBL
g1GGWLIVsokA4sX2+kdEw6+3GAktYlgqwrx4FTto4uoyFkz4Mndw2n+drUjCfGug
JMS/zGwB9jB6ZRhcAu5kKfINW3LTP8kD1GfgwqNvJ4s/I+DVkAwgFtEleN4xM9tP
uINTPVFCsJx/lzBk/QxGKDcAZkJhFxZNvzNo7tgIZuVzWYAq5BYKI6CGwRj7llTa
OZh1iRDKZD2Vo9xzRI8Gq7sFWbiMQDPuFKZYoPNQcCvVEj3TDuZNPY+69RhBxFTP
buksMp24LhczsayT/Yeb2RSuwekLQ2e+QcLXBk0y2QtjHclkNmW47onF4MffW/kk
m9UuFLzA5ndoxdzFcNyhtx/weIV3Jr45M9Tfm7gCKD7fRYXa47zfMneXc/IHpZ5Q
KvKdk6FxYZFxmZHk8F7MhTKI40XYwBmCiCEYO3YG3foNDa2rds2yhuLTCvUOPJsp
hXcr+FbZPDYtSDx6xdgnk/RP9eBmUYOpPOlp83mf874KrCaBYxgl9/WAmgr3tmZj
uMuJrBCgIHEWuGmN7h5K3xCP07xEnWAEZcEAAed8V8LITqvNet6TvUKVZW03uQbX
NZ3SdnL3ksEqV2sMy70TSkWP34vrEi7t+w4GNOSHWCW0lL6k+7Swg+zYGAlQHcZl
KmQbliYljxWfKGtR07o484z3P0DVnw9ESGAyKCOOCQH1HSRteT8sNC4GD1Fu4QK7
uyQqe5p+FlWuP4szBE1xHOpcuWeHrVw0rnvkgva+At1lb+N2GD9qnpjac5yFhjoo
UZSAJiKFYUD2qCh1u1NktLKz1k7xXelmf5ygwANnGLVLSZZkO2C9tV1O2mmYzFUv
zfN4D0NSx4LHOPi0PJIM//F9JBnzZ/1IiV7bHkVX0bJme33p1h1aKVMUPWEI/PCT
PwE2gkIvgfc0e+JGZDdk7Fi5/j7lZ8cGSyKVduGmXlNOEHVPx6TGNfwKBwFPl8eH
AuI+zyCeArFUrrRR0jCVvIRamN3rAi8rLiKFhmXVXLn1N33c5oyi2N1dVVBz7JOc
pSOC121Z+NZ19zU7ZKJoO5YIsJWf7e9MjJgNyU0KT4e1oQg7NDh/A7NV/qnVYFs6
K6dOzZR4gXvg0GUiW1n5QId1ABSLA8RHvOmOZutQ1f+KXGJB7mNIrOOGX2JEZmKX
bWvsS5tEFSpL58DkUJg+xUySGzqaf1elEJb+GYBUizuErrMsZekhx0TPCywvf5lk
DxHcJRsyDj1mhCkM9AuGh8jJ3wLLygdBdH46k08KYeTN6S4AQGjGHqUHYe3MRfTv
Rzq2JYSjhOGz0Cq4qcGn1pNbIEJ8wTWJR57DNClS59TDCPjiI1XlUBNoD2GKr2Xl
C3Gwh3okxtGtFMbqZM0DBSZUg7p3wQRygnKLkBsnJ2EuqOfQLsxdj9/tajmTIUON
JzMyi8nCZ1wE1Ss2GJRHt9o6LSk/OY5hAAE80aLTpKB7ewyJ1kPNOFPtlZ2gCp7/
M5ckwpFMGwzWC1Co3GJmMugUmfhsgQKXJbmYoJKC84o+DVqDv16JUvCJ74SEqvwC
Oeq0xoNjkdjppCopez8aM9RInIPotuf2iOE9lU18oCeLCclwr/2A4E8oklu1t598
euQw1/s+WTn/h0xQZiv1YGlPnvdNIFcJpsPLZNioaxEHKx/Q1iGVqs0lvvigQNzs
6A2l7gOijUPdjnRAVJmvLis5bZQxL7FhFaevpISBCI71zuxzHuP6O4K8vwSTyyNc
CDMSjOOH7ljjEWK2yx87oTQI+PHxGs0EZlWNiSfWnCfc9i8ejdtXY3oR0FokQAK6
3+P6HYMwPE9d88rSRCs+EQsbj59koWTKdBnjZBw84hT6IrEt2Ub1jVimdczbQHsM
lD5c1itf5RqxkextMrKYrSSbel/p3h28QJvhLhqPuhRVN0nWh7kdZ4zGYuiVZSEc
NlnhIGuN1W5ASm6RfhVYZlOC2rk88enhJjmCp3TVLYZ+rv+WYO2Y/0dv5pSOldsW
XpKVJQ8aFM/g5SEj8TP3HMPmHWPn4yFOmg2iXQKsiWz2kwxbv6DAus1eZ8QsoPBf
qjdXDHfI+YTf9ZCJ3MN3FlZ/jxoVRpRvpvS87eiUodPFrih/BONz1ab/L4uBfwsz
hyj1cxsPrzqw6eyfAHZxR3/7ZsJgv3fh80N8UBedc614IZKF4xyRblg4o1MkP6EX
/za0MJDBIz52QX1raW8VWPJiaqkUp6t3/yz13FsjRPGVt+bmibRqQ25zaX8Qmfe/
mizH1LkVM0xHbL6PMC0fEF3N4iMXyQ/OLo/7N5blc9mN0lt7lCbMm4aLoeGy155B
FGsb5Gnh5mNcSX7gy2dBI1XX//ofyJtvDNxorpy+jLELtj5K8RbTsbMt6Qvq6NCy
zJio7zAWtQeugF7GC0ft2ue1BcOgbGoqe7m9LdIT4NeUlZETCHsz5bFLzIRw1zmK
ciO4Uykn8B+ButTjSp7oWcyD/hdQmPt+5MQhoXbiZ2y7TLQbJ3cgbB80E0tECoeX
TSHjMRPUALItlJPSj5ywnQc9Ctz0KqhX9GFTYmBXuAqXO3XAu87vCKJDuzQMQh7D
sAiz/vBuebOGXybv/LjhUN5JsITbLyyM3g0DaUwQc6tgs57JjuwBEgdRff5YVvH4
YTRwYW0TvJbYRZjZ4oOj1z3Vi5+EDwveNIPcyYy+SyftUUTiGYD5lcFJrVcmkv3c
BmWrfXaG2HTlSI3LrTocdqj2RCJ+naOoNJu8yOqkfb03WxiApQ/nb1HTJrr9W21i
7RXvko16n4Ri2w+talQuL1coWWxe9NI7s7typ/89QHnh7XW8euMF6BQFj8AaSJqf
HuLUSCFuo9tiTsjjYHdyaDgT/saOXXUo4w/06vFAGPASV8BXPJ9N5YnKvtRGt/kB
AEqYus2bTt+LuXMhMQcR+brd3v61Yhj+wlXwKJozdoM+NkONeKFjIMHKtjoXqm9S
lO5J0BiRADYJhefXCAawzZTfN18uInuFhsHoLq70i/gHB0XgLD1u+lmfoiP5Y9ls
QB/6+r7Up4jXD7gcwpoKxTCdyKi5s8CIDFYNmU/SIkNVKIhx4FHpWVDLsFGrrLUu
6FnNRvbCN7ujCljMar64pJyw0t5GyY36PzxP/KDGnWW6PA01pwY89AgXJPo5wEdX
WymTM9jprnnDrG3oCj/QupmnHYNaNMT0p7nVl2U5tuOe/TC6xse5BAIt0w7zdDvM
BBawGgJyvVwJ1IbwsyQ/5SHVcxuk+RoPx17arT1oNCIAYV1AZX/N2E2OfcQTqtBt
+F0zZqNHGNsvDU2SJfssfk6AIOCm6nqha3tEdNdlptAfbU93mlwcV3bNJyplqQ1c
4Mg4XGhKyFi/EUia0ad4/pjaT0Brsg6DRfzjxPk78bKectSEwpBOnpOXW+SkrX08
tbasewhk18xdcU/9uvz494t4r038SaNaTStDAHC/1iksRnqAVaSZlFQ572Hg53Ha
Cn2tp3TSHveDkiWsTGWk31oWH0p3aSBeyaZv8soNHkGK7z827LTKECjvnHPTtENR
0LYDggHMAcDpBlv1p5s5xx38yiajQzDGH5U6wv81vGh6RUv+CTTNfV7ZICGk/vNC
m1x14rwOagwyFIN6LSmIdYUVzNederYVEs7lQDS+1f7v9aWFbSpClTclAs0JhWkB
uwyNX2x6I138b0ewmjh1q0XOKaNZtlKupgWNysbJFthiMjfpcW58PeO7dzxv0yVe
SVGkuplmswnvxc82r0tHCi3RSk1Oj+3sqFL1VmKlttUunFOGVinMuuMnvTXP3YnR
8iY4JvMTApKyW0tVfzuob6/fCehFi2rG+xFq98w5nEV+aq2CO/KmlWCWSF6sTzPW
dCi0YCEyX1F/7gdth37Rxq4/OT6mg5T0muLZSpPQfgkOS+8t0tyrxGGnXaevVxXf
MFD9coojEnQJn85Wo4nWONSDM1mjHa5A3jAvqmr36Vpxg0vr1WaDLDEiF4jcbUvP
jNQXFCKisFDPb6+4lQXAHMgd2oIXyIrgBn9OIpCFFpwNufpUctTwSQuimp2Nyd9+
2qGtrFI7FnvBbDMd+6zet3h3Y2c7eXLVyVu3Eb0RH/Rl+5DqbSe3yD37Wto9qPLn
D5Lj0Kp6Yrt9y6Lchvs2AGbOsPRIXr9ZAJk6j3znya3Ffm3/PCAEVm5FlwPin0gk
VYsmO2QwEHusKiuGIOAfDLbdQH4P0v8vaT7YUZDC3DFfDTUFw5HBWOOmnMf5BF3o
p+1ui/e3SOU80SVNawO/0GiLy+ZF6OlMkv+5SNJwNWC5BohzGm7Gkea/qyzNVaGH
yM4hdFcem9i5hUxQ5Ut7SattMrI87RcIkgiQFIv3w9hh9XabUav/8MPqmAlQ+jRh
3FUzLqag4OIBxrPXibclIVbzeHWBKJWeOO+vAi1NGUSdSGF9tM73fqvaIc33jl6T
qbOlIuCryaDE7pIckr/9HF94jtUM8XpQVm/vvyykxp2BlqNHOveBIocO9UU+xa2f
vQOJdeWHos57/zx5U3bGANdPkCuEVW6Je6Oap7pWmyeMWLrXobTo78pgSzI32KXS
ziFwFtRWE+zJ2xENKmNDwkvE29KxNxaBXwhTHJ8D0Xl+vYLidIcBYkVox1T8Ijw4
QWC2IBuQptUxgRJWG6pmf2beMkpZIdmcvHwrk9UAJGgTmbF6cnbNcbZYBHEh1Wrb
nRSPuRDkudg07xkE/zn6NYADlGPJk1ZfEBflcYTHGlfMTNmM/ay7DXy+opXREQpv
3wz/QObuKhKnLUV2rubGoqWUGkGgFOrgnY6Hzmh+5xY/rE5BGdusJl5SzXpsawZ9
DlEhodiBFrnNeWdbA+W94BNYyrDa+McYzQxi62B8DDlgCXK33ivxFp5wOTgJ+PdS
jCLUn/Jp9i5Os3ShYeoJBdMMAAdfgOD4gfOI4Yk8gE4qDSjr2XHnJZq3cY20IE6Q
AFOjuwMV8RNc79P0iDZLe2qE498k+dSE1HMJxuEm6k1gxw1vvqOuKIS1pgkp6Nqx
6J19K2EqsuU7VGlRVGQAej5a3ACAtaSIG8T0xZOq+qsNX25WZqhMV6thbpq3AvQb
srnQvqNAWyzDJWp3fGgXecgWFwBxOJCOwk+BWonu9ry/6D5iNAGx1apabt3GtbAe
/4RvJohXJ8w5Ll99PCq+yVFwZluZdBChqceb0+luxMNgpPd9fIktCTCih0xNa65U
yXFD+uQKagL7GLktyDGjaZnGvhUHTq9DQ/J5RxIa1z5sVZkzowAD6eniZeTSIxCI
2pokW9Y2X1NzLgge/L6mWesKZoD2OxSp8QLLZurROh2hdcGLbiBR/6NjFkjSOFoL
YH11gZB/gsI93c1vVL2OBBEWznYkm4Y80yH7i14RJeUT8fEOIlkU+I5PyNJ07Mf8
7SD8qUCYoTBRWVttMamZ4HdAEYpnCI3n3E40NF5buJTXC/LpLk6IoqhPYG6nKwRj
Gs/9HcYU7EqRp/EqjNfzJnrhEiKy89FShdHtln4n7QCiNoaaZpiOPLu1MmnZVWLE
+XLsvgiy+NAcXXleMp3IhJKcLe+gD2Oh/3118jQb+YVM2kWuR+El7GwhlR29PR6t
HCTEcTmVA1GgepLxN6PVVpBEuUaGnQHGc7RUsKELLRirCnV2henayFg9ITqAqkJ5
4ssOM9jahXe/Y+ZMjvW9f9FL5IcC4ZlVdTQfnQvKmOjirl0PaghFfrd550NBpOJY
y9XmXfP9zt2UJNkyY8jhYCluqIq8f4RYJNmsF5gprLUUG/6cCSDsss+KckfGVewR
zWrLRK3L1BTAEpvviJOVIjH/eYDRcj2qAKxBdWeLAVEjQ1ceIOnxHSmWGALhTmpu
rAHrUNod9fecVS5deMLnDhgZc2uN8NbwtG9YnnrdQ8QdM3gojwK58MYCinmMeoR0
P4WQH1LuA7wIZqnpIW2p0k8wXUILrKDjx/mF5ZMoLR02ypSwmeMz7JqXXD2vWrec
qu3mmEwrJySg84sSSe1NIlIspFJlQ0K5p110BDdpLvH0eL+D38SibiK7yf3fXsch
FBo/9N7WaRypBuqjAVUiyKnyBmYp+m9dERcfeI4dV/SlzZ0IEa60RoBIXsJvmhUD
3EltGUo/BNF2bxDUMx0JgfTRBuJhYFDvKdRjNKaWA7bRY2TBUjhbvCOUOp7l6my+
Sp+g26p9mrTqO6DbLE8z+qHdhMjjFtQwN4PHvzF8VbRgmZkoZk/2Bcp54NYN4kKF
JeBqyD8DPdMWV7Exwvng6JeS7cl9XspdbaTgGqsnUNTTVFFSUkPB/ULb7nAv25KA
v3GpH2275Ifqw37pe2d/6Xvp30mG/sQVF8uKL7h21dUDJp8qWyIKzIR5IJB6oKZN
t7LRYvp55IqBGbdziGpW/qmCVGnOtQ6ei6If2u0reYw6qVJtJPkXdjR50wRnycOM
JdDTk1ChUk8uw7Tpi7DcFIP93LwRNMB9Nq+RNu5TaypOy1basLCIXD2whgLjTkMV
XexSM21FNVWZeXZmqRhpSA5RG1NZsbOYNfkNRUb0+HiqRsS7nuJg92vd/s00PIv2
WN3jz0MG45WOjG4GFAV0n4XHdeWFmD9CEu83LRrj9MSeETTMgYXLRFBb073SEByB
yNmE/2+CnBp/iNNYtsMFIG7PVM3eH//VZcW6Akd0ZTPuXOP/9/w/uA8Ai5rj5Y92
9fH54gQcgOZAgnCIAkoKZxFeJwelyNU/Crb0acGPvv5TIJHifH8QM0HpmdjmfSWT
zZL8sMmJXhv96U9Hn560HVg0CtiTbIBxbld44nXHerNL67a9fvrQoDM9b+9iNIk5
zOew0MJPnqbESxag8bQsqnkuZx57ZQkMK4hiRWS6vyMDgZHpVCxyRE7nI+V66qWc
Pvg/jvp9OuVZHYulkTnbxA5Utm6ISLESCutaNUvTv9eg7CjaOfQO74yNNwSybwtG
o8byqghr22LrCd27OwENbGHuLkKfs5UmwIp2vrXfCnaVjpDwFdmH5BKJqXiXCdIa
bRWm2iDrchxttDFVoa5kD8rGrCptNnMlwuKewLa83ieOT6E/J+RSZa6Bi6+vvqaS
UXKSNGdTMH5lhsdJACr11cvmYQ2ZfuIXJ9w6xth05a2BB9JhcDzk/AzSsMWozJNp
ZZew1FHlSXBmSHxTBboDc9/mitok7Kqx8Naok5Pr7hwZGJx+14kZ6UTIpPuI9aEC
Tka1Xa4Kz9GzMZ/FnhL9C/J5J4CYnVt/R/qpGKBnRenrbIZub8+bG2kkEKjKejE6
ydGhGFoYNymA83S2jeMdKrjck+62ApCqEvHr6sRBkUNbUsmeLFY+gcPb7jFEJJH2
/fLi7tjNcskHdraSt27TySKm50OTX/Ga3ME3M/+UR1ttMhmMhFEXkDDDMBhDta41
vZw+dIh/yQZqtUDW2cyZsrncb2vUxIRInjd0twtwk+75dcEvxRRtm5D5sXzktFuR
axdZy1E2FY97AYv+4SOWG6g9SNLlPyfZCWS7AU+Qbdi/FcPhUW09aRICDc9Atlom
A3r+b2O8nAVfj2D7dguMEvt6ZyGaPuC+HRq+AjzwwTa8eSTg5NlnKwpYLQluChkQ
E+vFNkIio2RdwyRyi6Lr50DOaaFRIrCH9P2IQDSicvzlHpWtnwklUJgrCjaDmOxo
FHqPMDgqNi/uoIn216lvavqSB/t4aBAvS7fYgX1ddNw1D972POLNJrHpBcO4M/il
LGLgVIAVJ4tfy4oGx8pTFWfNdE598X40IFCgsPuOk6ukbl30CZA0/RRgfA/esVL3
+D6i+xdqS7i0pceW5KdldL7UqKpRychKvmQ9gVSlnrQFMhVQ7i4Xfsbud3yhQugZ
8aZh1XLmalMdOkRgQuNyvWm5LJR9UPBPheuL1/pXVCJeml4SrK/NAS6pKwlQhJID
H+GZeJje7gxSOWKdD7a0qsJTrZNHi13e53xO0rcPM0argr3+dyK/G72SWIDuQNEF
QgRIqf0+FTvZ4ZYOY9XBKsIUtuqHF8f7UmVyelUGytelVnE0wNlXh9bBidYE97bF
qFcp8S1NYfg2hW6Esgl8U9bJwfYlEnnFmZcS9GxZy4MpnFKWyVqfO5sq9n9k48/B
e9gJ2V5m7m6i8INmPBBpDnmHWWwVAa28N5TJbXPhGzcuKKyYNAj6moPtkPvduHsD
qcxLf8EBzNcShyvVdGjBXkKW4V5EL0pojd0+WvXC0tFq5l83c0hUHDJYkf8vPCH0
Bu8kD/wv3WmpQhV3X0FxW3V6tkegXJhem4Uaq6EMG2g0sJGowBK9g2e2jpoyTrDd
yzYn2pp2uWsVnwiaCCN679XoFzuD8yxiN+4XP0DjNNvEzLfyJ5W0fab3A/vWdnxX
HM0B8LeZQnaOMTg/Dy1RLAx5gomWezJQJdbC3QZg+KIiNl7YNB7V1S6781y7KMXu
hS8c+1dQBaor2+PkcY+NvV2z5NCce22BAs7+15iyIaJflgLxT/jnem07L5fzMBjG
FPAxieAw0uyQM0E6Tueu0Ut6JE6zz/cOKKICuCwJEtKk3EhwYrfNAKl+pl78u3TU
uB/l7agJG2GWHXneaROms5i5M9Jxqf3B16yX9AKyTpY9NAcz9BBbDf/pf54LPwhs
JSPWXzmGMaye1A9gyPz3H++u7o/Lb2lPa1PyEGBSKzZk0DInQOGVmca40XTAPpOC
01KnRmNzy+KHpxCwow/xzMTElY5kt8u3qBrJMhNODem/rvj42qR4d4NIjuoR3FBQ
/YgEhPlkuUU+QjC6EzqvOx9x60241dtv2TkZm2esu2inaTH1KH1F1TrVH5zZtmYK
Tq70tFSPynp7uW+8JWc1TrIkkQh2eBMRtSOUP0l0uFqccMmBvUYQJHeJMcfLKs1z
01jmS2HmffyC+S0UNfEeLjjGMDsPBRiKyWdIHVs7h3CYXgBw3oHsLUMF4/xnp3DG
iHPsfOQzzog4Ah65cQqKhjyjxfaJDwWFFbaQZGyXPpubqgY958bU9y1xSQoNi68X
WQyVmEPYPZsezWUK+HOIdHeKtSe1XRMbHPzJmNXCgMTQMKJ5StqvOsToVpp2DEjQ
zjQDqTV8C4ECS0d9tGeB3j1Ji1hgJ20zc3DQ6JaKey1p5YYYUh99TgQvXkuSdD08
JqbI4812Tuwf0A1P3bVaHa9v8hNEEKHRoDcZDQfEWQ6fvS/U1SkvxHPGl0tINaDG
Y0gJrtCpUdy39RbgjYWUun0yFcDG/uAYCV/0c6khawpi0zkeMlESP5ZChwmIvTvN
kUYhQI7UtA3aqoc64e3Im8pG5dyRWfGEt1gZA6IAfiTzfLo1fjrxX52JAKAMCDVi
YGlclobYiWlFpr8hv36nW+ZhOZpTRpnSQT7rATa7pevMfbg6N5P9+diqviPDW8m1
/zu/JVXMLqa7VDmvas7D2Axxk2LdHdTrK3WpRXD2//wRZiEwmlWAhI3SGepibsPx
6XX9/ncLcrqDzV5MjrU0x7C1z8bLkAlHARElIQ4ln2cWvUXXp+LzFu9dDqvmJbr5
jwaYsGwpTfeAXgnJ4mpww308e8XYvaDbGdhl00cnPF1vClABi7VJKYrJz3hRGqeo
UZfpp4KHKy57wUxsTAfP+yk2FQfEQjO6CgZaPYAFiBhED7sFtW2fqlkm5tnKzxzK
FMG/fv0iJk4hoLxAQd6D4iP0QZqSceF/ugg4bu100/G3pv9yaQkRWEFoEMEK+1P8
D9yN6axUX57Uef7yprjEcyohnBZlO/1C/oWmd3wYwrrEJ4luz1VcxLhLFu5zdPn3
AvmEIRtxW3P+O8OW8auvxjImbrbbSwQQcU7p9AXBi6K4L35UGg1+BUf4XA6IY+e3
ePLQaJPecQn52Osav+KlkK9q05IJ768XBph7U1JSnZ7oMjUN3uATkQOsFwjo3MgD
lnV79nfhrBx1vC7H8hSmxI8tqE2kykPKjnNnGI6yWK1DhjLx167S1gDu5Rd6UfJi
zOI7WorD5dPAew4cEACLLEjBMqPtXEBDVcia64vJwJd5q9O+TdCGp7NTeBxd8EcY
+vrEeTE5DFWHAzEWN4Vhw4xP++MGGVPUUdgnjP/Dpcxb8BPrmCf8zNmYRavFiyYi
jtp7qYuoeqCeIFlSHxqxPmZmUxMf1AzWQ+//ujVQFhd5YizLeQ7qkb9O/QmS1ehB
Xskt9Bo9BdMK1EznW8zws4/IgqpDkBacRlFvA4+//6qq5q5enEFzl1w5QRSivzBW
aXcF2+pmBQROJcou6jCL7s6Kwan1voZ+2NVg7mNBN+2DBYBVwMofqiTtuDeWssfF
OfBtYH0HU8wqb3TxlQM/FXFi7ZNpokmxftWZ5eDBGOJ4ndbR9xXzb3ikK6twJMsh
FN0TPejU7QdZ4beWMmTvgIzEVO777+Xrmpw+aKdQzj/OTkT2DVkZWh24KQzAIKXZ
eIp2WsrKWHHZiIVqJAI6F6XG5lPeSpoSbCR0M8yNSk5yilZPUkg7ZPU0VoQwa+Ad
y9pOorZ1neWzjJsvz0SOSVod+ZwI9O7hOBzYW5DUBqqOZZE+Vgrt0mTvLpYMKup6
HbZZ2b+9RtPNLBgZJnksUouOgYIS2fgmSPs/AGzN0wMUbFFp9e1tf4B8kc6YLV1m
+DT+i6bl6yLC57LxCFX/i7V3FD4udpIEwNHzqHlvD0hbd3RVEaYTDAatQ2ISNZYX
+XpWu9eWt2oqPl7Wfq9Ud0fBlqMyDCH2/fYCHkBij2uNLWtEJ6DCO04UBysrg5Un
3YLNokJJSXRICATqB4NK2fFEHX2//pe97U5Wcn5V9nbbXITBgKKVbNkoM1D3f+Mt
E1cxOvGijCxAnQbJ2Pp57txr1XdFklEFcovuxSB3WDOWgA7SSqBQ2vFMD4GGaiOw
lluwfDFV3aZe9A/06ablLx0uk+4KzZp1Yg8V+poiqinpPtiA07Y1a3hqBtkZioPM
8JVgUjl7ZBj0d3BJOxyos2MIxcK0j5krM1VrLRZzYDG39l3ab+oUrECVnwtv6XON
CYpj2niEVP/FSd3K8MVs4NbhdKgzZtMCvfcDuT5OS9iD42ZY3VJjSyD03E8P/DVt
kZCQoM11i9KfogkGuNAdZjy/DF1Nc8rImcUxfE0Noe9hsAHEtlzwHQUPaZ5azjFL
P3y5xwQckNJQTQIcF+bJiSI9OTQuu+Dse05HhCRc2A9GxdvQWQ4YeeO/HJoPM7o2
td4Nimjx95ldFcxZjOVXoqz7ppqHTz8WPrmG0Mjv3kyQj/zlSdDw8BzK8TEIMuX+
YKKmIZK1E3AhuGgy7bkP1yTjRgbgR5COh9S+K0PQMteFAdPgIjDCY1Dwu2JLuMre
/cjIKYCA/KrINGuVrDXD/dWNuWezqykU4rhqq8Q0Cc448P7JHzaXAoSJYcbzQgix
cCKe1QefZBVOuAxehXhEAALtZoh7HIDkOli30PLnxH9fe6ZP+O9vHmf5U7/uGSEw
DpwwqGlUleXMI4wlp96s6ZKx4Tmg01gn4IlVB9vGjAyJQtYlTVOKcoCiBq80Mi4I
1AIhGOP7yUB6ZQotmo8cuRLBRCXKV/d/KM3bbMSKW0TG31l12yxUgNl2YIvZFur3
Ph4JPgIbTwWZTuXEYAYZvCpe4Miamylz+8VF6H9IXeo1+Fr0VFVJFZ6iTWiNyczM
yvO/RmLnj8B6kBqVM6l2hVzylcBaBpwKDsfzyV8crTphGP5Au+l+XTwpsicHZS6u
BDrYwXYUZFdQmEOOeB+NiIRmJUInBFjKtAbOAx/N9+XrsDlYnjY0sJ1jJ77/5tlr
bixP/AHX8Q7pBpuviinOpQfoY6tmvhSs8NTxkyPk1B84Xh2ZXR4MOHDHGB1SRr/q
9YXPi8mL/HBeUTjjBYObuINjgtIPnbh+JukKPn/1RNLPDjouZgKW8Yh46zTyghEI
mwwaKPrpk+lcW5GJnkb76AE0uf8cBxtckx/nVSuj5pBGrUumAA+YKUGqohzB+AjQ
KYqE6ewDYA/Yr5f9Kfkoc/lmDHJptBoJ+Kszd5NA+x1HNX9ffMw8rQBQ6Bm7LH8P
O9cpaR09lmuxiJHtRxF7tldf57CXh8aRbSb3N7qFVuEo4vcm9KIMIG72grt8JD0K
cY5ZF689QjfvgiK585y2GYQg95GQzmE2PtUMy3nCUNEoaBXXerP2jgsokNBiP57/
VzdRNZ6Tr98bnvY3bM9OvoB+kGdwsS3M7fW3BUzupdCJPBaka3dmUkbWzdqSb9JW
Gyz9MQ/H+lxUMKV3TrYEWai6JZ9yrPg3KgA7LkE2N8qcvPacNiofB1/zPi2EveVM
gjessXocH/7vjKyIWzGhTRAggdrPVvnBZ9k+rgbOdlcd/mDLZnckiD9HIjEynEVl
2JZaut7FDi1FKhyVeClCGauD+z8ipt0G2ZBw6e7JqK/vnVenZGLGPRcalz+fBSmc
Ki38M8x/ERmk8iV4Yn1LIuwL52nuzoxJwsBa2QKsqTy88gfSwH1ShSeFOQz0j8oz
zTBOnezzW8+VuiE5iiK6t3jtCJClPPBWsx0eu5Aai7TVGgzy9iCHGuCSkP33J/UM
5le7AjOfaNp0UJiG+vZ0UdI538Z8m6Ri3Dj9PtPQuYh0jP2bMNBQ640f9pa7lq06
J9A9c4xFnIe7NQk7/26gxypcejYBxwi47Eh763MrorrfMut4BKuM1hx2kP7dSNn0
1u2aLS3ak7SyVqNwrQGwNc5EAxCbSUpydUSSUdR9s9CzjBhWttcRVWboGI0ejXdS
AzXx3uptJQtBmCEGNxLoU0RlH325+ug0qf2BYDs/Wn9dq6ZABmu3fy6kfIGbW0kX
8cE9fJ/g8cAxD1TlmGtRnH21vQxW+TlZ+x/aOPCZt0xDB33Oip3vmAp8gxHoWxx0
JO3+knqecBF/uwcuuUd5mSTebG6oqHtDFt+36/Y4UI0Fo9vvbJS6/DkKvGfXXptb
imZo7a3ts8kXosS7vDUFXv7mUaM0s5DPk2M1DZpJDguXjlw9f/hL/BwdZ3uHoj1H
7Zoduxoog4EdwHd8pmSHBS1jKqhOo1ADRF2gPUTLRQCifcSUVpaWGEEj1WhZcFCc
EAKn52LXyfGdoQbGsyBNoMSlbRnKaekjnmnj/FybnWbp7KDQpkWtACcspe1NiTWM
6TnLl3HQ3MDodKyyy1dFRF3P2IRrjCYMK4/t4WOgL+0Or9cMlamldbZcl+hpHAXf
T1RC3jhrut5f0NssBKSMNXY/ftxKyvFYm71nuOt1+GBeTIA8mtfn/YUHoLnM0qK8
VQB7XyMiRIk/859CzE3HknNl6Zozak/Iv34YA92ptrdRr40B1XO2SB51aajyoHLJ
lB4qxjHY7x5HA4rYHIPbQBsT9Ix9oHuaNJRGPkAAdeA/6gME0t0a+9U69yCrgfgF
rqu23R7EI/1t3rNmU0pO1qoWGeN6kJgpDMPR3HBt0WgncBGASbgvZdAxhIBZKMDn
VKt7A4MURr/zAOSQFpjIVoXAaKApQJBny6GHE38XpNYxf49wOiRov6eZpcK33149
lMdZ9DbdZFk74Fc/qldNBGFk3uW6OGxA59UOMU3Qq+x3s9vHn9QJEbgtaPHWI04e
cBYha8IRaYHobuB1GUWqB7RsJE0zSboNA2t36a1V2Ll1u+wy5ALdAHMdjnt7lE1d
ndZM3D+1Yh41FZryDV1XZhr8ReQlMGMtgUQvPS6LVaGRnNPal9AQBqPkMzpDidXj
Vsmbeho7sE4tVACtpqfkccdZhBOuySpsfki7T6hHhtBdkT+CK+BPdidNpQE25TdW
QDnB9fFOCn3i66cjTT5TqKmw8JwykFuWiLbTGFkGR8w+08Jocwt9jqIb8RWaZeIj
W7CmYK3NMhVBKiwX8ENIjZMgcJRWaYDDF2ndISVw+APkxqxiGYaBoGCdnm99CBLh
+cA11v3Vex0YuDkKG5ytT0IOeB6DsCbh/XpPgRqrDRLUaEm14IPi4r7Okb4HVeJT
KFYCwd/Pp+H2pJ21IYvq4Y3xc2WrqaTvlkbJhb/W/hWH6rxiO1Lm+WMeLAYavN/X
cOHBmAP5G93IcSRiZDSsFttBLigJgvY12vmgx5tk+aiWaxi/t8NF/GM9pvk8PXch
0x2IANXvO9MsUALpA8M5IQJSFDPwzcA2N+3b8NRQ92XIIfkMG3e3kfTeM5uAv7yy
VQ3+CHRIb+pAqF1C/CFGSUon4nw7PMLGXEHS3rRbVapSxSFwJ4/zxPP/pd7Ei801
VWVBGHkhG+UwCfotLBIxjEqQKJMDeVLtNHi7LqLuaNleMf9AQLtIaW2kW/IUDgqf
kHg5/cZemNyTGd+0bxuS/8296Jg2fUytX2sJZl9QJ4sicDW2YKhVjwzuJ+OYd8Hx
Bzo0ZdpVFSR9Sj/V03NWl3FFrZMkhR/ctZff4PM3/LXZwhB92wVvFWEcMk7Re/a7
oVPCz/7gqfez7JvFxuVp/1hreElMDkAUJ0DsCOoHZfpO1eeYU8M57Oy+ERfRmwPS
tCuMdpCY643FS6FALUGx3taGVx6yUo8biUFwSsQpbnnh0HIEQyAwiQI+uwhD53pD
8LZn4Kp7U0zuGfs1yjj9pRZHK6VAJlXW9gWQJtwltRz0fL49TQZt4GYjPuG5X2wj
Nc3N0cHPK/rqQ834CvM65quMPUK2GjqPoB15P9MZ1z+s0htmt840AF5ulpCeISa8
tSQnkSMw5YEzsL2JN6k+1EjNd90RKLffFqQPytJ3lpG3JCxcbvDs1KOFTOmEGhqO
04EbIWUlJnHzDXICVYQ5WmDQ6cQ+Sf4dNWd1ZaYJ5+wOWvOsMluX1aumFxxS8zlz
NyWrHBdfouzhNsRuIVPtjicX+amVCF7Pmap63GWP7AA9PCN2Z9ZAz65JC1i0ex1Q
p8zcFx6miKqc+d4kQJdVOf7N8jFOeXe0iiC0XgV35fwKDlkYM9ovKim0gEE/1uwR
J9rijPytsi2LIz7vAzNTGG7ZwKLosw5JMM8Sen3XZE/zu18vsiQc7URO7dKfn5FA
JfVeQqEqss/mCNs1/NdR855XypQkYur2j+6H3jaDDhyZCuFmxdPCcQAg39HgOKhb
6pekNgItx1oqp5wOBNuL9jMUgt8XrE9ih//3wJDyHl1+5GSF8yp59Sj9DldCtpsF
jDlJVcHCqZRJ/2TJjE9FLom+2C8+MAhjEFh/uZt3XuULDzC6uye9f1CDngGktDmM
klvmWBrovqvP9tmh6Yx1W53e08Vzh9+mGKhTq1LjFBRsGZbqr/82kovzRANdQR18
q3EvEPxILqADDFxvBrx9wIVPv1qQeNxNXZQ5N0hGrZpSorYaFDVLRsjvHZJF/fuH
hVSHYb1te3WPY1ONWpFLSXR954Er/zv55lX5gG3qIwbzajiqqIoRfcM+uF8ITGoy
RCbirz4150XFRwSitICQ6iCgb6xGgG59mQo8fm4nxtUijcYyCtunGrU/0u+oiwlb
uY0tAnG9YpJi3WfOwZIeUjHMmUoqDffa2M5RRlfNVxvHRhcuNcowWYfw2wk2OoMi
gOk8km2EYDi5HjEyKJN1fJ+MT/vQpWI/T55sH2vcLBpeUPzMHbS9oW7UDfI4o8nZ
Sg4RdUavTWTBilcG0krpx36qL7csu4RbhF/UOIbrNXGumF03A1Jwj+0YbO4WR4nL
Xf1wJkniai6XztW6RegxflA43Y3nihf18+O/794Fea0Hje6EUwSwZEx74rA/b/Ub
rxRshdBcefdiM6nT7ha4qB+Cd/r2eMRnwgYxOYMPuvzAgysyTsPvt3w8UduECDrV
9tVBVMn9J6onJHBJv8ilIXDPOzJkeHay9DIEkVX+g3ApA0cuOovW3IclVCWtxBWZ
N+gjg+rhjIWw+7C4Se4TT7N/RdRh5RvnkNUJ79mD8DQFbMyhgvGrNVvwN/u0YlxM
uPcfwf5CFy2VdHr8IHQmSsejZ09Jy9aVHHA39UsVkboocZFyfqetrcGzy2efJzLI
6fBXspl8njUGEp6hgdy7gFSw0kajl/dbnBIOoBO73kW4lSl0XPMmlNvOcKTztXlY
rVARX8xYrMjY2lBYlPlcpbpJIjdwc0Rlx+ujvfRLhVyE1OpGti/ivXSkN2a/BH8g
IFK1unlFHGA/eyAw4Q+e1tJJz7c3sWhIpEekZKAYJW4WYDYkzzOV0UJp47Li9Sme
l8DB8kOfHMt29azpnHJ0ER9VB8XKrLIUF6/wk+a99mmr0SzDy9/t/uqfV+Of/xJ3
/sB4xU/JyeixJLE5qU/tyY4Gt7rsr3Gh5FZU1CeHKQiaGTxbo1E2v2GssX0ROcHT
pBmtC3ZTP5wS3F/16oHsJNAs+X1vba1QpJGb4pokjBP23QzlHuz5IIIh0uIiKXb6
DdjiayGBecOkh5JUOyUSma+TBeaRdvgPwa4VVcplpcrrArCR6kWPGoY5R7O7KIUD
9yHs823C5AEiFimUrfMJOPaw9OFMY6wVWrjAiQBRFZvzTXfC63IXlVQ/3vqssChK
qAEoRBvYD8XlDBjSOJ3kTVNVz9aXkFj3SMbJNjs9FGJk+8nJoxLCXCWdJymK2vbQ
b9U+JtH/Wz2Uv9YAHVHVJbOT5kdJNlKoq+VY30gGReeCiHqHeNnIjwTh4m7+m6zd
AwWP9bbJxlFpd2K6vGf7ct79ND61QtR+q9qBcZP+uVQZOPmAVK48VypQ+RjZf5R1
NLTuKvaZZIloEbGnoKBpftW9qCwc1RhGEl3AAz137iFhTgvU5Me/IIbv+C5YuHju
hiPl2Pj1a4M8kRHeuRbocTQHo9DRCXR6Cz1u0mrKHN6MYH5sevEk2uHizdiM1yiV
TzxR1ed1wnoJssvW312wOaZN5roG1iewIr6bpS0/SF/5t4whnU3y1eU/2sQFDEzq
3H2zSJl6C3iroVXWZySe6fZijyfeAxtHf1Nr/pbbu9Rx12ivGY7MGFV1G1/F1mB0
iIgJZVfEt91lKUmbrri6GDev+2npn8Qc3bj0hUq/j/zTsD1Qt5uw2jmYaTax5IMl
lZveOMfzakkjh+DVDqI6nGfMNBWFkdZq2/2ndUHO72p6qZW6BtowZ4vREXpxupeJ
UrH+BxLCumhRZLApwpHvLIv98osPPFZ5G1v1aaNExKYw16a5Jw/U6AwgmrJT8SI7
TK+M8y8UURQzwaSIAwz/L1drWW0SIy8qnICAm+ZN8mBOI0gQ9ErZt3pc+ZMG/X2k
uBWI1chdMVq0RC+GiAhBveFjDvQlnuRMRWuCiG1SpcDfHK1SHXOzvW+EQ98LV//T
+9VEKX48RRMYXgr6qPizvZFLC6EsXMZEP+vpX+YLPlgnvt3WWNkjq5s28BIanspw
oBQnpOpYvcZn08X1JVa0XNPDP31SE2qPCiqHuYZgNdY1hEdvoLHdZIkYLCt9tKcL
JyUBCJ0RXvpbkVATImZNprowq52zbp/nnR69d7iflxS8YWLyJ9cRq7vFBdVzsDdu
84SRR0koGWKHj2SGQ9XbM2qwBTXqYuhtRVHO2lO53YpU/nLCZSOId1t32S0q3gTN
zNVFXGj3onDW8F8uT6Uj8JxyhzBSvM005OhgJir6+vgmzf8J1ktxucvEH4gonw0s
jqCD6QkZSXErBR7uTrRjdYGRLwrP7dMyxKL96qz/DtYl5hB2TFAIBS9lMXudg9ZO
gA/TOJZv4x9chy39h5vuje0VFFb2WVogVChHNsDuQ7tyN9rYDnnE1gJ84Po5s0S/
JoZULR6LX/W2+FyXcd0jZFMJ/66lV2xd0gshcQbcI0VNAKldiBCBoNNuWcYY2Ry2
lvLH4J9oLupsiJCpnnKQv6ZGRiAtndAMpZzgQg+auP/k1HNYJlwd5hgI227w2w63
EO9mXo/Y+bQoH9RO+9ZFvJtmjXEV/rtd+Otyvq9+US5j4UTtK6cD5oSRSLtJfIZl
vJpw+zX+KbW0hWHufwqvAumFK4bGT6l799sTn4MPksrXopeOJF2VKynx+1CtYJVw
ip+4pkdyF/ztWTF+pPb9g+lSkkhpZKTbu/riR1DA/HJcmoAAeQt7eylqGguA7thz
HJT8EBL3kXsn7KIYsI3WaglGShmUarCGsBFReBINFW8TkoJoh/hLy7/WVFWGlHdn
KYOuHTSML7M7iGgTmch3ReAQPIcu+3XWKod2qsRmY0jlFaPUmf9e6mt75a9mwCO6
H8NhAwqECs0Qpo204i7+8RUxbLvOdeLxXERakAfW+l1IjmRZEIYaQzN28OKfil0e
32Ad6HyKUIkJvtzgBfGrC9//HANhRAX+jX6JEks1qIA100gG7V1qt+DPuYEFHt0v
nL7N+kKyxJXDEfiQKNNZfLVPV2oT18sEhtUnHeCF8o937HC2nJiaKjCOdKoU/L4M
CfZxMn0KNXDao3S16IRqlYx7X6mAaI+J3OMMdmToOH5Ie77m6dFUdtrkXP0ikpw7
WkjOEPns/EAAipQFcq7gBkKNkAJ5FxD4uB+DVLJ6zieesCM3J8ByHWpwRNyx2nzT
Ct8YBUk+u05vitu2XXX+ZSPMKVJ37mHPuucKChq5YL9pSxjb7iRo6acrFJPM8xFX
1p9DITTleOzDVExearsXcsST4gTqdOkFUHz9xYGDT5e5OLubZ+hHdflJYpb/jbSn
1TCQNhlzmzn6GzjyVCLAl8FLv/D+u/hPZbpJnharICTxuR0PpIWyV3vE3bDe8qRY
dvcbO8VU4Lg/+mEoCKQv11fCXCEUZ5SfE5/FVxW4tfLsTeC6rk5BZYDnqvJC3jP+
snNpAYZifDK+rcycN70utLvFppU9EaciR4CsbadPQ1hK78348NE95p3GA6QEeRwm
tQqLPYqqGZckBqh55RSnar9Gwdp4F+Le+FTkx6alcbsRvt9anfENKGVyxYLsAEUE
VAXperyhtehW0qWjIge2pnr9twCUrKJrqMU1E8kBzZylSBYtXbrx3+j8+wR+cRWh
eUuepkVRjZPDwDONZIWkuyPUaXtnobupVI7D91SThE1fxgLtU+MXckrbr96/zTVC
R5pOzhoVV2Kl1U5syMj2oB7iTG5NnjX2/WTRQj0H2tm97ECeUKYhIn+OiPZRVfsv
4HgqFU9NFRTgqyaqmk60NpptUB18cAsSmbqtgXg0g/DtRrjvUFIPAl5xd2WqRbUH
R5NaDY2QrO+XGvorc4u3FoBGCadcGnIvntKbtPMaK1BkwpevOp6UJIdxv8O3xzTm
EO+m5KS75bsW0Z8HVfT6H7y7/KYG/NbEqnDA3/9dyPk+/DAjCdAD0ByvkYCLHaoF
2m94wcXoAnS6E4dDe1fOWDLjzdojDPAV0E0wR0/aS90JJ6qS/GVLrAJhnppiYdhf
U8M5wIRxfx5W68vQ904e3ka/PAwTRxdjV+C7wLr6Jbk4vLdqUuNyWqx9pDd8AZRf
TCF1M+yGPUCz6E0KhDTBpU0/UpEt9RJKZhtXBTIRX0vFXOe+o6DIBLXx3CGn5iRx
TUG4nw1wZxvhh3Ay8bLVznilHSsuZqZh58xLQSwxG4UBDZhPY1actSomkitANcRJ
ZF7ViLpUZ2BQutxkxv6JJxBaBjeOkax/qHvKZTQNfAeA9ZSX5YXKifCXzW6fgwoE
PJL1BhZogS4MIXdtaOBj/W935qBajx/1TXsXO4DGYUs9V77wrOMyN0FTVW0zquiw
zjlG/8iYGGelGYivzL29J4sNHQYULjFN/JWNEeD3Df4szMqAFNsafXINlchb4cC6
6PYoph18PhZQzR/nbGlg9MwQ2oDa2beqnkH+7sjYGlZzXhDK/UTf7EO5WLXCLMNY
M+dtgENXNPrJGr9/eEyHxVDcbxlWU4AIyAyeE77S3rVEbPo1NDudKDWi5VdWqf+f
k8BnwPWhNy5tZlaJmhQZ325LJqiUBX6I7mvaOvObr2vJxhhJxs2yEUJjRvpjeNAp
PQJJS7lMBJ1NOtB1tQbPrenuekIG0Syj/kCyqDkkglFeEnMSyTsl0L1CsHQhNMs4
eivUPdjiWPhzXOzze4nquXP+DrW4bnRRDLjMLXqdggOzN0WNhlPX/tVlUQ34oc7a
OCuvvNXBbXOTRXHH0ZBbgWDQC0Hwt0Mk4FfMrMyHIsU9OGSh4UGA/OCSTojIePRD
MkjikaiGjjZzwYE2zuf7JtvhfSXQfTMETuxC+Q24viEUqgKimZp4DfOdf3aqP/1r
I9HFJKmFpUDuNfnmC9pVrvuR6uF0dpimBIRSvPb0sCuDClHbrpirvzNe5cE9sR/z
QvGB/RdA59dkU7+r5KEzFM8N2NCVYqD48qfhAQmMflNby3N99WxZP7DM5pbP36Xw
NaaCeB7aXIFaVh1iFADfCb0Vq6k10nl37o0Sbqtw5t23I1ssFIC8Xqjb46BRouij
VWJEQjL7mXiiOZzHgJTHJg+skGE+ApvJv1RmI6reOsDhlYxEtO2odx8xUgdU5url
XbHUGvIj+vpQyDXbhJQoyhT+tJmhLwoSypRRrVI+nx65lngLJCRSPwBcg8bYVU1u
YEJj2XqtZnNaE5jHwleblZEZmsMW5H0Am5pcjxfs4875wvqaKHxeoCM0HpzecBQB
2uLjK1MjAF2JMZhxa+wXf1i6104/wIpJob32cCTlu+2LfSBbSMSsrXhneab9QAPV
ZnT6x5suA+nYShD1yKS8rb61TOH7WFnE4pvX15bgUD9coei/hcq2JtoKebuLNHXt
xD1qHntBhGGJLPLg1rcFzChfdbsJBpk0njySziSpQFOOdl34RPru9sStgZXPPgBe
/6OY5pBXItXChVueJ8OkQ5WUc0Oba5dPm6x9hMBix7c8WMdosfGIHl4U48kkly4X
w+wc2MKqUgqWND2k0/PNV3By0zSYKBEmzRGg96HShrL5GubnGThmDvaViaie7GCH
JgmJ95eD59ky0attudAKMRs5maCi8pQwgGVBUnRLDtiI85P2XrB3uVAJEGWnCkxe
iFN7zk9ttYeqv53d0r9LyN1S984ngEojR23tqtXR5gbX70KPDDiNmGJKfYvJVe3h
6T6mOKfTvQVOp5DtpEKkdufcao0nUO69JOq9t8rNhIN4yqBbcTWKmb2zZzfDOxS3
woDFuAK/PZJA1+Fhwa2yv9dG0V1Cp40k9b67XWFJrydJydt1RiW3caalXFljkD5Z
EnZu+pbKiYFZ/wzMHhM+/o++XgRwLeECQz1xGdO2sppapjeTZgxbyxlCcx1jySvu
fglT0vUcRkc50bBqNcM0P5N584mKO/vCjHwe3xhjCg5SNp/tJ3eV0fsTZkL9dd8k
6bj5BSP2wao3wrajSu29fXaR6A5+YTgzHMBlh1JTQutKM1PmzDStwqf2mA1K15T2
rGuYE++MIctH8NOc0WJqzNr+0eCvZgYyJR+qWoGSHTRH5xfCmQRKUGX0pdlVNSvj
SYrs0JvpB0VBeY3XOBn6uVFxLgYmV03wyv7VAofDAVEKltv6HuP1uNZXUicd5Dk1
CwuvNmIIFWjO0emaxBd8IQdfGqaYdBZFp2JvCuOgvIuc/JTfWuyoAQEwf8kNXMiq
oqh7bNGMaReFJobpVoo80zZN9rfD5gVUfj/ItIVXk/2DnOQQer5HMPk16ZzuRnvX
jg2CjWzmNmuioJHfaL/+PeZSxbucqHnKplFPVdwsl3ChCN5kMLnr6NYnPlxwI9Jc
PwcvC16PO+kNq0pDHh97Ei0T+KRXwCo/FWNWxPCMBJQ8oWugVKWJYhCPWgfoaP+O
Vujf4lPIubsqiR26Xi4wir95leDWdG7ETx/J94Cnn9odClI0E1AltkEn5JCu1VgM
JMnNHpWObAgB1+KfW5ejSBZJANnPQSTGwI811KJuew51sT8zWEmf8wDmhRQIQVpQ
PTomxqDWTi6zVeXSqT+/kT2FZeeKL4Dz9RMfRPN8rPVa81QmgrTe+Q1W4d19oDmR
FlZTOnT0N+UyXe4t6XJBFIuhtGSpOh4RIg67ZQ735fS+tEm3gsVjMEv7cdLFdMS3
S3ckDK2q1Vhpc3jpsM1jhGOyKlISvNsFiqgyW7vGhyijfk5XeZAURQEJ5paOjMJS
x6juAZ0hlRB3ZFnXEjsWD2NPPs66pews9XZAOQzNhGT07c7wSwfgmd/L2Qica/RZ
5pamVFCxDhBN/cskjs7tuis3S0PFxSNpfH9Af5xWxIYXv4tqsXQ4V15AMKcpmYFW
+Z/ggXVzmsHDII39iwysh1Pafx8UHCS/ORCAM88Oy9Cw0QSwJ9rpDS+qA7l4WbTG
CqofSyCuBbWut/3PB0x1bjK5TKH+V2SzdOWnv1gslsOc790HGpz7xkbwiD0G/6fQ
BHSJ+dTQjLDBhkMG1CczkxEQXjzTjXm8y/ZUCQKap/100wMhjEqESxLrtcQA02sv
sUzYrlXlsJoK7tcmGnu9ahXcqm4uHE6/V0PVzxMpLEXlgvrmWjH0pwDVnaYGIKTD
m2DpoDXopJi+COhhnPsDD+ixVDo0Mf6PuFpQS13TEKy281oKCAZ6WFJBBbOwJiP9
ZcK1c+BWQR7G9uLjrmuxwFy+uCVPuQKzKpYQ1X3+xvmP6rXvzv2LuEc/KWm8iGTv
AuXhCM4WahkzMTkI+nakitTC5SCSEa2BNA3KHSEzcXFZrTFAHXnKkLqtAcJV3S4x
YngXAe5JhnMz4BAFDsWQ0rZxRPsT/rUBFqGfqWoV2g0CtXs979mw0dzd/eLPKVDG
JEkDh/+v/rvhdHOqf8sK3DGW7Bsss6SmNPJK2nQoneGTCIgEThxYrGO9ETHHxo8d
veeVU4q2Wu7pmqXZGpPEeLKBqYEe0GvMJtXGLjb06YU69bA/kcoYlMcg94hSkBZU
77l30NcUrgzbCpjpMUEojLG5GeOkTArtqbRblk5NvWSWNl4yvUNh/zfyWB7o4xc4
NS4bYteR0CUxGwF/RUsPxdbZzGnOBQr7ehucKPvm0FWZ3ENSVyRXyyRGQC5vv0Rr
shO5whIY5UnjuPMVLGDIzcle25nFJQZaMNhu/ZMK5JE5SCGOJlPHdo22Ch3PIWZu
Me+T2++C2gZPSOl8uQqVn5TsEMZQUZTUQ0qb8b5M1P6JVfme+gnNprzFKdZ6qax6
9u6ODqhTvtXiUvf8Ifw8tifjMQpMOLWQNwpJ98BxAzeFJvspRUXqEI0YjpwpifDP
zDsRXj+BHRPW4pDyjS/uvweUaD/2+BxpSDK/4FzKWWI0BONsJzMiayj97eT55DvB
htO2x0lJkdjlTD9yJkE0W2lf4RxsC4pHLfPnzQhkWUZj60yDeQmRju0JLDsQIcem
yT3d2OcFwjwFv7/BKUn0ILL7u/ve9OzHBafBjneJsOtUODTukDdAAyULNbgffTKj
Y80t7pz+KKWoTD1Qo+9Z5pfyzjb5/QMykdw7CZElz1rEGWVdZMpbjppDsw4MkSD0
WyNRIC3iGJ+7KMWjTEb7q85xwQQ08e+tpYKd3Lw7jIbFVtQeSVnrJYefqy4LyLM9
aaolBnJisZXdmQYf7INWKyVf83EpgVACMSum1tqNvRUvjRByHEO44osVlZiNYDfi
xS82g1zmIYZs2Mr+vk0gtqLyDjG9kpP44MTAKvbAjBYiUHqR8qRVSPI4Tkl0kuGS
J+xWeBVvbHd/Rd7kwrY+wp04e11VnSodX8LW2Chs2NvXQ4YklUq1H0zZhdWOH4Dp
XpYsAmnK24FV/dVEmjuAoInq8k9FVeZVNuGidP0cP4MMr9FXRGbzVVAmYriTEJjf
9OVOcSsHnfKJ0zo3UEmH0BNLp4K9fa0oE30loOCfOofINZtGBOPih6gI+Nj9cJdj
AJEq7JWgSrHCDllBLNxzCv4N8k9/e+NAg19OYnQtwTBVXLLpimziW4gG0S0ZJu1N
3iN7ddps6nsU8wix11/GtGFpy6AV3KOb1cTD+NF2NaBIIqGkxR1P1ekWc7UE6HDG
ILIGUrSF3mNAStgbbvGqcMkKdoPBohVORdv9VQsarW9sHnHxjYX6fWqgETAu6mvS
VVQpS/kEpjsprw1/4BhoY22OUIhWQUfod/Y6luJa1XFjn4/jYbyrtrknsg25WV6S
1gSaUnK0pR9xw815OnNx+QoRomUmZQiFoFSABXEEBlSvLkiMl+Fwm+zHEu9a576Z
JWjSTMOnowqHcj1X53dOQbdsnKrXEmqDU5+5u3xhI+9anSTrxRGfhZzM8E1I4JlZ
iGo5lgtadyS3PVEIu8rf9hMIWHqM9OCqylsl0wd3GqJGAievrBT+JY5Ai1U/enzm
L2q7GyRw//PCFZ2RRZLCb7Dw4XuAEVEaKFVQzHroz2BPS8bwzAarlgi+L7/GIgf3
nzHeePH8RqYqf++ipGx7/iN2vz2snwwH43KD63vtj9XX8+acn5IzUU9n2gUcJw2f
+wqOHBUV2aGk7x9Chis67oNkhAJR0EW01bqT67VyeMlgQs3W7gA1pzsHTK4sULVX
fhMyP9txNPLfbuClhYicmUsfmkgV/wrRzEthi/lXiohsb0LCNI3tvMoN/jg6ZGiQ
SGhbVNyH5tbgZXBoQlinz5tU9gzH6LdPDNuHWzyFuybKwm0V8lR+2ObTt5nirC5J
+Q/vGC0U+5KNeOlV19FJF2NtuYc/0bpsVhg4XoHVomu19IIh1+i31r3O3WPI/w1V
Pl6wF8ns76jaycss8aN3DnnwD2IGrLgE2FxYXALo/PLpP3vcQTJx4d3UfXBICyOw
P9wE6cxkGSwMxQD08hOn49GfsKEOn3bKGQUCUd3VzjtxjZGMdKSMrU5ytnXq76eB
EIReijWwnJYBYMR3irho5WEczfALVXB08t7LoeeoZtZRgDuZpKbzQD3EYEpToOWf
Wyxq36gseN9z8XjqcuRCiEeUXj61O7O7l1tNC2dggUqtkoaUEK9t0dOGAM/HwNp3
crglY5vJv6HO1EAZ7R4x42HLgHNjec/XtMDTOQN7xAvDhYxt4ENvuzyAzf9wZN1j
GI62S3MezE2c/3b0YCKO4LSM8ScGxPPiPYJtiGPXvJem7rrJPwzUYeK9RerZovtx
Wr/BVamUhYnBlc4oGo2ou6IrnelODBRyt0rOecow/PS3CEWaus0Gam1SoE3U+UL1
wxvbuiVnFBXEFaNjYcIdGP6lIsSOHi0yhwHASrGE5QlBfBD1JGGqJT0zMxl+50zv
g/xVhUyCLFXw9yecNX/krH/F47Yie6hqAsFfF172w7bB5Fty92+G0OYGIxJzoKSW
ZXb3eOep+SuTAPWnfPpk+wO+mqUFoYvR21pHQuZiUQ6bpPulJRiKPdzvE0MUXB5P
KPGXB2lXzOTcI9SkpR3J+oOK/g+6KdT7exFMNF1o6vzhqZPmoTK8j/zb/espn0rG
CTz/Faw3BmIL21CFjEGha6g9Jz7ZC+SQmMSjiKsWWHXyMsv0caZcaGAyVfxzRTEp
6leY2sRaU8q5pDF3DR5QFfXKmhqilwm4O74qepaAAmEpNLYYJxaSX7vdUN59xHJN
WmL+4jAtj8KMyGiSdgRE34VEUSOikD2+IwaRntbpmqvO7y9LesZzaRN3WmmB6NwF
8z+7cJjbz0ZU6T2A3Sgi7ZWgcEx9ccM3w4WQ7L9tQjIea0KNB19FXrtoCRc8a502
so/qh1Jxgjb9ci6Cb2Ewl5099JOkwyg4RFyMTxfkhaSLf1CjprqD4fbv8tvAoIrW
ZIsOBgZmqnaFaTozLAZ2u38fSNWoRunNSAj9fINtfW1P234JqR/P+ks7DDCtg8R4
CReKm4R3mV6I8xNfivJVG5i9bak5GghiakbcC3VZliqUxc2MCHmyV552xumX2KgH
Wyn1D98iMkvBEeJ1pZpfvROD2I6E9PFJl2ESlrT8CHDJJuVhg8KJqfC7imYXkPn9
PaOyKJdsxG44pqIHgzshbzgzwTItx2zHkjZhZGRwpwNs+0jxu+WYf7jQ8CqKDXdL
ayZxxhoxpzhhD3f/aPN07kxglUrILvrl8OX4QiJ8oPpjoU8RI+Re53h7pmGd8A0Y
alvi3SCiI25oDbox4G71nQwfY9qQM+XvW9rs1lwVp59lkQhSoYSm88M39qAeizcO
MVKg46uiNKu7lQvilkuziBnDSdqHB86qDCifaFXMME7hXyiAN/ijpS2HC8bTpu+H
SsgOGq7c01PqOoEuGgHSUrYJnHqn/O2ocMmfFtCpNleb++frmzUcO8yyJ++Lv21h
+DnJcNT7QrMgZxRy7AdjZMmiCrP3RnwM+z9UGjI5rjQpsWig5OF7DbdFB65mU6BA
a5ni78C9O5FIK+Q+U7zvff/RmDoOJKfFAKsUj/HY9shQ5XuH4tw8pbEbqbCyyljI
34hrqsKK8k2NtYGJS32i+GThAuZjz9+Bm1XDgRpc7gVCrEMjML1MRmq458o7Gw3b
ORD+D0XgHaVjUQLO9DOV61YTYG+9kD8lgfZUoSH7aZ5phFEACkVsaxN1n0aGS3si
p4jY1+irF0dIEqpwvZef00wD7UzloFYfV39xeRFpNaH2WlZIhe2Oq8OHyMUPVR5+
dbA1nNBlYL4RU8BuPp2rgqB+7GJ/mmYbdUn8/2brLQDy/MwBBGxyVMibsrwR3L9K
Fo9FYFNJvYEt92hO3LyzGKYNyDjQzmlUqbUEaCzvrg1Pza7JaJvhtD/OJnimoifE
S9mYk8t9CsO3FgtdqdadGAevoow7bw6FC9In8IC3bEemmoZcTykvr+kIeVGZuzK/
a2lW6onk9cIqS9uGaiFmoZ8ZP31EkzmL3gs6Lh+ol0ZIg3VY24wdy4UfuNxpxfgt
SHLsIIIACfIeX6wLQy7jWQpW7YcY67LCqEVRBeUPuGDpzdlG0eTOUFpCp4v4XHn1
rVjvzG/TBFdR/Tl2iOXoOGEve+iLO83FiYyc+NcR8lWoP9oUXkW3Gk8kYl13psnR
w3Z2Klun/NURnILrlsAHQEhGHz8tNwAr0ZYmEe4krFglxf665O3LlSoZezfhWrgF
UzVfIvMH8nkJt813bsC7D2bw2KxE1Cvbi618EykbQc5YWB2+Ritfadb8H6GUomWf
cv8VUfGUD9shAs2vtaMSZXaQv6eD8xakYbsJ0S172TOQgq8P3+PQ9HvkSTsjq/7V
AHqlOX1UKD+7oO8+F0UkVvhhmVLkPYoy27kfo0hIKBO9IJnwdSaM6y8r5B9I2Vf8
WjJvIz+O3fbobp6EeBFDanV0tyUEikNIdkoGSgJLanF1v2651g2ASvpOgwWtf5gv
KftprIt9jOe/xoimX7Rsxsv0PGWULXN4ZsDLA10+H7+ELiATD6lJhuRH2a5wVoDh
z731OO2i1ihXo+GIKWw1x45I/eMay/FBzCk3+XWbpzfapYG2Au2s6T03ZgRlRbZ/
Qv+kojF77wD2eqVNC6wKGM9f8T+hdQ08nEWkeiPaA2LRVsns+J4hmdhZ4qYdS1uS
yNiEKEQjNOo4YJeUPDEGvc4zE2sRJczp6/jieCgnRVgNrJDuweS7/eNYX02odH7x
A0G43wfNa+PGJZd9DsM1Vcsn6cmsqTzZ4VgLepd52TFrPLqdJ1fCSiRKUqAJszaW
lT6jHnalX0aOxhHViLpDj6xXIdz5PTRJOnpZy6AEkmI4qfXPdKMRMXxoXW0TRVT9
XKiEgcxBVsvwyl69O/djc4MHer4FPCLjD7aCotKQ5P9n3dEomS3KqCGDI2KfWaIT
N5RQ/9FDoN2w8Q+A1mfaTbSPl2TEHiStd03UGr6UXnJ+EWHXu4Fz4DkKmL22AZ0G
LZSAdywL/8vrSKvEHwDHETsC5OahQ3gR0BntgtMczoevQo52FJqRw0kI0ImSTHl3
HDZKny2zT6GPzn5dE3kzHUndrjr1T0HO3KvA0uF7lwBv06sHv/z4PbZAmPrNKfHx
PJe/yBIuAcX4AvB5IJtAkDjBLeix2uDbinKrp93R8eftR1nv9GUXjFKkTvqOJbnc
pCgISufcf6+QcAY7oCFOZQYz/FnWq1rYl51XfSK8t8RaBvkkw0LMJnQmtqnaIIr0
r5dPdfDFp2+hG8FPiUaQbDbLsby3yAi5vyeMZBVhlmyrOMbHRo5ykNufKqTZK+Xo
F+GBNJze175ZpTWvgpDYAG4FyhAyWRg5DVgj3D446EhCs19N5/w0knB06RFHr1DR
YSTlyNr300MkSWa7LhD441mekN7Drg0UBuDc9DeRq7pa4p2Dn3czkcRwbJWMR92I
lP3QzeDvc8libhhlnG0yyU3DxTNm8G/RJQrHyo6gWXsY3Y399R80vzMNx+ud84S1
w2s9dpYdRD05bCpj4hJV1iapgVJcNytrzd64KwmQKkhCjAcK7xsrswMSzAwAWln8
arysilNM+dJom6qBa4/wFA0lPexyZNyNh0Py2lpe2a3TuykTYIV2rtL7IanXYIn6
3byuXdZRHuq7mY13K002BXHo3E8fXqE84zSTxKXkzd8Gs2QQ61Fgk65JD4NNhuow
Mbt3jRF1eeF+K8OoVRpj+AVx6pe0zL/jUo7Vh5BqR6EvFiUdaS4WTtEtfsOQ4G8J
DD8q4CI2xTRZE9vPlqyip8DYF8zAUN3Xz5e3cn8nBch773o4WtVi3i1MWHIWE8sf
dkLgwEZVUfcFtFHLh+7fGcbPgZPTArGIS8oXo9uKLT9YoVVfAUA80dbcHdsuT1L5
kZSnB4f2nTg9mU8zTJ2HrkVYp/ibo//DucPZvcHIcOyE3aKxaFDfvdJiLLr1TuOm
vpgQthEmqyhm2rve0b0FC3uUxQXAzU/LJb5ShTWooEkGRS12avJDAsrmc/oH9+rv
XKc7TLeZhgYJiN3VD3SihbBNQfrQipYotXHQBC3eVaHnURmBJK+e9XajlCNGoY8R
M4ej8ohM34qGN61VSSOggEqdnGdDLM5uxLZjlk5Qv7EvmKByDrZ+l6qL1OB9HGdQ
YvxfkVIhukOMCeVvk7zejn8HkzZxTFCqYeEUT+3rCek8xUxE1TXJpkKYJOTg0ZXW
c5DMYdi9Dc9qORqENsqE6eGNkWFzCCAu3/9d7lY6eqjJrsGlqwTiU+K//22eiS/U
f3ERPUP14iG7KEkn8D/xhey45hgzpePjD5KHnrD9K0Kfm3ngGAG8ghQOJjMV3Tek
+XxcLqjYgkvasUQ2BJ5PZhbtFg0gCwnJKLpfyaHMyZDf3Ewbt7mJ2dGyKrENuUZT
wk5twkJFtMEaHejAvQxRCizc8SmkBHrhh3FMVHAAiJKYsv3QoWRODIagS0nkZDyo
CEnaNM9bVZEoqofEUZKvg+gNzlbFGKZ8K+8+R/XbeDLMsj8KPXSjkishgDkbGNSU
UKMyGljgY8icI0KRniS2UoyPcV4l9jia2tcqoLg8BFHbmXBgdVeozv9w0rHA8B5n
fzea9+xDnywqn3KYgncaI2MhGASHS/BKjccC4GOPXjqJj42SBujyT9iXXTXj6nUP
skwM30e7fumKg1huxtPO7Gth06ZuaQ7WuKvvMpDU7IqBX8yhgMZoRXpFmn3uWXac
gLsphMW+UmsWK6qOpa8g5EVBgBs0StW1sN2vPgqoRvX3iilPzsGIt8BAxAH+uVxC
9bdJk6+FZN+vc7nCKLvYaqoFTpoPvYC9KuKb99pHcBE+1INH3DDw4nnKTEGNSqJE
NdJjKZaY0ytGXXioH2e9M9dlbhfCvCqzXtKINyzqhZoinGFh2dgToQO9vdrl1d1W
cLbGL2LudpA8tZg8WZNGwwKvAfonIg4LrfssCnRiokDAnv5JG28FYwHzrSCE/Wwr
osbm721MtImYWgpZdwzRBKg5Mv4p9Ck62srRLp2GZQDSGNsNSAtOF2YDDVQ0FTjl
Lq3qqrdheCIS1py/KcbppKquIY/qcP00McTgMGGl/Vrsw/031d+PyqN3oPiWMPjK
sdHiJhsHFqL+GhT6BghtpLkwtYIQLtxR4KxbXnbqDo+9Gsxhj2XmxLd3cqfLrcpL
rZfulejQtBc2SttX482Flvm7DyJPyiihvxivFwYxCqREWHUiy+KHi+zj6FqdsbAT
McPB19of5M6gXnY5e8y45S67o8kEIGxt74GfmaF9CmGgpDyFwPKiNh7Qd09CcWQ8
7nD9hk68wcrUrKiMAAlnZq/vVlQY7X9JLlJ01TgMdef+VTtHJ17Sm+5hgHodtbz2
xAkIL97FHczHCY7mL2FvP2ZD8toFvRlO+MN3hNlfOn4mO3fwInEVIygU2mNniWsT
09cTUomTTGXQHiQTW8SbISN3glKkA8m0zqwKPdrFnTaIk/13NOsKNOwC7i4sxgy5
4ZwlREsBBBSZrnILeot0pR+c8ScfP4/AxUJWUytrJj+2JdtwOsZsijs/3TGGI8BG
5lrILOG6vq3cjKndytgfVTW+lhM2NQ3Qzd3zBy3xCram5bJgBVc+GvGRQVzwh68l
/OD2cuJEgUGHAi9LLEFL88PhaGfTs+3b6uVGkevvqPOaOWc2odKQws/abiIxXzlH
/w//jloCdNHG6K37SkRs1QXQn2V3+29QpidB6PMobhCfn2ztQkY6RZc/vpSfHZmZ
fn5HDEqfmY1fUe9NL2KK4IWUGtZs5mtwOOvmbyYRJMEH6lv+IOtFOGuoSqwcpAAI
iUgmgzhg/OPPn0sn3VIRG7jjGqALjp9e3gE8dOA5NnLZ6SsegktwX8xVEQWPx2Q2
+vG8nJl0TwEwXBPvjGBrnrQLkdlzlmXNJltkYRgiced6QHuu1V5siM5F+xlIv3az
XZMg7m9JsvbN6zKG8hNvTxVRo7WctkvEgwsA8WVYwW9iuDeAkO5KEAu6jD+diBWn
SbsUJiJH7PSlc0pkrge5PSTizuSi0lqLMFFgUkoVptkDrbcf7zNPu4g9E1eK5uoi
qx2fF89R6/FUdQ+77GRq4MNksOzUeE+DwRozLHfFGsTOakx4ZlPYrmdWwQM8JhDQ
3/1XmcyFU/E7i0TlW/ZcfMHbMJgnF26eFTdo97DUVmiSZ6/ZzeFYdGfuxRzu4REr
HzZSyy6qhPMIt8Lz0f38UJ8J+XAp0Sq/SMuvcqJKd3gjsZ4UfEmneh9/SuE7iURL
GJbRhiai4myizw+WWi8QtZnkRq9wvmRkRdctf87UAka/BHumbyf4CUWXigM4dkpI
9U7LjTColDXilzIsVAYsyK4Xo6LS/Dhs0jo0vLq8tRL4mqLUlRUy2yblvQNHRQtI
0ULTbiMccC47TLb+oa+OiL7bMREiceowZZD9kRzXOueCfoXuVGBDoyLNHY1EDqTr
SWOCdzBODaC3DQwiATLGZnB+3aPnFKlM5sasw8ZkyiutuY/GPbknQFNL2N1PUjPy
G0XXXF674pogbeKGdX5LVUFqq1CoAPWyQnWDhC8pZSstu+1qWAN44mdRWbckcACb
HkVqkb6o51LJQJczI0OMhn5IQqGtAM4kqogRWMQ9ZsOU0YFmmE2pV0moG0NSS/dZ
33gSUmJeCZtwlzuS/SyJQDUCyYGqUzsPUyKAc9M+qhzyPDFPSShsBheew3kflmlN
PLFdV/oI0+mSJ67jt+kPLTzCInyztlFy1fUh0YZR9OV9X+Nipa/P3WfNrqzuGdKT
ee04tKKd8oplcGUCfSstbywVN6crb7tYwA9RlvBSAYlKQOzXrYGRjTGVAx4CCWFo
3azdJmBT+zwRVsg5tMOBLQTkVZZaLUCQ0YJhImXPOtIzQgyC5jdx22GGUtw/0DB5
98v6/f7p4nThudAuoLoqfAUf7oZDwzfy64ic6/5Jr2kP92+2bx8Uht5t9YChJbrA
5WGcjsJm+b4sB6/f3IRf2a73CFOWZfT16K9jUpTJQ6Dcm8irIVwdkybK9u7KpuCM
NZ/JmgeZDoH3hFJtlltwctxhE/Bnva2lndx3kvJ9MQLji6L+W/1K5U4+5jqi1+Y0
YLVf02NMh10xsGT4tYo+XTzVTxgyh1KCz0XS2d4FteL87Q0ESysz8Z9c1O7+G0fb
vXn43T2rE3Qd5KoWZT0biJFsVDMMbirwc5e7Bkdx3rTph3r1zwf8N46QI+PuMji5
4KLywbFb3Itub8ogdRUQjBs8Skzukdgyw8rTt7WBn/QZhQhlEN8ZgvWkcmqI0yG3
iYfwl/V3DWSsDfhLbtSlZA+YM+tyUJa3WLeX4ISYr1ayv3M+GjfTkQxC3D2jdUyu
6gd8Y0BkQoNmyGDG6h81cXToLCzCm6jAjcC4eGFmVRn3ATaQNCjb80xP8SXtRbF2
59tGeWoblxvIhQJHPyCZQVplIDRhp5OXRYoGeLZWnsBuSYqVbQu+VoC/I3cFaZJ9
fEzlxMJDTukIKOefb2D2rof1RlhUv+88ORAZ5I9TZfqFnnaC+D/oHgaqF0afiVcI
/8txXDCNfj4ye/KiG/uCEnW5zq+i22G9aZDtmn3NtDu7JXs//dRSbz1J1SEZm0TU
FwftMgf4Noa28zy1QepKdnt5JlYhvcF+6J7xrR7fTnS7nD2H343pO2kD29UNqEPz
w9B4L3ksrlKDHGlBMEu2N+10Xhi3e8ZBXewYwyAtgT6tQXpi/fPh3wnx38Bvb5ND
UKSe550uf6Pr1VNymKc+M76OfLjNL40r35AXTUoZP4bNVoUQLsBgy1h1/n6hnqNp
RaRW0QRMEgNZi+Ro9i9KwZCRRBprg5U/C6DZSgCErELgiR35exefnBvURaSfEamb
z9L9VqGTpsQEezH6sAh2lx7C6qwQWrrDlaI+lyG/fVOu6v+j/gCBf5mtX6qNIq7g
ZaYALaKujZVvfdplNDlZn4Rz5exwmMHyiDh5afyqVD1O9kxOo/K2g7M5lGjdoS4h
MzALzHhJmush/WmZjawRa2c3Us9uzE8lPdPYVQt+XbDeTNATWBs36JPmHH1AA/Hw
3biM2kQrlQ6WQPVL43i1eV79U9sEO2tzFP+obgv8zROcne2iDeAh015/MjjOK+Qs
zgX408BHDBAx5CSDJkDrhVE5YYs1R0K/p33/6KbOXEp2l7xZudw0eeI/9ZusMwmX
TfcmfmXLuZaOL2y3sJmk6d8Nfgt9pSLy1NSs07ihbN2YFUweU4BWujBQf/WHnouF
e/efcbTWH2wikxE4iI/fBj046G8gul7AOs2embmWorjpZmOmMnEZCa9+QzPPcbsJ
C5pXbtYQ0aDbHLqGXUwSBX969K4pJ72L/L8DaILGrlD5ilyDEx9VOV79/q2Pd7lr
+Dibim8UXdHbfbcu/MUVXQ2/PFWToWyDjja9IjF9lveUjveVFSyb4Ejzeda0k/D/
G2Z5tP99lhbewOthWGFQCbUO+Kwb2buwc4a6hmFx2NfNbanKagOO5C029KiG7QmM
q2gKUs9MYxHnCL++sPTyVmEd/fKPlgm2ae3A9a0HfSu/Fqv5Yqy6cWmH02QskktC
CfyQHVKXuVlNCtNtCTO/5hE08x0E99fO0GmaFPXykFGIm910x6kbb9uD0nDseJh7
5rWxtHga1mMQrg1YTJsyhrKGZfoVJoQUJUdZepX7v2VYiG6h9KunRVP7AIp5YhY7
0Opz2Thjul7OfReGxy76jKPwRuQNLhzVyskADrc0hVjW26K0znsjVfY/WsOe9C1n
0Iaj1WTWUUM6mMjoA9Kf+eZsaqTqh4jcNKt8RApe27nF3ewKrSw8Ea9ERHsMapCz
ZoKpYKmS0iMlyv/rMDTwVxrQu2dvZJ380cBwzd0Y4f2A8Cwh1+TI8EnuyCqM3Epy
nz3tKxFcWy31PRX+MsgTxG7pIQYsC6YUHC55xE2FGqu1rsT0cHYGrt42WsPd3AsI
f+yVhcY2B6veD1zYYKxjBYqjpHGHWQHdh7w0lC65Owb7Ac9cRWEZ0R2tapkGF8qZ
P9lG2IbS+1eJbAouyDKYY91mT8nsKNRWw6gM/EwlBX5RtQu+XN3AWAXqo3YZVmSA
tWqAAhDiRkOFPv8F5UOA3PLBqSQ8jx4NYqv6J03RxoeTm7r86WabZmI/DsXTo63d
8OnW7Jq+UpFKWLnHRoM0OO058BKdu3LvdI0SiIF+W7Hyf8yXM5l1MgotGIqpWZhB
exOTMj3MOcWJCPnAFFTDuuZl1irfN0sKxXBA6jg68vRqXvRaGg5Aiytf+2emYlsl
Q0mRFmp25O6nPGPW1bDifJ2soJmGOLrpXt8k9M6eBKWyqgQUqfKiQ0X2MEufs+nr
SkHcyChbOUafQSpe2A6uIe2X5VUm3Vkyxms12/J4Av/77PnDCgR85GumiHSoJfdf
/BZuHIVXTJm1gRLVfBa4JyoMwH9MzwUDlD0IlWZNsgg61PYNKaJyS6HYis35nffU
O1K/hcLq/hjLjQ+/jyR5dFsK5zDKr39ldegFeiWD3lNZeoVnoc+NhCJV7bK1EhqE
7nd4sHgReOXz4yCd6tBpvctFJGmRcxirMsHqWOrtBWKneKdPwyyJDAGK+bMGqS/o
mzpRedqz1F8lonsR8AoXtuxFBNOZaFwM/xq25Qng9R8qSsirGSbETfrG0OzhVvv1
MRIj7NvVVSGnCWIUtrA3uuHjAUELsKARCJ/KkvwpjY2pzcNN+Jt/wNgh0Zi6AlGh
/ZVjBh8WNzrlIdAFy5JcihuVtqaluAaBkWjL/nvCqQcrGXKc6RTMLrGBXQCEBKq+
3S1PMrJBtLg1eEEmOF81MNxsCWRwuMcGfyMtQvUOK82Afj+JUkM2ALoXAdx1Dpo0
YSYTM3T81NjjRnZOYoJiKlpVxtvowEdRdaasYg8PtJjYF3N4TkZw0wYazinldVM6
Ol8MgrFKVZo+BxkbVSWgRMTCo4+3lZfb+l/5quBH7qcK+zVXY/xoXp4lX6SIt83a
qN7y4+Y/DB23qlAHwIYCvu7e0R7GSaBGMIO2vRdcWJdTpt+nv/HhKtCMcp3k+X38
nyHawdvTVdhoT1MQVPHv0FkaKPJvCMKftnUBcT0kUv9Uro7ikZf2gf4XmdUaewhC
G4vFNxadkTn9Mcx0Na8gKobkRT3aPH3jAtLjBgO+o1rphV3tvpvJQaI8OtIXtGV6
MPQs9BLcgXXB8GIs6yuZQ00VOO8tkgF1RPkRv47WU2pyuUVYVXTDDMvp92tA+1f7
JuAYW7GOZHbS5/SxThGUWdd+d9TjhqMidfPvteSfbhai1VpKT6zvq592DEe9TRaH
Sqo/f44HPk34HFSZxl7+4Z0hlPrltV+oavs7VmufbXucO/cccCe/zNm3sDCs8X+7
boEtcTQKfiQmi/VfNovz3WmpttSeOLIw6y99sQU9ukSDlLZ1UfucajBPtfoftok4
eBfG9u2J5yzfPAgbsxMZHooe1vFNiPMXBWnDYmxOm0QzfF5XbKtvPOWFrVCuGmxk
01dQS7JgPP+eOibfPAcnIjt8o9Azub1hd4M7gvghh2CeMaIm505zapIgnHXhDzsJ
FTm5CFcHZTYRSiy2fPCNP7pCjAe08JI+gcGm2U1rRCv+PzEcueCEm/61SIzxTJ6T
9ehmkmkLhxH2TdBsadORGzo7rP/1ysKK4W7QvfYXuAenQhHhnC6jS0W9PHsaU47Q
L2M6V6bNi4oRY4QzXQwn9TVFBZWrYtpzDmMcJofwFjPr6r9CuUzUqvZHTDwOJO6h
egY/vIlWAbptCyzXLl3qEDZ67WM4vVy/nlAhP7wqijADfkL1W5rQtSCXUMjvs89s
2aQm/IZGXqnZP3rc6pTP4e9jUKpTEQCQ6rVzYC0/ZSyVATGLvtexpL3UE+FpNOHV
2ep9sN/JjrUemqB0NIuPMydVovO992slTDfmh/BumvLAM4nLT+GtG/G/3hFuLOr0
usx3F5gLrao9Wg+3+/FN8h9ZgAbQiQ5b95g6Wc3QmzD3WSDY18yutVYiI62JtHBc
V/Qi6N/Q+5kZuh1eZl0KZS/EvzGMuuaeDFnyLZxJMFFB2EfF/NH5gY82M15iUbT7
WIDLDqUGPzalw1Hs61y3VUvkfTmvtb6GMMXx4uO/WiG+J/R4yV8J3hinu4YZxwip
UsHZLxgezYlHabHSpRN2T8mlkMoaML/amw5Aut3PhS4BFL+rMOdJniVqyZoN24kW
ytInJvNv2nSZnd5SCRz3jdcBg7ZbnzdTwGCqut/4q6hOrA5k9LgLviGfwfQRdJfy
rCKaAEXgyEF/Ly61ZedtR6xop1monuhB57KPkHJjSYKZC26IEauqFu90ixdQT+GB
sZaJV9tdrpckuuTl3M5TmGfL7GimMHoT7SdgqP3gxwqDQQ0upDAHDgQgG85eXs9k
Of79H1cnnFQ33Ou7SJVbDEY8pX43av9q5/l7LeGtaLBmMRKzF7zduj2HlifkNbYh
QmwAsFhmtiCs1lkoTnpdL1awGkp/NNhhNIlJkCVpV/idzajcP4gZ4rXmXRGsscKb
vGtCbhgzvVeQ/DLNvcU+Fm5V/L1Qm/jNPsz4GnHPiP1iDfR1ShkxBvrwmXPactqg
2vqOvhQqyxhO/RMQFfULvKQMW9bodwtNusmM5EeMLHYAlVjhxQGiJxPWfxUrhlhC
wBxy3mfTA6D8efjjTyj03CzDbFIZgE3AQjybYksFLUhfogMa/tpFmEJgcBMbGnhj
tsyG8PI2kCQI4NtkoK8ifI+M5XIGLNA+2NhrVELpTRzy0/tesytL558c74Magxnd
mNU+THiVX5d9WCtF0q13NGpm93sWmJhE7TlLlYW87V6+F8mphRpuSkrj4qq95ESd
vS+FE4jXUnsmgC6Nv4atWEw+yhZIWGwegvwv2/918cXNHHeD6Gl3X6jxdLUWnLDQ
rDsxLXbnldciIk4OhBYE6KvVDc0Qq0jrw7dx3YE68JAbqfLLdV41qYxc/U9g9xq8
b0tWIpMCHBghlj3pAlDSv/vpFDBvB8nkwvOd/nCWeSf3N0LLon0OtLlZ6av0/v+8
HgbyObctno8Gwq3qVWHfwYvdpro3L+PqRayEemf9/PWKzUb8R101cUbmOorWM915
RfNXPHkw0WB7/Jj73Cz7E+b9SM88ro3SxMfc8ks9X7prCnrlaxIug4m1y/oXdMCy
Y/5P75ECwyPiCTgxdEAMO+FKc7FbIDQaOU7zkVKqi7lmuxcFp03rqfLxSlaySa3N
1BM6PSCoIXDfzUIMNXOxFxg7fXTXBylvn6w6wGehNLD7NoFg1XgZ6R1qZNESmaIM
1/DgXtbFxFieh306KoWmrgBBzM/AKmJF6DkUXfATjfUra9nFXQ9QN5To0oZRuEfy
IFvks1d4T15BghB1SYpAcCtzPEKnNqDZQzE8P7Ma7magBonKeUYFAfNnAziaIMxu
m6NX5SqC3RcOXuK8gmoMw54TWNGtCPD/ovFlCxfOfsAsC/ZVQ4aCO0spBrwqs3fU
Z5lsyrjVUlkVjfJEKg9FjmrTvhZ7wds0SyvDjyBVpcHEt+FejDkNRPv7Je13DKAn
X7+4c52EOb3y/pGYmsncD2/PaONP7ukD4W+ZLbaSkEvUMQLCGxySPG+onynghma1
3WtxyZTtv2HqqqIbXhXbsVGiM9xPRbM7gEATDWv+3frZwKYN+LcwNsx/Pq6AuM1G
9zhFMBG9Qz6tSi4eI/f/hCjIeo1FMTII7ZmLxZ4sYLDw+LkQ7S6ExFisVAS5Xlui
JP98QjL7eRDaKlYGiLu1EqhwRLiIys03ee0f02u16x21gOX4gREcGXz5hAHyphXO
pOWgeJi7Aqm0vL02AKk66IIh6rDcyxsF07rQJBOFlV7Mt6x4YPro3FO5INeEB6KL
HwAOquVVU671lgnxbWCyS7ns/t+FQNjj2xvxn+30qXz9YvTAbjiIYMZFHayahzh7
EZHPXk9C+Rvz7vlHAiUd1b7IIw2KDCzohk94lQhnQiy6qEGj2RwB/Y5Y79Df7dZN
xxI7YQWsF0bSsrKbr7cj7L/Ribj8zD2iuQl74wHeyuHEOu0sPII+lj5mMuP69UFR
GkerjoyUGsMZSZmwCDvOFpk8vSmBLAXfLiQA2jwM4rJOcNUBoy6fOxjGcEn+6e8W
o4re7Fmq8WvU8h8Ib+Qq9AikIAyuRC2IimMPEZtCHgdjd5LHED0VVILx1QvnI13W
+4/HCCA3tLtFMdcqWqsAY6dyBOqU/lIjcvUoLIbgd+CPeTbUO9A4vUKgotfFTLJ6
zwgov8PlWoOVKO4HsPF6zrSTuNejDzpUWPlG51Sa8jv3XApprHk9Io3vzSTSsGMJ
FEMHi5HWi0HRrBHraP1IS8hAqxF/FsMYmMecSv3Vtp1bASGg52975VvENCpFmd20
w7YIrZ+AP88oKtS29l0if1H4hFMV6K/PTh+eL3EywBak3pyVlrsX2DTelEMYJsyl
vGexfdqU5rFg/n28AZ9csw9Qcg1FWegXSkwaYXIlqiWUE4Zu/IWhaFriudS+LKel
AwCtm3w1QF/gqfDHZzbu4AbMB7gecMRm/qU2lys8SA9y/iHNuKeKTKUqH8d/MdGF
dyDGmvBvRTSWh4FBIfj4RHV2ZevewW6kEr6YxTlDvEPyLI4gmvbVeiYDvncLswjS
ZOT16fE2YONjKEx8UcBQ7gC3GYZEsQZdNOpNdnXUYprlla/XO+ZgQBMJIhrcMGqv
oti3Fl7HRiqZAlZIWbIfEdBKpGvjvFdscbu9HKMozvsl7ZY3Vf2YjKgUCqwnAA6e
bWl6ZC3Q5JFufjSGiPM6M0aMFY0JcpBrkYqu2erCHK4imDhAB8ghLuSTMyNrsGmG
vCZWtYVdJqXCdPmuQeCLORkzrvbtC968dlpxAspxrSGDxFbJpeeL9o3+9j4Q6GGQ
sDca7nuBAo5p4gI0cQxBNhZeYYwDqWlaCMSR1Iz5nEv6SQtqiBcGj3g8HY4crgO2
6t6cCGbKzGLh5/7h51MBmCt+XVQRR1r3/hRKO2uR1+Bk5q9z7WxEET0zIqLuXb5j
htWrVxyULGaiNw7fnoQsmaluVec2+MgMnaJO1rTZg/0ZcqYyoXrUMmo4yZ8TFbcF
Gbr6ahomWzvjKGa+bLYd/uVCEaAgqzbkhkc1XweaK1LZ1H5HWBaCaSgSg4WHxMtO
Gk/ZTXIjnx9bv70U30Wn7Um/9kaNZ85cf0Nop8n9bODboAXZnHoxAVm+6CjVAkR2
4FBwh9T620MqkWdw0OXcmHR8uQMKK8K5simQfwRjcuE+VS9JzRjlNRLTReBpioLy
QVnsyeNY/SN6qQ2i4AINhafwakLOLDTPROSEkNmqXPGL802kAn/R4KDu8cRJ/sMJ
HSw/Ic1j+Wv/3nLZCQs/iw67G3xsmrNxPPyM6G68FxsWkWEvODY5zZ114Dv4Xpv/
H6mU7pwxqeI6jWELREnHBzIil2ImADell5pIh38P7V/c1Qonn+Fifn+3ShyHTdb3
++AnBIhlCMZRtTIMtZUgBYSP31Qxu7rEW7XZ33KwNyY/ZsyUyWso48YHB6Z/wqJu
TQ02URqYIuOB2Snrk8nI4FtktpaAeQrsLGgKjH8YoSKswMZX7HfMMiyKHxaWq/Km
53kvEyxeGT4Kp/CRzrUudiMqiK54l9VgPib8lfOrj7SiEwvdmNSmVY5U2aB2IKWa
896IVWw4QTUnHbbZY+521sRjTp8yKcaFaQ8ul03xaEm53LSOieLRGQUpk083yOgK
KvZGoyGiKx1bQ/SXAWu7WUdPh/Bp3bFEMG0lnjL9L/EONR8mbmddSnh/yR3Pbt6v
Ft0YgDAntfWhMHZ6iqDT8Mt22OkY5fEzVqx5woHFFnqtVmF8mDKckFcsAZKs1rHj
IrrCp+qJ0G7DRdWD1Pr3mTlrGMigpGBP3p5OdyZcu9G1Cz4Hj9CRUXBk7yfWYeel
znS+MU1Vo9kJ5doc0vE+TKP+8xQdzLYq87OH4H8TPIfeoV+3j2nBXbUPnUwh132n
4x3S7W8Nte1Sm9b+wputt5MVjBiainqyOdnGdzWo4Fvipsmug0uTwCdQp27pxlyM
rSvG/+dCesjnq84yuuFhQdONGNHfRDQJtv8mIXYMSBTaNbHwL0mK1OTUh72rcozB
kee3M2FKSfNvUuTBz6XCelNS+OqmwG4+pkp/40dj3YkNOcnEaEy36BMM/PD907qR
Tbf20PRdZKhxsEEYhThOsRYPQDWRYlytuscGqe5jsBiyKYVFsM5RTtQWE5ZOUBkq
JGgMUv/PAdAmBokECPQwAwDDBT3D1vDsC0mZOWVBPihDRrRKCGNHaw2ja3FjPH5T
09XwEHae7Y1cIiwYznD+WL2hQ+VvBZzsDQ7SYsHUzgghX7fmYFkBbXcRa0eUMkdk
gEG0aNoDup/EETex5vvh1OVOjW9fhwogME/JRMjZzDcoqZfKEPWHPAetqg/D1DGd
yQgx5FoE8C/WWgs/GxLj63qpmcEWReCUwPDkeqUrIZwT+cILLfaVfQCiMXKo728r
BxGzT2uUDvLWA8I9pwyOyJXFx8caiN+UIGufdIwJ1A+dYesS+5V49YkbJK0++Dyh
ibyNs1e9DVi2FPhdxyb7sXFbVnYD5ulEONDPHl87xZJhWl+fvH2hhFh15BM6be8X
+SPX2NC5dAaw/aopRDX9LLVJP0UaaWQupVfwX/BsJWAfu7Xw6kk0ECEK6rwbGShO
nWaWb5dazHF55kqhJpdOpNf8ls/pHplEblcKcc8GIZmu3tXRfB23ISIpgSl0RxhK
eT9IVsIrtu4QJER5XnwpfpEFf2fGQqs3uay7kw2USNI1fhl6LyrDKJZTQd5WpssZ
Dp3v8aOC7jSJyRvyDt0f4qcCt4g36OpEufsIm4VogLgV5HDeG+3c+4a2oKmVCxdT
VjQH2ZLIgGpdtWMSG2kL177JJlv+fS/xdQcyVWHSg+m4/pjc4sDyoqOKAqFhMIRL
5r63D6I0EeuAWRu++DFS4bY6SRqw1b2gRGtIDhvdAD175uMowOjaFRL4QZr24ZjN
S/fUMj9Rt2uZHhvP0a+3/GHR/3fZE4lWhGLaYcg0UM8k12gSH+U/7cNX2Imj8TxT
5+lG+J1TmXbj0xld55bzMzLq9fhjXuavXpj7yg1GuPj3AhfFJSp+pmzywoVJsCYo
VzY6DScKZkqLzKveHhC7UorNI+vykSUKwNAg6K8QNbTVLN9lTgC/jyC5pgvelH90
6+UvGUKrTbRFWI4lli5Qw42P23kANDwC1Ksv8hE65eNymaIYWLiZ3WFhGm4f2C/v
Py26C0vmWNsHrGENVHn+UkN6tbx2MR2PJSHpVIkdaOUIxtST6KNa/EtM5kXMp9jQ
/yS+tGMBvG7w4Ql2d0LElUw65eg7wv5xFO/yrCnEa3P8NclutPeMpJbqvVIpCFcN
tHTbv+2ycpJq48jMqgj+zNGjtFg3wDAtuuODwxLa7c8n/kmbzOut5xeIRgcA6yeE
+JDUpKRfiCkQvOhPE11MmYHO4JTR7LJVweTSKZ/AM9pD+GUGrqXTitrHgV0q+yVw
Av6nM9Lb0dtCv6r12No/ACiyA5v1kwkM18kGXotCUXx8hJtPIEb2Zyi1sHQ5XHqQ
oxELOZp4xzD4z8hRhKH5TETbRY7sY5V1oNqM4s2EO9GhItITBWUiEjQc5KtCXO5b
fz7nX5F3m9fT5HuaigL8QtslwGL4CSsYBEFY98Iozy4sXhu0nO38PlsvrRmL6/Mg
vYzEHmspjsL6DLzM90JtmvApf/8RmEmxPH0Wtx1afhZRkbvvxTRNIEqDKy/hagec
kwS4iijCGwDEtm1zZCR55MsezQ+arDMlEuWGbjJPEBjqfAmfaMAdBflz3Md4xcuw
A3TTxAXFAEBtPlGFItt1/HEHd0UANrjlx8RLQVIHS/pYWx0RTa68izpxseiUYRZx
lACNQGDkqmN2I5VspxJ4xMVeUXozEr3KNxtZI3dTZdcFO3NpVf1LeCRyqRdiKWO/
lfx/KSBpBYzLS0V/UU9znqMYyGLqUgI95+YWOBehhFLoEn4KAILDtc2Y9pTkXJ4t
D2rn7++l8MGtjCrL1k92exNrusJk94O6R8FZfI6JHSIMujus9PteUxrlNY57pM1Z
95rJ2hQym9DIvjBOyuL7eMUKnj+mnpZ1liELkKdA4eVOb/JJ06AnAPbj4iF46SsY
bD7JFI0XZkmxiSD9tcH4vLioncRuit7DwfA+cfbzl+Y/oyWuzBGmpST0h+jd7h4d
AnUPpxOeAbsODsD8TLFu3Cvqy/2msRKrTtf+/dbOwqG28YnBe6MlqcEnWdoKg9+o
ddWSLOEBdxtrk4TpqrASjLwGa/S03wfshelbP1oRmq6nPnF7qOBLcFUmmm/5cB/1
qJL2l6OTSI+2H82ZYVrSpFwGAsN8qahldJbL0R6CNWIzAal9dHQqsWr2AfMGhl5U
0iPxxOxkkB6ACAYatjt3la+ikHdnfOazhs8Wwud+nw4wtwTSop+Ega/bIwvdqnyb
nBA0EDcxIWhtRX9SJNsQ9UD9Md2SMLAKFUbChj0XPUQEwXim32hv62h+UoecrI2q
KIzfiLg/y4pXJBOLjVIEvy2cetkUBBLg3iKERkDsxxpWi7Q7H99WR5+veU6JIjow
HFNwBQAZFNOdNb/BAC8qLuJy8p3bVFS+oAZCc1M+CYAYI1lACPA2SsYUBlNpKNYw
dykIdKgETs5jhOezpSp+E5hS6sqcHlg0PARZYIrunQHsR2cDv13iqQQow0nLjO+e
a9h6uGx3aEsB46BD7GwVfRPaOWsNHh7E0WmWJ/fnQa22AEKMWrUv+ylaY7NlCuci
99e5fcDOLRdYpKGfc+WsTFjuI0huVyz98wmmqeEPEFbYj1R8SqMS6NFhs+jQzlcS
YZLKzl91q91s4YOFM8wfYHE/n8PckhSwsWJqhfWVkRYnrlrSeFFn0guN81jbOHMu
fVNqNNT7kH7fHH+W1aR+3I1min3WEaqLBJUBR1BMaM+6l4XRM8nfsio0Q+zal9YG
H3CCkA3k/zQvDmSM4M7OAWwxZTTTB0AKHqlauoOh9ELXkybTk6LrZKrYZRoW+ByT
BqgpDv/rWWGrnQZ/7upsggOyneMVvsf0XndEbdRAPkQxbEe+CVUuoqGR8BvYNM5W
7ypeIwwGhJfQ+AtcavZLFMMCtStPHIDvVgvB+ckM1GodamuDPBnpqNiBAgSiki0J
IJPr3QreIj5GwFhAqExHXahQ0jahpsFSkELeBwpVU8dCNp0G1bcgr7GHfVmVBvlV
3HsHmzUbPHnRieORNxRtqKUjRUatAf+pU70g9n75uKKtYnDIa8ZDVQjltO7tBo1G
zH+IziyacOdRl9hes6mwUoXp7yn1Akfy7ykja5u8lAYU7mzspJAidztWBTazHSZF
TeEbGRLPSkxmjDktcdUPcUYGYlC4eX1XVlqLsBY7Ac7OY3Z+Mb27EvsBBqRWQFIt
B/MvMViSRmGqsbrd3ySCioWDM12a2oKGmQH19PICWLVXd2keCyw1OGZ+b+j7C4bt
nEG93iClwDM3/Y3K5obf8E/wCk13tAEULwJWUYHi03wDDZsUCilUabBQ0ftaRoAt
vBtFG/AVTh0RtoXzmN1HS5D73qEcFSjY036JgaZm9NLmPochLzUMHnxSmDL6Vglw
2oK/IED35ZQZyGcqURHpK8nWos0eCgtW3neqbk8d6D1cFosAgZcnMstUAAfXTIAt
iKuFA+tzjcxM9egLw6Pn1P/DUs4TYunGz37JzoHRJkPt64fzVIUk83d7gYvBheFD
nNF+0XhKuo3DRe8pvzrKC3Ww7FE+ehf8TFQZFOMU/BcxvhTf3WKw7Iezd9JcmPZ6
XI77qwn86OVQJlO1S8NN5TVH8QDrTbgyFF7pCVL4peMuYXurdBgHtWU2K7YGOAac
/oLgdwdfNf4/AcNbESjjOxueVcVT8t2scZVlcCDUvSGcnDApiwCmOrx69zvB5iY2
ozR6NSJyzLhr6ayMfvWYB0G2Xo3AtiMQpQM1/Z0PxEPWP37GE2ryKtk7MyzfHZOp
JKhHUqdjOac33iHf3l8TJHCsqOt9dN+716IiGSRN40k5diyg7uDsCcuUSDsyCDJn
9/kYV8PEezRjErh5NfB8FwNlCgvY3yLukprP4pOHYb9Ij/O7TajD9Zz+9BXrpNCJ
L6dPwMYHQmBAhm9XwjFUVUvHY8D78v7hNLhSh0U2AZ4LZfd8kSyekKAfzDqlEPls
y97xz83VlwbrSRM2zHAnDnazGWxE7cJdoCitpHLZLB+uAxmzoVAxy0Jmmg3nKXyc
C35CXqMd4W3YbbBeGF7FZhQxuVcaTCajO6319/2jc1iyGNuHaQSnOGEaEZOP/FKI
7E4YT2O47zPMJF68UwKV4R4gkW3MnNhWE3O7uJe4xZrEGLekve6g5G3xAhl3rEUp
IJv7DDxEV66A0Xi3owXBlEnfULPpghM5N3/23vgMiaqXzZl8K/gBW//zZfXq1gXW
HY7IiSQd/07oWu6tae5Lz3VKn2+zeSnlNVWHAF5VwkU8OW2pWYkKB4r0CG3LzKiC
CMUnUTlLaU+2w8oblu8aDBJ407Ss4oEbxrEi0DbYl1SLW0yPOsU4XYsFY8aw2wMx
28U1OYvfWkq7nyC4l5NwNMTwsPXwX6SvoRCk/Fqn+I9WOlst+qJBFElLz9qqhdoA
rQ+pG4hKTSlbcXbHqSOgFMexc5guXX1fZmcxjWX3lfcoFU+8Qyy/lhphN+3mbilH
+rhtsXO0OJiAx2jmTUxl1+kW2zOWXVl5+OTLO/hn9BPlkSCGTTWZmVttBfGZdM9R
zobIfOJl4VjNttLMu5uNoATEGC5cisQkPAnYwz9pI6wLNmOjERVOFX4by/t0MV8H
DVhjU4NQIQup85/dK9uQz98+D4R8yCN8+JY/+X9virhwAfF7GhfvhU5yWmeFhYjo
D5cJr7qHB6LsHVXzrGfHZDXLeMRSwSUFoEK6ffka6DeosykU1ga3gk+KZn1ImRrY
OLvdgL1H3nSBz292NIh9aLs3h6TinCq/a28I38u9ZGPkOiF7ZBKG5l7lZIbRYSjv
fanmODxo8GRNULmzgzuz7H0h2fserttAFuAMasCHPqoggYVUWDjuyHeXkanFb6F9
81ec7F4tKMKgfhQvYcdA9OcG2mriTr4SadF9QU/JaazPqv4KVmrB1v42Mw6pclhN
0hEBJO2X7V/2jmwWdJZtexY5SrcjgZiLc+fawgRgkBGVgol/GBlboabeVKnPwpIQ
xpMJX07B0IFegvlVNFequqqRIqNlKJBDDZ4WLzzuo3c+Mk8JcPAHhkH9L2Bp9DQ5
sh5lae3idcNIGTyMsy86sVm4WzC6f0iHY+BHdHyqXw5SmlQbfbkOc0sBWfQvqLNs
PkYSoTu1lWekDa/PjNQnjh6zhloLcTHdmuq64x6bbyva2BuQZb2GqFtwYqlp2Aro
JzUH3fNIeYg0u9aPMPVtxjq2GQJ8u+HesVZCu2wVAAi3cPVc59tHFQOCbHEtmiKo
P654Lid31M6W4COz9wGOJPJXon+KN/iZssawI6qtQ3xzSE+riqQDAYdKueRkwMqX
8XRjnLljxud5jUMwdrz2PB03u5EqWOBS6qnZTFP8oIg5WopqZjMAnI1tuqU7ls9r
C2rl3DZ0EjEo45F9JCZ2Uoj76YP0NmErjdzHjEwsU9IyqwYzFUopB1K1G84sGpzK
kr8uiFqH8sLcreSz6eMFnAungGI9+1xEAiTLVtGCQuUAJaMCLDiHVuiS1iJqY5JI
hrjxEhnFgbZ5AatjdRxm2gsPhSjLffcOrJl68jhZpokVwP3G0bcCpuLQxaA2rOpK
E6RtCR6bwT2mzAEo2ZFTD6hmMVoNscTCohO0D5igCNwfHJG10DBAMxnJ5hb/V+d0
8Wx16hB4PEPGnSCrjXCdn6dra04CcnIqkVX4tjTtTXt0Kzz5bylA9N6MaldIkjDN
VjDEHdej3gmhNcAihWc1SVNfJlJz3aSkBGQS3hyBQUfYnKFt3WeA/yH/KkOx6Frj
9RwoYwopztro7Eb+c8GnVNILSHstn22o30GaPLHhdOmAzPYNxFjlHI/77dPx6peT
ugX5oJS64pIoB4E2fiK9F2o5gfNmdpIyyDCx9HqYyKzjNYiu+4tFk3h3N8B8TRO6
jk1L2IAfFV558WsLDxtFsb/QeCA/m/ufft0C0KsRFH/tbDoxyO+mNOpd+h95viPW
U9WdmxDxxFYb6MiexNc0T9ECOQuZRwAOn70OYd3ir8xirJCXBF5Zcza0516O29BJ
KHynMMVjhJvcoZpXm7tWmI/aBCOLGc8yWCxiLThwOPQpO6qcY5hvLsMnJaRzZnVi
WhVUWNhuxp0J+GkkRhCMrGEXpko3CQsd2Sr6KArwjpicX8VE3V7Z/gGcEx0uORf+
OKQExkcUZIJ8eQZJRvZuGlhThtrp1W7YJy1eZGVaVRsiwAy3U7zSPfmVNTc/EQ/i
Nt6kvDjyV2BaOZteLLnRW5Qf0h6H9/UQmWzk3By5PqLVZV1++fxKckSP6B8X1xAe
vsPEJ1tNLwFSJmH+odFoqzybDmhg/w9Vj48VhIH3YZ47mSaRVbY/6njgGLTIH9by
UxDL9kVhEqKsrbaB8MDJ2GJAbLoB/UaVHV9+9cIp2+lm/sE7EnGoqirvr2Hnbza5
8VsS9da9jLO1vfr7af1v78VCyVnXIE1uFTT9RSfe32/OWhUvfXi3xccWiR8MxiEi
KkCtUSGZFlBZBQZ9o/8HdYUCEn4hfpEjEbgiPy3jGS7wTIn4N1EnIPCoWl0Lloht
XHAk88bprfFl2xZl6g1xnYfjwqkpR/v70Yega/of5SB9YODk/VWv37Ew+j9Iv+Te
35rMvK9+j6R16p+xPLzXcmnAlyHz3pf/ST+I5MhEa8vP1EbnPu2Qn/3bVPMFyMuN
SBHsqaVf4TxjHTBtkLw52Y/FhZ4lvTFrY2I3J03g60UYfRIh2lLv6F7iACO41raI
Ck2CML+VgvdO9iEgYLGa29ArTQXmN0b7prawQEyXKYMIvfBUO5nQCqiNcUlLshS/
RdE572fq/ZJalH4lTA6xjrOF/nrFttPru+GPA8f15QPAJ3zdK8ELuebkqPh5EiDI
1lCW/wVEU6F9QfoHTf7NINO4oQxlxgiO1NzJINijKBBeqarNWNL+GaAiVnxP7Hr5
az2BVErj/tpF2ZqU2n/QswwjOVXZJiLbrMsRf4eEcVRl79Aaiyhh2ehrlUM9WZ3M
TOaL4VLlm67WJCQz6otuRzlFK7SXkNLiMZHjVugMUmdOYfE7a3oFHZZGdSmQwOC6
Ww2lRZHjje+cqgf6NvnuELcVZ5OZpqofsf9W1saJWxloe2nCnbxZyxxGwXEsGxRi
cVgtap25cJ41eIgzaIcsPJ7i2EzHKgLFXkYiBhfd2wGDdsAH03gmCpyBJTc1yNm5
JXu9NWPL0MeNN4kH1lqnWGboAXIcR9WzwSIlKBE74C/8PJ2HRHyaW72jb9o/9mHh
Jx8Yg9TZYc5CyyWSWBi6u5NZcSkO9W1kj5SWuGuqjya+QJmvEOOFWji+m0z56mx3
DFk1+OVSA97sOb05NIL+3QHQ+RhVfuU1GB3YSUk8xTPiBNPT65/sA2ZgO+xc1jFm
BG6erHx6OXRhl2Er+VK2nQw5w91a1ZI4qm2eAJHY5dWQP9pM9ettP/EhxPnDyCeF
XlEj6v0Xj/8+G3UyLN95vrfq+82kTHbixqZKGbDNl8muL19amdGTkWZxg3UvzYYf
6PRxWt5/jPGx1gg15tb2gX7uF5VD9t+GbCmGe9BuePfASHS7Gmwuk3FJPyss4c8j
dPKwTY1FHOD7S5t1Efqzwhxqj9hsXhyiaOqFFwo0KgvVXtnp86tf7cx7odQZrvl5
9hO0/ZfYMsSrNnIN4pgxw3wAEcvKsdZuBU74zhqCvV4mslfGDonDl6T/LanUEXb5
5rcJSPFxJmIvIcJ3NXDYEZndBUAwyqG7FnrpCD2Pqz7s0ZZqOkBBHlpdJlZAV+F1
UAXzbCwWHtPLbJrazc/c36MWkEYEQbTF05V3YOO3X3rn47hzSCT+GEpHmz9pn/Mx
9WiZH1/cJePvCzZvjRPNNTDicEauAwf7Okre46PBne5wJN2FjT9iYPcwnCym90nJ
IdAuPGiExZwBsZoMzqYdQuwNiKj71u2BeeW7FOBMvwgx5XrjJmSZM3esAa0W0l4m
ESEdrt8UAkcpXGEDTqiPPTR6aBnUNkH14O9mowYT2nm22EFC9DV/XXpRedW3dxaI
V6NktBI28VqcLaO2h+HsP5kcarRuAg7AxxsN46JIBq7K/AaV8I1r8RoK81UguM+y
yrvbtIxEg4c8YbEbF+kohdhki2crQC73SyvgOT0gwAChDIoo0m7pieceAPd0BQas
JXWIRX9FDBf2znDfP8otuElS/fjq87TaRls00P4FxSG1bGc9P8oi6VqNl+a7wbmY
2xqsD6BoubbnUwWd2x48A3CV03/UemcOEejlEZTJfaezWTKj0unThgweHEZ/XGYe
Xk6hgIa3O8Pkm4JXlghI0r5v5AOkVvvzVRxGwq8q/E4LbInmYJymkBycrrpdSvvC
ttnTiOcdSgwOWv82l6XJGCNBBoJQdtCH2z8RKpCK9exAffR4pmExNW/S6vm7oKsj
ZwFLMSiNSG15AlwCDxULcfXpoZQq515Ah72ldFfjh+x537Mz31gtfgH4Hr0e4UvS
glj8ml4eQl7cnomuydwkx6p93SbpUhm5aFMN3X8q2XbSH1amfD3LZVC/yEgWE3tv
/MzQ2ZkZJfphC3mPDi0CaaQHPs7g8hzLI6NWTBbmujSiVyBjEExErMmGm5NXQ87c
Lx/mfde29hITq3fMHgvUjsgbfEZ/Akh6W+gWExxrCBLadlqFSm3n2cWYlwaNu3RL
Kn/a7TD6Dy5JUbATheC58max7bNIqZbrCrRQL7CJloPX5xeI5egYV/gDgNkN+1O8
N5cZbP9O6KcW/Ch+UhrCVd95t5D+faXJnOOGzhmlGCv3f/1RVhsli5LDDJLr4uvZ
K/0ZwwVfDS+AIVnlbavMwrPCmV4iHpyAET/QUB8TdQjCg+hZh4VexZnEmGsFsGhr
mU/mBN7YmCAjrJvbquuDjRVd/PlwqYv9gm9vZaWCFMUmv1SKgtKxCgpk4YFqZzps
8z/mwMe2oC2JPtgfJ8n6nmM5RgO+DdQBdWNKwkhXLqz3rH5oncMmxZ7LtjqIetI9
Fp/YOSIVQcu/DtorgEokWDCstqf0rg6YMcLJ2C2NtUrZ2BnOIKD3THE6usKT0H7n
gvkt2n5GzsuSQkrIEwHPXoy2AmNEII5ixXW9kJFyR7gybQ7JszJsImve5XMQoo/o
5iZKZm087X/rcnTmujNCzUb9kmVK+3fyfwlLvvvAQCSY+eFJxepO7ioZNNTTswv2
xiaBpGq/d3aleYDEPWw8OY0sR+iN/MgP6Xxi2tbURQcyn0c+17goua3giBG2Uzwy
DyY3yPARoSxueT3STnImXbzPtdzIdMmCyKAdqwqM+O+qNUGniP9MPcX2nANSKa2s
tT04nDYnp4B+q5k+dxQqi5+9YRs+8uTI8e8WIGOYX3gV2gN3reSK2KWdLTynwWf+
Rrd0zE8ODiYhdNpjEon/bE6ybQFsirz+p/zQAi3RWT8b/HnJRqPkKzAaEgkvqTFs
78V31mg0FelNlN//aXh3lWrNyDpAy9Z7O0sTS61e9m3+XrMit01vqlBfqx7YM8qP
MiiXpQ610fItMcBirhITJDmlNUKaAMftcO+0aApHTZUILpeK/vh9Jlzo/qEC1fSy
/rs+jHxVulh9TnfRMA6l2BKOHWS8dFcvNwjf25e9L5rgCEGDnaigAEo4JQMOHStc
G5LNfNG0jYr92inmEuschtTwnXKcTTtu6Lnl+Blumhl3ZMbPYSq4mHLUObDHE/ut
daA91YB+5XRPrvuRDtEY0ZJu7uFG45IGBET2b/YImO6CyZynxtuVEqvjZTrLi0n6
+9cs6HTMFR7PZb77lPgnRS4q35j/in0I485mVpaGggj+Pixg02A4+b95F0YeoYfx
DkNbAWygKAcB0UZO7AxDnp3KCbmihVwJIgYozV1ptOtWNXsfXdZf8wRRrdYoNLJC
Pfk6NXFB2x/sARrdGgRsRZ6V8fHUflBHfdZu8mP9/wkIbbhSwseTH3vyuZG/Ddw7
YMJa62AjikJmbHo5LK1vOVcSVd84UYv/VFWAED1t+1lkwxbGxR0TBN4w/H0b/74+
lNyKpjU8iTDHDLB9O7/h8cRRW1i//DZ4p5CoW2jjJk1YiWm9K8xdHmkm6t/7tOQ0
+TIBoivezm+9TY4Wn7OiJpvlx+6akxZ26FZaTE1orNh043W2JkAw0Ci55D/xW3nV
2GGZKUHbhcjUPwVr6RCiu4HKjm1vmL113ZOec98tBZMe8bU0gLRb+xnAqKdhO3b7
OYG2a1S9IhLLd9OX4wJgaWAb916U7KajmzTGjGHN3EfZlm/NnJtFJpk0nXeduQpp
GkskrfOyPBo/r+6XuNbhCTNMszRJv3HsYBz4C0xsgjbe0XUCtjgjB98faDArvvW3
r0OORZ/sFS7a2oYALharAd970fCI7zjiYg8TlsiIxsxLZtShIYUseyE28RadJErh
m5ob+Ysq4FSFrywea1BPbxekih813bZ+9qOWb5pramMhIKeWa2JwPNO3NnroJFS7
poMLUt3xDKlsfGicKs63zIzto70QmpLkFIl4nE5jF877wPYeFMcO/wwNscEoF6TX
yVk220SwF405/+GqK0kKa1iRCOv1xo9FrCZ8tZ/L9F7YAOjpXxiRR1FNn9HpUu91
jxgD4G0Lxeh9xYrqQ+Z1akw0zho1id7NBvArovdIKS6ercLoxpHeR8jUSlTWWIV2
2v+oi0m3rVPukK0pqjiBEilrkwN2FxXdw04n7buK/oeLRquXaQRHc3PuVz6N1S3B
WjKpqyVZlDepYybO7fWx4jIM8PEMV1HbsiYx9PVDh4i6pbjRylehmelbgKxliR4t
rITPktytsOrmSveumlZOXAHJk+EJ6Ca/vedK0ql65CDc8KLQ/PPh6vmCOIdN8xVh
gtuyDyTFoiVsV3kw3vhXGAisY1cxjQpsvniJ2UNhu47cj6WPGH+4FW2ABq/VJ59y
A0pkVbEH462O2fOudnEToGApgjWKxu7mZx4LeIBPvtCTke/hPNm0kZHoHSUUqWLf
MrsPR/BJFjVbyhEWUZ3ph7Bi3I8NS48jWay59H9Te1jSlsomTm88QBvv45BUCg/5
na79+REU0QRspL5m/a0QN7KjsAhRPQJ4G2YY3vPG3W0/HMdAuCuN8hiLWLj4NlEA
N9pSA1EereqxrmbsnFa1vJZrUHAEEhMZjqBN5WUW5aUTTJsGCEWwUruiTFoCezid
Qi6mx9ZYQWZO8ldyGkXBSSqAWmkXtNUkOyB4+5m4EN2apii+PAU4LLLjZd25HdXT
wLNls7YV1JefUyZyM1g3MwtBe9azATjFUq0469gjqur4/9oXnIamM1xEUTF8iV/F
vLpsNKNfHuvMWAjnItWH+ujFZaGDC7y4shMvGw7Fv9++oFw5B60etJnoiRzwMiT9
bLTIH2eqd315V5JEbadDy8h6h+Wwwl27Nq1Pdl0UlQgCxFzCoULDlUaC0OWsSBRI
bgEOU1dZctT4r7mNZSlVz8roGPswrD2FXoMGttJw8krnIg2qGcMlw+tv4JKVM/9J
c9tMDCgPB5UkJ/zPJJfhXRn/I7AyjMhQxyHw0qz+FR849IqyTb1vfX4gKkOOIRSN
9lD4BygTpIA5NLAYycAifNUuc+eGJzz0/V9g007jVSC44iH5+g6jnJm2hKt2wXAd
ROFZi0xUYR1N1B75QRWTT4kTRYAh7vzv1xOmKjZsDIFsufK/44Xkcw/af5emUNEJ
objnTiJ/Uepgrz6qzHEN0QTH877wrAg0uLjKlmNBJwOoUN4E9NlDFrU3hz+esDC0
/6hPYSvkrzrOjyUwjpjz6osjeMuJeebJJSREjjR0d7XxRUk7WIDdupX6ocrMPAHU
/MoylDLCL1ljYolfLoxswrt39XonoYCs0ctc0VBldz0EUBRVG0o6/MkxZO2+IEVc
jq7gitlGG+qZ2IyR984SF+UsQ4i/351CQfqDU4UYVPhgHjqKoQMl2/b4TOxut/RZ
LybTwXN7kz5G3aKps3lhL4j59yiqLVQ0FesAbxOeV8+XW+9oSEADxsUgdBHQVDWB
23yGiTCvt8icgXzPdrB5aT6RwYp45/upvckfjH2j4rB7wKNOVWJXdZnf7lhVQf2P
Ziw18MOp4Yhz+xuwOQ/Y9w12PXhfF0q9Z8UGk6iBrMExPwnaqevnXa0DfwFtNGXK
xjoWxrMjgVP5eaMSX05nZz4FPbWGDCUQoWYmkzqMdHfHagdoPNW468mcfohU5xya
toGk9/0FQXzbK8iuIN2NdsByAmPTQ87DCy7WZcJ7vfZE0P8qzGFEfd4CAvGMearh
niqMX4qcwaa2MccL7nDty6NIwd9Ic7COp7q3Cf7BCpzgGc3EyZLX4Te4j/Lho6RH
+6jv8oD/7bN/aP7Uo5Dkp2h6p8qaZhcc6EQ4nsvkYbNcJ5+zMt2fBxpjiEDrBTEj
sRpyIL5XJTPFYw+EXFrdbsp62n/ImW3MU2XHdmZJszH6jYphP2YtbDQi0g+2vXK+
AQ0GuFMZQQPtPUFCFCLxIEECqFmRFlscFQcboX5dGHuD5oAnIAX+4k+f1D301Zry
uUax9JYqE62WpE14cOrHRRY5hLdTUHbZiD1x8h1PdtsT04RHn0BOTIlMzq0mujLe
vANgZLGvpMgqMRpkdyJnFVSoEDaBJa1JHo7obt2FIW5toWy0zIw2W+xBxZYphAX9
XF5THbqd97M/Q7/27dbv8L3rQqVjlQsPJNWy1v4E0lJ900o+33TIV72ik4zAdEKq
NIplGdJ6PZTkaNBdwwuhGegoHuWlif02+8Ap4U7WLMVh8lbA2X0ouAhA3ZZLCeAJ
0Q4YpBccbiu9rdsG0EzopRvZQDf1WBAGDzF/p9/gdVzd3ilSYGh/2tQMqdGIQaTq
eZ6usR+NijFurDfR8pmEym92H9ivMtemNFWBC6iqqyjG+8/4nBhY3ovXtOiYAhzn
KkrmtkLFT/1r8kSeRbXRA8gq/QZMoYRewYzrnzhUa6QRbFQ/PwJbYUFIjR4u3bmU
oDwdY9uPlNq7QlBls+9u9HBKQvw5IyNf8NTiBNNKmzirB42YlCHgSeCn4GEGC3zB
9VF26R/G2wjzc/h5nRcZYvHHRgrjWUWRImTWgaZrXUVPMPIoARgVRmOomiBYUgM/
yLfUIB/yMgNf2Q7lCHBEfjGZZs6nNWWGzz0w4Hx2+jgpo/70x6bQs70Klew4gnQ7
lTI000MIrpAcP6x4heUzXIMLsomP/RmFVnonQ5TWosuJ6jPc3P4GZXStAVtzAOb4
rCy9/0v9UwT7IM4Hg5siMtoAjkvyjDpLtPKSPY0QsESktavWFCSUhsuIE2ARiRat
6N/AANirtCG04/bp0o6Suu11BYnrTWRWXSf/VY+321uOBesGARQocdiJzAJwgm2n
W/dfbEAYB/QR5i5dG3cErZTP7RzNmH4GK0CYlDh0bo7fE+ZMsdqLAECTO3jP7Iyt
Gu+dZGDWSn+au/hv6OSS1kCKCUyP2MfbyunkVit8Wpkd0xIf857C6UobpmcUIvTW
0aoLxUkk2+420FwGlDfPMeygK4Zj0O3LQwPSGlSO0yU81Px6Un1yFIdCahnut4u4
jIlHGvqRQI4fqhPsGQ3k4pXLI6v2SvMg6pzwPdAvPRNhYVsJTIIptfmo9Gu6kZtl
hXCshJ+k2g0e0KTu4O/JUmxzXjIFsGHmPogt7Il8A31PwFj+J14m8d6lpyvVfRVy
L8JMsXGbewkh8n91kRcp/+ch6fbbdWes0SlJlXVQDUs3JPM2d3GHHAXkdBAcPVp0
b8qR9jIwDKRcv3kdXaqDYEM5DRtaLxURkv24bqC8ZurdQ5R75lmM3HLLxFQ9yLy1
4emd+m9Z2WnJ3jhJUgLPCGHWRE1vaPjCTqEhVrm4g+oipcqm0cpjd0RSF8ZBzN/g
GMXW7w7SIifLeBNlmwbhnHDmElPJC9BSzCw2TGCdRF7wbdweNkPk1lM75Vv4xLgW
66jQMZzV07b9y/a58wEETCFjTOXDybVri8uSifpJ6h+jNEy6qh0r4IzD+MW+zR2d
CYgcjkFLIsNg6tmLpW2Zz4OfuvAmEwwA03FF5fBqKwSGFiIEi0vTTeqixXabHApe
dQ3UpsdH8rAlIHr4w54oCcgkpXMSVsRamcL7vhBTkC082O+tBrTd4XgjKQWRzvet
vjCk/a9c92eyMpjuYN7MtApFxP9HeA5uTzFiIV4HJR2dEhMJ4SbR6B8IDFauwok0
RopYYiDV0bNn2LMW/ylGjqw1Ic4CIEF+gpSsm8iPFFBjzZHbXVaPwAcLNXA3vgCV
7Jd/6N3eHlaZHynLPqFDrrXSSX28jeZBXvncDPDf5qj3l29xAItAxKv0/oqO6ApY
r5wAuXneFIy+SQRFousSzJavjP+DU4Byg15Io33uvbm+SJsu1cfkMGnR3HsF9jrJ
BMNLSCXpVHB3+x6PX2lVXZrzDkxXHePgF13bqP6X/lJc2kVuqjRu7P2+vxoT096W
594++1aQwrp2lUBJbBbl1XLN/Loeb3OOiniXH7uKQ0ga3HbHpT8wlwnZmXkNFVlR
/m6WgAFRgh77jZqV1B6vCnzRHW5G4lai6GBJg4rFeJnf8Re0fCADKwD6Sfv0UY9f
pods70Oncp6862pu8WuFSkjJBip406LTidJrlieuKj3fHgwCGXwnQ7AWgG4G9/oA
cf0WhEZcOdFcvhcGpBBW8h94la0yISilNXDhzCv18Lx0BGxnaKsrkoZky543sM91
rb3kSOUVoKRJBkCoyYoISNFdcPfQsuwogPbJaCUZSRtS0aO+qqGNhp5MTlSExWeg
req00GOYnkks8lcdNfkHf8jdcJG7unNT3GuSzg0aVsKvSMsFW7q33GYk8gY+9bfj
I0IkG4mEEzXeyuCCGuOAn+lO0wBRk5RiJKDxE+askJwB20Yd85D4ZKbRFedtPjuB
c5Mm0DmsyAQT8gj+i2xWds7arHYDXs4MbfD5fzs+cEBXx+eE1Fk097JffCxYfuDr
aayp0yQXHmY3ylqrEWUkzo1xt1VjNEasCrGGqc4LPgOK879VP252wPhGmbGJrRFB
x3s7WcbzgHJZke24V0oOEpQTJK8j/r4F5yPx2KuCb4TN3nIybhgYg3YlPfahmp57
K6cBPYs22fRqukFBaeEE2ydWHz1Te/jWh7ZA6PTrayvUxUSEhn/DK7luKUUIIGET
2Y7QA8Pjok2MfHAJdWEc77hkAtAEI+9b8InYqLeH/zjoXGif4kIeYCpRsUfqELf2
wRiCuUnte4utl/xSAac8YKo0+9w3V+dmhhoQ54vgOw/i2Vmun21AHvRi5t0PM1p1
OveNNpMjs+knChi907J+FWKOyn/2zgCG9W4iu42JVLp7JZx3F+BdwiJ9BFVrUHbc
1wIGCSL8UZ2Xp0Cgj+3hPJIlKoMPX1JoHh2cEASbm7wIMx4/AUVIjVRliMcVDI0o
ycsYF7DFVvSqXzACXLo6y2+fgPQIhFmK41GOSmxLsIs7yoEgSuB1dAD+D51wT15B
PNPRKt+sdhTbW+IfwXDG2OdEtbpXo4ZDv1+Vd7PRKJ3pv5FXSheYZ6k1EtsLwCgK
jLW9HHNo+h3DZkCUHTo0O5N40GakVKZpTi943RnT5hpfBVG3W2ys9P2LLSx0Tk4E
dZNCv8BmNZLERXl8kgD3cdG9II1nION+ST9MpzGVwEgPubgeFAtEZGpKmD52TCaC
V4vIE97twW7/jryIBtPY4zUcVZTiqoPk1pbvqIVjyP/w3wVE9dHkA4WLNwicZ1gE
3lJAp//g+tE/zgjwxqvBz7VwsNdmh7HC8Fusnw7VvCzL5hNDHQm1kwS36dnFV4vL
LOALCVpnpRprwbpzAJRi5pm3ID7z3x6pbUNBtwPPopuJJWI9Co6WZzNS+cwoacf7
1i8/ybSUnufKq7pvyDtX05X/M6d9PF6lvYE41piZv1GerrVQQQEtlQ07RGb5Bfvx
gYSMihVcRXvkFqt81h91MZkOXYaUv3Yi+6kD7KToGpB/UTy7054t7/2OC2mxhQW2
dm/3HTz/gSfS7BFE6hgW5I48nTMJl1S8coY9KVnbMUd703qSRr15TQxS0ampNMEE
IdylL+JdJoQ1QKVjSsV2LKPOXJZaQf5/ECGAbHbZ6HSKOzMEYurWT+p6NOamue6V
7hIx1oQEDLdp3BWLmtUVvE0S5fV4YMuvdx/1JrwfUMisXx8EKPzD746QY0r7Orgs
eSdJn8dtS8BZ718Lo6loMJ3uDOSeLidk+g9jWdGiZY4Ty5eGNdz46qCN1xLX5l6Y
RyHpPQrJ8mQx9vtE4lymqsZn4l8pAmOe92p8YBYdX4vfIM+FOx01c+qhbpCD9bEk
+uh8N24eAxNIJMHRKkdzaRUj4MRoqwHeFJq5fn/AZQ8hzEa+beTwVUrnCfFhiw9F
gED03CE0lNgsg6D3KSMJKv7DpMUDKt6qOkHpFPZ7ztS/Y22TqxDiFqyUKdC2QBwL
nYTBhXSVH1ceH/C9JR/wqy3HynyZz3VD6ZIZh2UQXjDvUZTH+sP9BT5CEMpprG1k
nk3MMYrmvfJWmtbvtjjVcljYRYwwfCflKHtGY9tmdSrX0Gh1sZ+gfOMiUQlSShck
De8TYIIXn4haUwkqYvP1Up92TAUBGxqBc/ppA5C3jhlM96B4BT8tOpNhwvjznxT4
6e91uGNN9pfCAsg1qn69/LovrXIOR3U0QQf5ySOW3dSl+K4/tH9dVCi3leX4pVFP
fL0kVDlunmb0V5176EzOvd0qdp+NZdIN6oumYqMXU4BBh20e6U2eZgjUqRqNDn34
ZrQwS0tSHQ537Bm6G5DRQed5PhylnLdUyv/mLB6a9nGQNP/nqyLqqaGwFWS1brYY
fh/hXskiNxDD05Bl/bTsh5dYcP7l8ENnr+U5oSCpx6tv9NgcRbmSY/d1M/EjvjOd
NzfeVawPocKn3wOKxn0RufAoZGruG+uH4IPEA+CxkmcIVfBV60E9Jw24/BxFhSnC
Rx3UmsCIbDKV2Yk8idan6QonmjlPZwj0AovNu+0DKCMcrMH2wVYpeM0dO4gtkPBr
7LnvyD6jabsVi6wRCZczfS1ZgJXF95Spuay2Qx2564Y2WPJG8OeEBgNgh1qw7X5p
7chQSOOOl6I+1H/y5dyViLSuPpSOj4itSNN595bidPDI/6kq/ys6w/ICqI9NpO3j
t1R2Nxb6K3Vblg+FVGdSa7IbDqzzVC7VK/TjnCg1m0pymXNmjJHDQyNtyw/vjiiz
Lu13sVJ9TO7J7sTip2GLIlOSmOnWRRUT4L/CgjtEuH1vWxnm0GEvcBq6dUhRmcnv
qvZ2Jm3fpcvGnj9rC/RJpCJOVelzKga89IpefV0curZKo206EL9C3f/BYBMl75cm
HXA3qtfY1RmRyio7LqoTc2ReKqU/kr/tqULEI9F/y3eEBLa9sHKV/6o5JuEf/JCD
4f8RpRh12M25NXoN+IVZmmttFwNKV8YXtO8tt120olGMDmi+N2j9ZzpIA7gGGv3U
AXSPJGsTWsXb98DQT/+O8OBaqTUNtbpwszJ4isQMMTjgKJjSZTD0E/UcNT+0jc2y
e8koRSMpLE5mAcI1BTf6lhjc4z1b+ororQU80J/pQ1Zp8yQHazKyeGW95oYgztio
X/CuvHX4OT26mf1zojXw2pxABqLHKEA4tjoDWKbebfmWnBpNCfDegdTLqA0uTV+R
Z6NaQuEl2Q++C+2RZCC5L5CS7AUqIenGBluTGCWtA4tBKKZaAH7UV1e7IvxyBZDD
t+4Cyn7KIJAFv+EdAzmDG7ViorLPEccwtmnX3IwkxabneaJGnJ+GJhQyFmMQ87Q7
s1E10yjo1c7rWK4uAaezWPFZRi6Li6lLxfLkcoXUryGglYGp0Cyk6s20n+/k/hN2
NRnAFmOL2Poq46L2ys9tzFnq/R+kkgj00yKPdUEjNWT5SqZFqfDE4o6jh2d3MPvA
hk/2oGs8MMF4c8uCCPt3LD1pbvGZPiJuKC+fnpIJ/w/dHg6Tt1QjgGD7zTzEagXQ
M2aq2xhmtioY2RULB2xM/xNfPnJvsvM/OMeDOvrCkJCfnmuDcTdejZU6P0i43LkY
OWnpfKqNAkaaKD9a67H5ZIT5EkK8+skijxcfvv1wLpLQTG+lxIylsvV+XKfiYx7T
hOdW3VYFIRBmABI929jDotso940lZnS77kNGunBK2M+Xuy2kOwRxSaQ/XOOmaPFe
ec8pVaTwIeWzzzho/K5jTN2n768d0PMFmxoBxYuPGEB00KQUYTBobQ5MZiA6nszQ
mN5ZiUP2ie5meOIsgbNTnj5gZTwgv0IT3WA4W2HNAVnaOAn5asfhiKyFuIWX3god
3PTEC1QvU7dnzAHEQ9SYB5ho8O/BjIrmZT/2YaMxNTEXN/SmwGlVluqpHDVRkfoS
ACf+UJIYp7AbyGYBac5uCOeynkqXz+dLN/2fSPLCAeYFUU0PyKRPCxjFK8u1pmGz
b0JOFQpzDOaKajkAc6frnVfgeOZxDNsSTSi9ziyay7hHIKIv3c4LB6X6SdUtyj+a
ufSYqQKlMw8Eug6wqbc5+XAkhq49ln0OiXRB5lLKMqH38NsNLpPvbYXN4SF4uxLX
sdAfTW2ujIqZna7WeJ0eKLHUrk0UwSLzSKlSo590TYu/P5vuCUyOe5bo6zCAbpYo
R6F78U+iXGMI56jAtD7rE+gKh8P+SrSQbJUhT1kvdWEmK3ImL+hPsgu+WOjDd0fN
acBLqtLONQmOvX8PY4sFtWv6A9jzvLis2bTbKc3qfh6jlp6BEQbVBzp8lFdnjPLj
EmoALM5gRPTtT3DqaVfdYTPJpVa03JaYQx76GvpEiCFhUOXu/zYAsxa8b2Pd8WVX
OD/UsK+UzfCMNIrrxsxm+4HRh5B2Y5sBC4HnaX5T7ZNoDYYC8eiUgRB4rtZoYQUp
HlAwsmZySaV2zXhwKYBuFjhlY6y/BcjuZuoWfG71pp4RZF8p1GTggaouk89SCd7i
35S3VCGLATlsVzTxljkGsJnPe4FwYQJJ3gPvV/Lnjo53+hUiNqJFtVWsxjMwT2jy
ZDoNIaEIFAV9hfZoOYZx0ZvN1PwUdflhBoUs+Z9HUdK8YQ7VaqCCscKrhn2XrRrK
TLzstmRdR4aFzlV6M6xq/1ECVY6Xv89kMTjHdeSU5TOL9SklVgjWdkBlQb/Xt53/
JDfJaH/J6ROek7NM8BzKrYEeLY88e9jhyNWYjXA4UBcoluUQ8Y8wekf3XTHGPKfz
uw2A/DzpQFRnfW+vn1Vxb7vMg77NeRf0AHIqPUUovDv6oHIfexCjD9O993Ztu3lG
K0gMlBKaFnW+63b1XYq/ilR2rDsh+Lc74/AeBYecQNXljv/+Scd9UUuqBdPWI1Ag
cn2OLZZeDcjPBbad/VP+p5IlXs+Hoqiiw/3xKDExdzj86qNO6BSoGVR2POr5YVLd
HfZmn5Gtv+Ly5Lmoo3D55wn2FFVDUwX+UUKwRljqp+zqlumOKD7cm2KRwfzSeWUc
jf7OE9hODHHutK+5m0fw0Qz3PlHHzZA0Pa291Oz+igQn6lAdObIflRQxFk1DoTyF
5Xy33dbteJDH2uiTDcVuOpwvQl4OviNAKaXgoHOP2X0W1Idvk5kidTUzGfapBQRB
nbH1Pe4bpaw38t52LIPiA3xyLKBXlZsRBQ24F+ixnDpUI3YUkz8pc/xQp9+y81Dc
GUcZQAmOsjlynNRjdsaoLzu96BSlAFUNE3CCs/GlV+J+VBtt2s8H1NpNV/fa+TeC
9cc8+EbnAxPmMtCJdRQIxq7suO2a5mVOzdgi21EqFYCpObPihdy4O4Bx3B7vu8/D
r7lFOgfcMQBmMPnovM4sKWRitrl4iX7lNhecbJTqS6mcE/cgYgkH2gLCPpizGB+7
Puvp0UBKj4L9V161VLSJ6rTeMrjDyBpCnjoBDe2U3eDUJQCOczewIi1wSM0vhjfB
ukzsNtkBjdWzQSsImeE/A3+oG06YQHNK17m/98B8hVgVh8/RYuOaAl11NrQbALyH
1e1vvWZtIh0+y4VmKHsoqS9y7+kPfSIFGlYeYDlgHKdQp+PrabQiw2bwsOt+WTGI
OR8Q3yl+375WC2WL95F9df5U2wgjSvjJhyassFs1ZAbYFb+KiUAxxoWeb8QOoPXZ
LrLRqmkfmHqWiU2TrgnEzcpC9YWYk2NuI2CMD3zBhYiVtqQelzJdoZJBS63nzCgF
hzuPWuhgbh8F1eDQeZamOJRNRCEDGVCWCApodhiQyQIxwQdCmFkI+Cy3ghBtwQPs
FTTDcOOtphOwOsx8ze3xu54IStXoKPrgWVKqTHOK5j48FXX6u8I3BsGSg4oOY7gy
yZsdC+ZW42qgqo+LMRAH/2ZgE3avQ0jFJsjA8EdIxngPth/0+bZZbF7lL5tFqaND
bfAcrB/s6kgv56C6mmKt5ysf2rjbKxGhefGtw8KFqKizZ8oxZHp7uf+oNJ69FG4S
BmVfq2CstYc76o2A2G+bJIhc9nH+aFVqfQ9G+DTpzZ7+bWQ6iSImQprB3zSA5iIS
/wBVpTcVuE7zhM5TwIcf+bZ9hcV5L2nGQxYizAeFaWmkc7EMY7kdH9PT4ktvv8lB
o2Vj4C7tkcW5SMMD/YB5doJSfz6zINZKcqB9Gw6A/pAxo+JloR37VKMvFnwwfQ31
/wj3kPKbEZm3EfiwUbuIXjDv/zQli7bd+0jsSkfwXIfx/sJT+JaxjY7GqrQFHMLw
EOgqR2E6+uJBi8zFloqgq1tZWLXJgcGIk+cdouev2qD0K9kYKgWnXqMB6jsvFI5b
ohqqBdnNUM9KtoWuYdPA8ZIKq4qQeUQ87NXQmHsjfWaGzQNXHC87rnwRtPFcGzb/
yvE4JKjuNRvMuyZA/JOzdAUJrwOWhetMGHpi6FfwM9w1+kyICCocky92r2xSgb5j
tgzF+T3kwy6BwMFM02495jQYeq60dmkvFCPg/U5b8MY3bJZLypBsTU4SiueTHmAH
gqqad4n4XPpRLonuV1mVvlsOB4e0FuXK4sBzoqfPA/6/BUg30d04f8plGooARSRD
qJ0/oqU2HJejOZUZ0LUlYxEAtApSqUIHCw2p3axQOBXCDZZvbn3FPoRZnoAuPHXJ
hcfk/ogb3hWp3rX6hu6aJnWEHiecHC9vPnlJHdVlQVeJDR7T1E7IZHb98HP2DWtH
Ee8NQyt7vD7LIHxMbhKuxsV9Lzafk0OEn78ZRt5LkMPaxnGl31ALP21fxualfcAf
hPk6yyY8drgOEQ9RTpEbNVT3lLkKl0w5DLtb79XsjY+RSsXTvDdN1pFTtcCycU/g
HXj7jaQBL4p2w4vXeQReFMbmVRQgg0JVAMk9Fwukr3EBFyACGU2fStwGlhCqi2ki
rNeSbNCkzWpOodvoGW2+XQX3GST4iIfJ9vlQN9HXJFIsfzHkP8+APEoRGuBnySrM
hUY2ZFahZnQpcLpmp8OsDx7b3m3h0P9smJll7o5UemCe7kDUd4SqZ/nFLywCVxWH
wAMUYvg0hbND4xnHC76UDU1TqdSwcvkC1KaTEALt5FG93EFJhQP51mFXOC8/I+/j
DJub0KXr8cARTybtxhLHCREGHBNJn15SYjxQW/j2e16pcWr/WBvyYU31Ic7M5+Eq
aSYcQwAl6wm3mmSHNvR0apTghmhx2frcdb1R4B/JgoSqVQd2MslpjIKGxsY4zMXH
JaOsyqiFGsguRAR4dmSlB273UWnKHXe8gSJ2A+BbBy3RMt7utEGtxJylOM74obmY
NpwLiknlaqoK07PrUV0DAtszr3vs/PXOXas4TaUkHsUlnNXMchO36Ty0cF5LpR04
PmsrmAShuwYKGuZm/v1y78Uav1vxWbLnC6E6L2WCkVh6nGxPZyndSVbs6zpfpgLt
BXhtst6Fkmmx6iipWCl9XrkL3BfJizONvWjhMWInH265lRyisv5Ihjz+XR8ixoaG
o1wltEoCzOHcy/6A4r/NlBtzXxB6pf44EFjohxbuOSFGAtV8sgnYy/GW1tyI2JxA
O4L3SyRUgxcIcydFjnZLxZhfH4PjBDCMceE7sTKa/ZZ1XpE13A91aB+oghIEzNcx
38JEX5yuzOXmQuVb+nkHgMOq6DRJolWV0Ol0W52Dc8fA7WZY7xtQxrmhfVQ94p2I
3GrYQbYwYLPGH09n2xzEzMG5Z9dg8n9vVTDAIJk6M47lmUKCTLc0XeDv8vvx4hvh
oDMJkL8CONpBq84dKIWHxgkl1/QTNqhXD7l/p+ai9bkbBvfTFys00ox/gEenjOH2
gi71gQ9JZUQKenQqasE2KZRGgKWOer1sbXxd+7do5LmOY1Vw4eWjT7HcQVmNNxpb
fnTHjb8PXzwBAdCDQtaPZQVdWKcfjIBv16mFfZM1mctiFxgLZy74CMZTCY8x5dj5
pK9jQIAfA3fvOdQjPucJJUMEEC4wvOFeDL2LvSwNPMjWkBrS1Nerwv+H1+Rg3f4J
KQUhmzXW0BGJ7vFg1hKejEQsIr/Aqd8+sGHXWDBDWRnwI6Gbpco1SQ9uhzOR8Rvv
FrzLCIRuRFyUEhYllOCNRnbS7wYpVWHwqqD1iLpVhb7W78E0J4bF4GVFFaHHR5L1
LiPmvDo8IdYl/I9NHyzBzw/mM3O4DZPDeoqIo+vLaEO+vGenaCBmG087MYg74Zf+
RnbCOI+itfHfOfQVJ5mEcGXMt5X6eTIQQ9ByAsMlzZHkp1F+ryd+gEQhJa68RKMm
N2ttKBvHK3/6PxUzj7nmz2oc4KOXlV1m5fynD8n/qWnzE2DQt/YajTh7BRH+A/Fs
bBKp7mcwAuKLniRo9tcwZzr2M2WwuHWLsk9j5Gwhd+WINt7MbgzeWdm5Js0FWi3n
4NUvyYgAOuHK/dRTSS0CzshZJY5g+jpLOrIv2iRr6BVQz77geQnV7hL7fNcTaX9B
RTurAFZImGjZeXgCx4OeSt0QCx7vPVBewaXoK57TaTc5k0zyRlaOBVgGnZy07cDd
mTU/jqO2dreQgl/THFzYIgd5LdjoK2wTq+lYrSceIw15qS4zet5wyjcFeay3JCsr
nU6SzCVS+ftm8ZGvo1yMAbxASKQrnMlDI1xZypeyKkTbZUqU/Oc1jkvrr+bt0q+M
nOMr8atseniUct2AU08yaAtc0bZ7lwTfXGgMFdWTaaqAJqp0jcLrelHWZGiGAjgr
krxPCuly1vzC0RKlzla+kBkuCYkT0OhgP0PjWihpRhuOE+hJ1ZOJNjygwF0jA6QG
mFp/+loeB3nGXCTKgDuyw71p9kogOvxCHnx3SEeJvuQlMF5pF++xd4ssPFoPWEjT
bNbJAokMUs/TYhPjZs3Db3Jo5oEr+iL9IoZ8eJpyPS6P6c+mpDBXT81vKBTKH8hl
MwOHqmDdo0B7COIvU95elYEgvH00DlUKUmewB8V53Wu2nATvx2MlVCCnmQrR8bpQ
5KYV4p7wIcGHvkggA3V28k3H56tTPIBc19GPbHDq4FOBO6G6NwTGOTF2zGQkkOa9
p8k9CsjPemlCWFmv9szaV4qQ7RGAHE7oxJL0KJsGr4h1lYnZoZ8SoiVPO1Hin2U1
i0sZyM0ux87zhnCSDYGl+DM5BF6GGdNR7hMNLzcDFSHBJ4oCJ6KAl7b3vArvdT/W
vUEJ1xng9FaMe8elp1+qi43fIxazExDRhRdzA8TKv6BAEUIXFlfPMxq4WahyZUsC
GHyYdCmrE//gwCYhf77JO27C3H4jUS04fDVDI2aWoUb0L16EiCAX4VPkUoluWM0U
SRas1efsWnA200H6KL7/JRj0SLDwbrzf6FKFkAJWMP9dv/D/u+BqYA4/oNXyu4b7
Cr11seJnDS8/mEJfFyc1ppjn1weFBG4972wY0TuensC7jqvZFxBky0OFbyp6bX75
faCWB6gm3WGAARG0LK/x4m4aRp3AZ/xTHxIAQebTvVX/iTJMt8uqPtkF0yjVJde5
pM3iE0mR4KYi1juRhltWsB9i/yfIpA4eiCMmWjx7aYpwdPqg3JdkrHL/8BGgDMD1
G7aoqgiHd0ob5PFtLFRep3Dcl//EKEnGYYWPKvzDPlu22jWlj3AL12ebJazGUQkb
EQV+7purp6jbuDNXXQi+g7QVXfYCS7MbpKBrE6mbAG6oYG7G7XChasoGxrS2PpHe
/SXAStckGrk/JsU5qJEcuJ6/WN5POMLDfYGXLikgWiWsT7sZbyU2mzPobZi2C8JN
v6GXITw6HRhlZfy3cD+ZX9786hzCaqadiKZuRsqk4pP9WzahSFhU0KmAX5KvZdbP
r/+j9I23QQoFmExnx0LJd6vJuH70xLBvKctUkweC4ilv+FXG2eQ56JYByW1A2hMi
HbvT7Lo0hQcZkKeo1Ql/Ow6Cna6F51yy2Maay9f6YaqpYq+Tr4b9uS8xhY+O0Bh3
1esF2o5UuCRwBarEklAIs9xK8FRbtTNPkh4c2A1l2N2EtjmzoGO1FDMG2benKNcb
2dDztuBwlkwHdf/5wS21j9aJl8qeO7hNCcuRfHNNFYI=
`pragma protect end_protected
