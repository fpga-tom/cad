// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CKX+6DBtKeoKIsjRvNtEZe7pXJ3K6haZYSKzB1hpFZYg6TnGn/sEWaG1q7iEZKhA
P0Ue/m/b7zQNzdT9eOXpCkoS3sA5Zg6X8qtPzMLYV6GTPw53AFezYEWaB/frTi4Y
ulL1ZTJ4DG9mvFbNZsMVQGjg76uStDBD70iBSiWiLe4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 70016)
pJ4oxWXyLdfRlAmNE3G6xJzM527+QtyPf3c+eN8fK26wcalpKV2z11UsDpOrmSPT
EpJwAAARk/Uv4zEQ23/FDIm7BgyxPzfvHevKwF30aqbMwSdNTNrsj9eHrIoLMkab
DD1jBgvJIZx2MlEgTT7IqFL6cFwFXC35IcTxYyiShFod6LxHDiubkweCg4INASo1
l4FxxT4Ajha5YpVF2pB6W8MFrHKOjoidCcum4VvdDgRa18BA2/oameQ25TSCobRs
F7PKokG0ZgkaVHJq5IeSJ0+K5oWCM3Arb/757L0fz691NcAg+Nhvy1gHontECOfn
Dds8TSLoU3OHVhMHJZzmrIoVvZg7sG8ORi5PyecMrx3Jrf7MRtt0qKaycHda4ci0
t6P5zLjbVuNoj077r5jKbrFwSNbbN6/+/t4P72UGnwdDzXyLQZxd+x8vjgxWIaBE
fZ/sLM/f4gInSmojitlEfdukSy9cmqrIO6GKgz+yefO2X33LXpD40UrXfK2miHp2
BUz9J1EnCCrCd0cTt7EdBbWm97ClG4PWHtM5+MsFdaoOwlUbhViKwZnP93icrGxA
V3TBS02lLyoUZZTAaDf4M0Q02lCsRdggYqTk5Ph3baZSdzd/HQDi0xP4u/PjZVPE
5o1iq0ATLnbnGzdZWF6bZ+9IiW4nIBvW8dwUB6v6G0UhFgEl13CSjSHuLHd1Oe4R
MCMXdF9oqlpHeZr+GE53UmfLryZuW+Xa5J+VGC+/HC5q/vVXhH1gG9AQOy6z8YJl
reT9VyNUByGnbGKwZn+Oa/tD7jccxiTM9WfaOXI4bsQEZupu7qzEOfYDuKKiEz4E
rUVRRM+Zaa3pWW9MPqqlfjUNqVyDnPSdE3pTRJvrDtX69inekjU2TDuzWMxN1epk
LCsRYPl/kVCY9FBblp0EWAx4AfT8pt5YivopXcIWBOp0eSZ3jpc73AgHvjhTMqRH
7JZoqoSf+Gl8UAWg++i6IVgAhmBgzInqAE0GSWKcR1MzNX8eXG64qzUwYVOiFYIb
Bx2PbkdljUxUQ+OlIB+CDn6Eii7n3UMlKJ+kPcybGq9qwfD9EP4e75K1OHiIQIju
lxKG0zupToalESUxDWWvEtQoQOjMpC+/EmU/+05Q+/UWKgEQzqcTYg+pq0Qrk5sb
QGkzLPf8Uailk4l2TeNtiLshKFyXiCLWHp2ydWEs2a3hrhPTTiuvr6MitpbREqwg
8GaqoPfyMiUUZUzgvtic1X867GHPPxyarykcWG4cUCJWlB2vq6HXeBOh28/vE61C
rUiFY/DqDO43iR/d5Kki2lm6u7djY1fq7RqDE+cYZZPu2xv4l0k9W38zKrIskrRj
AkOSFuyzWB/CJnnC3yoF8SUSUHg6+vj4znRjrmm+Li6PBG196KBW33QUjCEet9eG
AznlezKdrPK1M4CCha74Z9pStbIkoUVAo5XCVTX6IDxjlg8erB515VXan/3u32HH
Y76yjPYI9YLbdiEGwAnIQoIN3xfvJFWitv83N3eprf8Weu9qjotO1Im4HHAIra8f
RzfhWbqb+vnXXEBv7h00LTq5IaORTZmveyu2kJ7SHUftSi6Q1YKt9YDT0XvVtRk7
2BOyXNiZ+lJv9k+P2MIBzCpKW0/kSml36WeiCL8cIGPkRNBXOW6g5d0ar4+dGfUn
Jpjw/+cuhq8caCKgbjyThhQftC2Ydu8uwT/rE8VS9/iY629BEYw6fcEOrDJBag9I
DLdy1JJ0ViiYGcR317bfmAN9JRZ6UR9HMJw/U3LTJ7ubkHP1n9blCQGqdi1TBfq4
4ap1CtgfxlTHndbYFtNwdzD8VtEBXpJMJG/D96yBFLlbNnzxYtxZF7eaSTMsQBvd
2GteTCsx5DqRxq3NlpE0M3dBe5vI0sK46Xnds+TxJcQ1sCzNblZPia4UeLzVKuwC
lEE7jwpYauWQvjp6xU2mfahcRw4cuQa1OhDW68p/WCBiyE1vQFUAbzFnMKJGmuu+
suoS931AZPOsYSOyJ9DJi164tbqqXbaiR4Er2TL7cOEcuTLY5FxbswlgSA8ICmjr
ZGaEpj75Bf+XdnJt4rIzY49Hooq60XstVD4jOticQXaGA13c/Bod5HjZLT34m+jm
AyFeWHNUQDqv2xwGB0ZAahZNGYGmKZk0LBKHqyPNPl03geSL2FJAlRgWslFHDlvs
x9DE5ffBNdAJ5qz2RHCLHhAxNFyCeBZKxrGgOoON/u7kQyUyYQ29lBOKBrnI74kB
H/b0FPHVYN0OzGInsFmfvfQGmeLjDSwnNvTruasMJu9gBIFDEB0Fwq6/Nm6a4z5Q
ScNshODRlAhl+LOyMJBwexdzbmxMN+cNTlHfhRY4BpSjojVq+K0SEXLuJ13fti98
mjIT5TaZEhsPHVdN57+gea4VxMgBMDBdwd5zg6PoQoJAzNEF7U0wy2laRIJVA7he
h97iMR/P+zy5Vfb7IPfoPyslklHazMnUTaGz9j4bTIPRtXnj2zuWSyP7+Mjf8IxZ
IJNYoKH+1H9GrFzB52DqzYmnOiHoCEc8U2v3IBtniX42vJPwabVHP+Y1HAIiwqqQ
EyAhtLRv3Ons8eVku92NvNvU9HQwow4kEmXY/iZPq+dM6FOiWx4ZT/rCpAnGTAUz
UDC6swhhR+FX9Li2eKn0ACBSgU9dxUJ2C4b7y31cWxTBEAl3S+gSaPJ/DrrbmAnK
o1NDyc71sQeoVHaYzopn1s/rgA0JMApaamMs+q2VslCP0c1sy8hFlAfgZixocC3a
QmhIz55nPfCKe70W3q6VzTP+7LXwdfG35hFFhfcMJqRnWB62Isw8kOz6ON0Fq1MA
wuvAgylDYv/c9NX9FrdNhNi6smFoEa8bnOSwWv7XqZyBz2x0c7PMHgSTqltx0i7Q
/1Sk5/gvH3xThIdlfhEWjPAYrrQY4WEEl9hf5hwPB3+nbT5H7UM25I9O0XVdDqsi
Xd8tWEL57mLeZKhQXK2zTDYAEb1Al0WoNsi/3mNlnelM48FW+U3jdnKeTdejFTTm
95gQcgiA8cbKkGzGiijEGHtCeJgssyRuzyLPbi0UxMOT4sx6FMZv1Cc4z9jRpT3c
qATf3UgvVzDEpQVTPGJeLGlBl/dr6jDGzZssBb764WTdb4eQCaBtCqbyJSAwvhOE
w8h0/MNKE2Qluk8Jgcp5ghIFH5IT7yC3OpHCGfZ4G5hW8iQ4/D3uSsrHRT+GWh/v
K8eEdY7K5OUv8oz44ZzxlDqyG4XFXhaf1biKd9sroKrOJknWQjO0LzKZdvU4XsL5
g8QT32B676RH1QZHtQjCaTL2I/8EGL7tRMlw2FMrzDw67FPeLxvT21pU290Rgtkf
vlS04VJKUulNX3I3Dcnx3ttHWQ4mgq9271umn2P2GMlNmmL6Bgfso1bd2sWFzVW1
aLx8KLFbKTGWXDEbX1caedOHhMNX0o5e5csjw6A4xorO0fQiVuagv7PoERAZPkG7
Y02kM0JriHL5pUH6K5ldpvJqwdtBPh6j0MCfM+MxD5seuAff+eHi/UzDbGlEngQb
4OtVMMezO8Efy5XfH4GWgZiLGUrsoa7sC5Tlyt9KJXxfI4AIfI+JSvTdQNW3v+73
JdKagdffzoseJqw5xRq68IQ9BLvgZ0MAN1KEtGfyE+2YdXw0GWzmzllunX/skLHu
6Dco4Kdamosxe+p/vGMu5LuDTWTQJWyi70WGdHkUY0cJ4gaOopJKPekBOJcZCjey
b3iKOx2PtiNQZMJV7CU0QdrUSLewkRgWzfHu1bhJede/QK1Q/bGmqoflSXWAl4iq
cmEPi8qKk0iPz3l38k+ov7ejd2YEa2ycuNUdi9WKJ0iPHnQZ+dZhUzyoFlmj53bW
rHzBABJu02I64aXDtfZA2Om5viET6+pqlxre6P2i/ALA+3R+1hVlw1Bnlh+bROyr
XsVFJxGS0tIbW+eqqPIefPD3i/MOXXYnWRm97zgmHs+SNL5ety0stzNUlKvIkGUb
PBekcr+FxP4XUXjKob2NuJQq7lP0bNzoHWOhvRrMzOe8fpFYa8vQD/LVKoamCrz/
PWhx64qoRVsyXUkvUWgXABws4IRM0l4HhhkUz35PVlDyvFuXcasaWu2ZLT/pXqw+
IyoZNjR5Rv0mFxCPRMbPFhueGtrcnKkydL/8uu/gq6l+0fAgzPiyc2eqFQ9hZLrs
3S/gxx8EuB7GeqHB/AzY+1WHo8vN2Ci2CXjxuFZYdwP2LIx9r7XyaFeZkKIvetOk
DBdNHtyVlxbFBj144kWWvzRQmyLOerSY63LQWlX7qX0KZTbjVATaeZ3jF0x0UVFP
r/sIdFsOdtuwySnrokHQg8xH0vD+cIA6jkvsnRS8+f5GErqoHvVJ8L6pRm1/kkmn
6BxZ7buglOzqgu2RD0fYbtREUZ4bhPF/is32xl4aR5VktMrg5oAlX7ztpxbc9xvs
2RPlT2PgiwAiXMSR015VvFsnFek3TYbpCkFWsiC+VbyfBGvDaOyv47peJYte0VDn
kB/BMNpCvKAqoCOTSkPYU8J2HmTkjQGhaMBBmq5nxXG1/g8ta86oG9MvdBA4a4jX
uSrfkSo2CSttLfU58n5bSx3zAgxcrLwH49Q+pn/tyoAspQ0lcKOcQ/P5YwYfJWqC
cxcs48Lw4HA0ZbN//YA5mu2PJkc7GXm2OGaPk6fcv5zCEtBqwX/RR8DxwNuS1zYW
HTPx/IY8vpLlQuXwJVNF/bPSzuk76mZ+Dp3MhYhG3xFsMH/+diCT6tpkEGHZkbSC
1aNx2MAGf7fVVpJg+ow/JprN3bnv9e28xNry1vcgtBn5crHwKfTUKpRAI5lsoctM
EvyWeEof2FyNsA0ZMbg9FgO+jMDNqhx6FCG0Sb4KDSfVW/5IS+NeItGHnrnhjcwg
ylQdRJiklyXARlK5u5rqbzU3q9qSybyjIc5/eM0KpzGIYuENwvXMqUSidR+Eoo9a
ehDcyVRgk/QToKx/7/kgq3w3ArAWIQVM7eXpVi9mPwPmHL/ia+DCluUOy2+8u8qI
Eg5TAQrToNLPp7vfGvd6lvP1IuIGpo5gzf18gp9gmR1G2zpH78fa0DOEZJBL1XX1
ngbVG3XBUCFv/ZYrbOU4gWpfF+Z3R8B+v0OjmlL8LYBggwmn6vrJAlRnXM17TPdE
cIaCp/rZEw6bHi9rHmGpD5mEE0QyeZMpZXunZb6ZNsbHlrzsuK/bn11XK4oIIK0W
z1DaxExxjtsOYWEbHWMbYGTc+RJem9W4BFMYNmvln2jTAZkUcjeYOQjKDkvL2inQ
GjW5vxyLRfBPLJ08kqHe9/h52IPVc/F4tqP/MOXCcYHq/ls4ICFOmQW8n0Obb90Q
IlYGSAbmavlPei7jp8bc2GAQMh2PHJl/n1mCyQR6Wfz4yI6rTE+zMz81mF/REMqk
IsdNPBujlteWbIJU3KksfGfofXttcT7uJV6N/IvmMTNYI/yxX9GK+YnWUivpb9Zi
yxidOEDkQaF9adeTMxA5jXNOTSM0qOyOnc8j89TGjT5tDIjLr3ywNYsrC7yGSkgQ
w6njNkFpzwiwB6Z7/iI1mFpZpN8vakysr6LD7Xk7VzifBkHT/281QKddN72HD8om
HpKxZhF6ogQJft4LgdetZYsir7IVmSrtrwOk1kBPUby9qkF3LXeCahC4S0BosRF0
hXNAddvVUvHnNC4npbarcSRaYydMkztIbgKLXqaAhIhJB3not8yJpclqYgq5MroG
N6++mcNC2MQMrHW5OZpItmeXTbyTOW4wrje2rq2XxuUrwR3CDPMmO+mb4sdw5Iwm
56b3tlaMNAyLR9Pn7NBya+syZpd02T5Ja5dF+HdrJyX+uxg/6CMbEyPWyaoOA5Wc
nJi3G6Jp40olWhE/XmRGEPfLwL9aWIZuxLksBvpMYhPk5kAz86gsnUTiPPa3zxxk
+It9nTIu2tKy+m0cEXd4sZLy7UeY3JS4eVWHVz6159NAS4cxb7w8LfseZwlafMCJ
UtKtMXStFBjvqVucwQ5S+MG6xfFj/5sFIGqiYLw9BhTmqCMjKWQ71OYQaqrKglxk
L3cKucCJyShZBJHy3xZVLRFTCnzTpvoDESVW/hveKUmvUkxYGgnoTVQQi9djtpx+
cOTW78kFzXon4cTlv4uoDAqSJtB+lj1xGVmIZ3h5mfntlN1TNQWr/KZxWs0bDH86
nLPJceAseqFqJTwZPBhCqlSPa+DC/YzsQQFcMsJf8JWYczGnoIIktpaQZ5X39PFj
qbe689LfLDgdnquxf4WUcAxW8fktOBgGAdZbg2NiR3eQXeg/2vX0wRlGtrQj3ppk
6Dh6xgOdTVwGYJ2cUe/Ag78xMMgod1gaRYkjE9JUSDLKECxsoStMbdzWoRvEObzq
lv0+husKD9qpUKvcI4Qgxk24MfmfD8AXWor3Bs37tGsW0oJXUkglrJX4WgwvoKXQ
MHIPWrjv7tNjDjt746grpScvB0Lgak9oIt18sCKpT2fa03+nA7679OwpQqosv9Ks
mqdddsr08Dq2CfNop2VrZ/rwrke1zgs1R3MtUBAMHadAkKLWMJ1zExi5M4lcnFXm
G/7wS1mdEaWjDK/CJ0RwLUCfDqJlZnvolhUb906LfPpeVum4M50n2KjQ18eL2TO0
+S+cx34ydEPTjR9TJsZiwTm9y0K2eggXU73d+o9On8BzTBpP0vns4QQgvyB/twn2
lR89M0tiRx6aMoUDiO2qjRIrTmhsiTYkIxqv3pJrSVA62wqVe1kbctrO2sDcBguB
zq1LAMOTyVMALMiBFTXCzco2NhG304s6SKAzq25HWd4zoO8N02XbenkJXwB+Yr3k
HMzCKtJbExVpGeipKXSSare6l5fKl5F+5ZoOwWng7T7IVwpfnNB7ofjqmDSqosR9
ngrRK2udruxrHdGJ+AihpEB6uPk9WfL7XzjQiyaJWw/bqtfN4qeicASLMsKkIGVr
RZRKgJnkPdsV4RLusj0k4ocq6gnsAWiWKqUJh/5V1qiVktDJtah7iFT60/mpxDgp
RPVU1apalUTNISSMidvk+XMliEtUj+5X7AiKUIpt0CCy3lCqNEe2eXCG6kOrfsL0
bv1ghwIrcnsMgpXYbA2P5IwYIDFLjETuAFsTX56l5TIAOv03w2gXl7sa8xQT1G+a
9i3Mo6ZbF+ojfUgkopTlsMiviecLqoJDT9fE/f97/cvDDxstUnOP86lr9u6wmYSE
zu11EzRFyQjC5MqnQvVtOS2irbAKoxJnBQZU/HlxxQYPJKiIb39g68pad5mxlsQ2
Ifmdnqawsjts59qyxQkalk3xkJAAWCx/EjZ1j8D8o2HSGH8pZ2ic47Lrxl5m7cZQ
lgixOKafWpmL45KIhP66BrxIJpztiXQWTLLMhPULxB46F9bqPYQ5vSQ6jwNlwg2p
rT56eJ3rUrsaV2jGmvPG2VJISTwtb60b2yQ2JNb/h1gEHEzWEIiRlK0HDaLZhebl
ukk/qq0SdV9Sn50tNB2IrvJF6hka4QeRqpxDz0Qi8+6NRaNfxC0HKTh+eR0S8QEy
wU1kZy86C1nPjy65LYq+k7CUs31/XKjboncPM2zWv6jYN5Veogzn9K7Y1x/4gxH1
K8PJA2VVFdRL1OHswiAAcvn4g351MuAAUk5O/M0iLMO4FS4LCit4LlZ7gq9otKjI
R6rndZuLYLdzBc3tEfSvcI5Ev9saR07ozXs5o6WG6mkdHztprwdVBqdopmIakS3G
iZABE73LuGt3tatuo9+n7RRsJN0Ua36+5GPyL15DlcTCVnjfUWvEZ092z7aUAORj
t0GRvRsSnsWo7P9wg4QdDHvi8t3sQ194RwWtUa9ZVI/Psj5srZXpeBUlNvPiiBVi
j47RJbJtS8rq7B4DEf/UQa4JDOls8/HbLf39UheafiwLpdoonpVtOAjehch3LdE/
sztToI6XGSZJgcQJuJ06xa9j0FanaNOHIeszmnyoIdQ/hhCNNNUIz8SzorYj5eBw
og/bZ3hXSc1fdzpPSqanlaAdzpR2uxomwQBb5aFq3Fq0lee7bCnYV9bj0Oerdrgh
IIIbhGruub1Jv4pXN8PrNw868bpxE39yVwSD1e+4oogZJ23AF0LyE+qdk/Epmm9a
qO0sZqTx3rPp6aW949nfYajx3d/IDoa2N//PeUtBgmgUIS5b/FR1nb3jWgXi0Bhi
PvF2pU5EPwGqNVWMAi+d0B76nYv+mekxMOs+1q+BDVEUM1SDuFlztp/ijzqRuDdZ
m0kwfnILBZoCDcr38A2HEiI3QggUHbRFrBw1xIrHb7608eZfNkWaT/wzsFm6iykb
ffEuafZnGyLOCDzGkEYIyvZ+3L/s/AWHNNia88Z2gV7r3JPsgCMyA8ciruwU2gwC
LE/eYEjb8revfLx+TcD/Mj+2F/H8KBD2DIfLUn5Zqd7Ey8IdtyurHTiOdvpRbJJv
2kA5a3/D12+QD2XCMKpAEwyb5ROwVCcFjFwpZdXh8Q6n6iWtDM/pf7H+Qvzq9nC1
1LalzjENj49A9UZ245eFyYKuFFSyN0cDZpHnlsQI/8nGsuifnNNVtPaN0WxI15OP
Rb0LLF0XKYbghlQsJs/ttIBWR09Z4XoG0dSwC1Rz8RfB9EXYEV+JQ/KJUFdqT8Aq
2FDPxXkRPCdFYiocmd92CjY9mnmFf/jZMCBKJuGLn4Lgt0EJ8wddHqCRMfDEiRLG
PURWCaz1zFj1AApIW+mOnZVO2Kgfgus3e3GpgjgnQ1vTnsWfaofk6qsOV+2k/hw4
vLl5uDspCuHpp2v8nrZutii4aoRh8dJKVFyBiiqxQnjqURNT9k8fTJAwYWWT1Aj8
5B4874TDkco1bjNye3QUDgRtclvKHc1nWSlHXYPNIrjVTUuC1mlm5WI94zsysWpE
jMTiEk1gC62afXG6z72RxPN0KGtXJmRrHRHjIVM3OT28CzDTfvM67TJ9hYh7/7En
NsZ5nRrjxjVbumUN1n/CF7SSf1ysiEUn/Z8+BlQqoFc3RT91kHR0x3d8xbloCcEV
0KJtMk8GmdMhHDQO49Rr8Z48VwCfPeMFYpFh376zJL/DcHLvuAVFqXSREyzLdkEK
WvFouyxC/7Lc8Uzfcc/AK5skuZiSi18TVA0tqZsFMWRzU5RLKA8f1wwaDCA5Keib
JNNRRnKIVALWtXwhdfwodFHy6mN+wwger+lNaKRPTFtoLAPntUD7bsYSSH5la6Pp
53ZjOZI7fdubUpts1A8KEDdHxBlRxpl0DGKZI/9ESsg5fTmm9Zag78Y8aUXNVDFy
n9j9E3NdwyDCRLxyNRyBuKdZiurpf0fQJ0NZXRIIeVyNIIIXaR1/FPu0Kmb3R9uK
Oi8KxBcupty2pPi8K8YstDbfihHuX47y8sFR57VnMAivBXlZCVc/+OqTbiK1bsA6
Fy7+wntQrgtKPvsH3tOF3I8k1QGJpQZ+512U8ZDpOowcuHNM0hyvV59+6lIFMlyw
zQWizEZpaEr6hcCqu9HsZLTh10WAqk3J3WmRlMFEuHEmi6iFOXREWQ2qrFL/2amy
bWNhZy7CebWqW/XEzQsfSi8ffRM1jZ2iwcblgoRpfqSRofT+MebRBCMvz520x8R1
EAnIgXCJWFCcKBykAcENqtcSV/fLXYwm3SrmB6dqKg/7b8xYQ1wDulzjZraUrFOM
+b0okOlXbuW0gV2HRTDr+MB9K+Zaavs+T7gyPW+PMes9PXnbrUeLQP6H8+zz8MNE
XOIp621T9jErXcGjZR0VmyWbk3rAY7+1cdW29i1+QuntmnbWHxlCZToOveT2Jl/A
NH2wGLuEq7jm8eci3slF+Bhh4S0T4KtrYmCPYOPxnnZ4GNltqQF5PyihLrgsv/mN
1f+XH49XkyCfoszJ9JwWGsjE9eAeSsPyVfIlWj1CfpZwmO1UaEfieuL0mHiwJMki
9X9cV+So+EdATiszD1VRRNxap9DlYvGRZS6yvJLAJqkwOySNUk8Grc0kaZpmKOWu
m0fgIbfrXBSFwQ7Vpku4/0UzHcbn32xATcHDdzkQlXIiToh3dgAOIoMhmBlNYQ/B
Y01sLbY0zn/IkRNZji/39c577158P2xTFATqFYGRtqEHSrSdAD0G1tV+oTYiu5FP
TIldGmCGLUYGwZKQuHkJh5T0IYLsFajDzQEbGULc645DrCMltTGBknw7NQvBZ0Gr
ZGVvgt4slEIIPzAtXIALoPFzKXYO1E1XfapZt1623dS5Q4YDahUkE9eY1KioSIKj
4d+NBXlV1l1nx3kr4elByhzp3S4WxmNai7h9pNiJAvWJBjI+4Sudbi/jfJTGn47D
+uVQ2HiUjLbSA6A6rrXD4AFJ0ERmBt/F4lfK7PZpPmOaWKj9jPADS0AijXnMyc2e
MD1EStMfWUC6gITSE/WIuwIUV4j+k7wCWPbt6MB5ALfC9T3PxIK+YMbv0lbBeAb1
NUQwtV1MP1wFodho2E54wKk1djBqM3Zkh0u7Dl0MxQN9QrBmpWFct0fKJUZp7RCh
Qrd6Zh0sgIC1e4ejhMWA6f2X1okuRx2Z0auLAQj49o5CW/LKiR2uoFIZqAiviA3w
TSpQ9ivukCi2cij/6RUNkr5ObeW+tKWPjqN39izkdXf4hoYdoWIZIQMswdEloyus
NpdatkwQ+8i2v3f6A7Mto7g9BcMl3yuF7698xxowBD3u4Mp/ctrMgo/2LyLYSDU5
N5Op94GYYphAcetz1VqNBvk7eryXKgdBOhGL2BZ1Byh6pKC+Daqq9PXbEKERHKJT
DRz+c6FfoHzlDYYiCkXvyhFdgQh4aC0Ionya/OR0k0VuMYgGDgbuh6kwNryM1bBv
KHBCuojiHiFKL2pBLIrUkxTmhkvJVp+G8y1BJAeDWGf0eb0csMXCEzUCS3i+K2T0
mHBJD9Q5WMucuJBZ1ju5Yjkem6CYZQ8NvsGa4/VvljvdDet9ZN4DrAi01xlruIjN
rDQG1VgSG/ReLxuKPoJQ1U7JW1tRcTzu1HvZ0gleWILo8h6NSaQabPE4+y8q1/U9
PhX3xUbgFyF4V6r4piplzmUl152oDDFAB87aDcA0BP6aSUhFujSCYkhj+qRMwqaH
ay6hEIRDRPceIbG7sGPxMsgj74WMMXWlX39najjMu1oI2JD70yRl57fwsfhZKG+M
YawO0QLAk4rimwlGjqpEZwn9BBgNSfsBlSCtNXypvxYRtV/ekwVKIqHVIJG6G7QM
FD4W4aFzO3lHMHh+h0yLFIjoS9/JnGOxOnrESB2FtIHHdjeyQxfbfLhtex6cU4jM
MoWoJ0C1e7CL1exvM0DtUPoCNaSl1W+Lxo495FatswqOLlGmxf1ewnBpQ2pFy7to
mvRjXm8cc9G50/L0Edg7XIqU44TfCy81uKv+p4U8S8Eeixms7SrujekYaHDVdhAz
eY6RHbJ9KGI4fOrmtpRzKBWSIeOlyfaE8KrrCY3Hit3csNJGbboTA750z+sM3gAn
2me+6HjT4L3oJqQhJQipDc6kB2VKhw7uexfbD89t+xyk6uOrVIsAoChfdIyvjJRR
E/gkApwNf2vGV3kE5d+scjVSECSwB+j12KdlNquUtq4gcKinPS0FGMTchhHP7kYF
6c73TAydBAuOFeCqXCgQonm2+Pc/OnLEMcDUPfpBqrR4MGyJDSmxROjCiVwGBTQM
PWf/heEU8NS+CKpbx2gY8ycQqz4dQJnjHTEh/u/1ni30tXAaG2cThLqAXUhppENA
p8vMqB2tjjabIcVKqb6BcaEZ+FRkREfHm1s5e958X2PgxgcXhcj9nyiTno8b6TbN
LBQBMNKnNUj4yGksl0xjm5JG6nZNB3fGZTI8UMC0Pw4npO54hviYl85lJ3vTCMZr
l6wQzllfG46c9Qh5CuEdqpVV6IHZFalbVSltJHxj0ij98BiaM8zm+oZYCCuPFEKf
ZGF5xitCSUySlawIOpT6f+6s+BIcf+D+JbLr5WI5AkDqUTqIkDbBk+foxaCEkAro
Gez+S499Peg/z0JVMVERCarcenZ4vEseQ7/pYH2reacTdJ/3zj+7QrUlA86Jxu5S
YYH6uNmRDUbBWedqCjHW1rrvF+jczl2oWYRvjjirubSW314Ivtv/2iGEW8QuDJT3
ibP4uWSQJXCwVNFzsLSc4n73nwHzjBAUOKTo2HQtwVIzsHmoVtATbJWxbeAjMT9l
Yp7SRPtXlY42Rn5ZsqFuHQE+7XRFn/uGC2w0R99ItS8XrdcBPYnQs9mNnc310w+A
Mv+bljQmINhXq2QJEqPbPtjohkc4BEqW1ztfRq8hV8P05P1MCXb+pqu3qS4jo5cX
b6yknDffAkHbAmXYpHeAIlr4o7A1mN7lFArJJ3kx24ZiMIH3OigaJ+QlIW0wGRHJ
mF05GGTztxtl1vWKqapdN15gG2yD1id9Gs4eoHBwWiHA/V2Z6NJioUlMENNO5v1U
7rzgwNMwr2i8W7YO48h2XJBeXMRuzkLaE2V+DLdFdW51UMyQfS2FvwkaPa2Ndt4R
4IZRQfLaUpcm6sSJA78UKJvPvBXcwSL43VHoSg7kiyvXPukbCwjtoECvEJzfRrXF
FuyG5JimsE1RYULPdKCJplOk+JRmWHItnIFHcW2yg/8dHwTIyhu97yF2r+78EaLZ
YV2xHq64crkiymGjO15VRIbmjO2JpHvvZ587MHwYOjRUew0rBd9b9crcyq8+1pC3
echYtBbAq3CfxNNgLKTFjOCqgdipqQqy/bjlRirKIN+23J3HkXX90Qup2sqnA1iM
qgJc4EdBV6S1ycIS8qbVp/CdNjJxJn1EFh2xgKKIWx66Qw0izfnckoPNRi31uevM
NqCJ1cJVRna+tZ7efwv474hn/Fho8wj4mYgy+KJo4rV+H+VWY6J+DxL6UyInhX4X
reHT03BS0xxENI+bLuxrUSkyedje4QYw3Gwkmhig81xKlzC2Ekx7/frCtAkWPPjL
I4CQT9YJMLg4SjWAe3CmRmSa/XOplXHtFV9rKtgFM6UGqo2SkOXaYXgHG+Bhrxr2
QhjYmw5j1+WRiOf1m8p3QHLdpNF2OKjkOkj8QIONYXnWAg5mdz6zcHnQIIQmIWx2
mgVyUguyvnKiU4Ur2t5golvmdOpT/IcG/2u4ZArCqB3C872Fhd5W7WAr8i5vQ5yJ
lJzGK187j2xQ4b04Ib1YcsH4g9cKCBrcN9M03drn2WnxNquyCBolvDnDJVJoR3nr
LAOT0kKMD+Y3RS2MApJ+PCKc7jXmPIsXgNoNg+iO4I0vc0L2vIDSF02D4rzqwSFt
v+ekudO8VGNXVP6IiqS0GTme3Cva49BuHybUFDXBtImjklYhliLJpaJcdHyNqcx6
Vo26Vjm6Wz6oREnLaexwpieer4U3nmA/4Dzem769IPCYfOtrliHklT2d1dmgmq5E
ePmxXfhg2StFZ5XKJC8r9fJD3e8e1kRGAy6TpqeYDziBdHSlgpZyipDiUHQcaKME
xfZjIzQyRTYsVY3vLxVBvLEkCl+CTnaD/MpKCIXLP11Ljru99prgExTwQNhWGpzH
6XIF4YdQm03efhoBOj6nTxpj3wLggip7HyNqiXJDLtboKJ1VekLFbozdglWoKvhj
NWEwwRJE+K6ppICzaBzkRzO92Qzw5xTj4gbupIp0v/RjaiYjNBnAiuDSFMJwqfW6
T6K29NaMrLWOuUT/8FnlbEMTr5D8CGrKJRGgg7TZY7z2KKIXeaLZx00o+gYtda3M
pNcIHJX3Wr02lp/qpYOlQKDzPu2Lg3jIJecwtAFWsEkTD1tFM1XIur5QOK8dX9KD
BIfu1YVo2qE5y0RoFpO7i3tRSTGhNj4U04++eKSCD4LlGyTa6gvJB1BRDqH1LRCL
RsGH6VPg384SWHH36cA+OAR94m1RE8fnJ5WyAX7r+y81JQLibeWqLxwZvBYdJS4/
u1fVc9YqjJQuCNNA01YicFTlVKQzj+NoRW2xGkaCndSn8KjwIN1q9yZCtGks+8Ap
MiEelCOubtj1O4SYAc945NpZTH6fi7JK+wNLlLTHjHBrUEokhA/mearhqe7yhPKP
A1gea59i0nZb6lxJrVsFFnO0DivYaKSz+THR9KoDPuDxgFAw7COhGyD6jNO9pBER
958QNmeM8OpMEM/48iiI8kVCpMwGnR+9LbShe9Hk2o4yUF7wfEaaA96yNDJDBR2f
oo+vAYUjxdmDotXClr010/2u/rU6IEWsw8VD0anLLuPC/+800Xiw9a2Slyw7y4cS
1AvxInNmH75Jqj5ZEto8ZfoHyrSevdSOuZefYYkiIVfGjZxOThF/Rt4Hw6I+8+Xh
VxqGPyS1VHZplMgwC//cBSHm0nW0Rz1QgGlAKrgJhcBg4aU3CH/dWtmb4STBnpTf
oai41XjA7f0JUTv0RaEyvnKR2U69E1HjMg/cFxB2GS5Momdjhl+LiC+tm+6ZKwSU
ClQt7r10iBcAmek4ARZJ+lUc9ZbCMd3Tcus+68ksLw7SVNk2AtdoqIh8BsiJV9KH
GYxDCUpSqc6Lk8xqNBaouScS1ZGrSHIEztdmgIr1HFehCDYV6AOzKQO9siSxOSM+
orsqR2+kdja+FCEBfijp0uDCm1kP/6N9RG/RGLkCHCdHty6IJKF5cfKMTnbjIXGL
QCsT/LbmAIF6PCokclbWGAIkWSdBZV7293XKtphQqQHYUV2sbauuQtUzRdmiSw/d
9MQxqdoO7PUF82VtO7o3Uv2EYYNmld5BvEC8LkHpjMtwG4TbtVJ8qiKn5rOFiyM6
dX3e0ROjaClgpWP/cZTYwnT8pkS70UWw2qpPxfI2CPVcgLNMME8aLrI3kTnAWHi8
53G7yvmiAx6Vp4cUyThZezqBHQxFt5lav1kJ6DaQU9tDdCdGPi3VfFTPwdiRcFnY
zzLVFlAobAqpwFSx68UymGg1pSZrg6z3vgKAr6eEO4O7p2M4XLzuKiy9iIDLSHMT
7xZ2whGEuTK7pEXvleX1b6VgXFUryUVSVcWfu/sRiYEcuy4bLaZS8OKeLlSk8Zdz
efcg/ktvVGJYGpCbqtpcBSZ8spmXMs5lEVtigNMQmtzi6XRMBXkucj9Nww/2yR8J
dUk2zpQlo3cqcy/A1SWwApuPExkRuVUGzQv6ptVJalvZpKwawdlervYLC36DdqOe
EIj5t6PqZr7qbbYeVufztHZxoEo4qTpt6JYGxxNC2gExQRebv3SXrKs8BtBy15HZ
f+Kmgp9gsX27VKP9kiTIDoOvHm59LUVvvRGHlZ95buma4BxKEpds34oZYUXXylN/
l5844oXPTrDHXVZ6yjuZWXQnQ3lFybl1GVjimCNK9LriXGbcIFFcZv8/qw8eqCOG
Fey281WrxqA/g1lTMnl1oql5neVufRzGCdmpP8lMDPTJe8xU8uCo4Nhxhdhz48/h
9MQl49U6SBuZBm/9Sb9SnLZU7UFL8g4jbQAFgmEMr4jlrDKydwxUn6tNSFZNOGAA
TZ5wmwU3lHaRoW1Mf1pUtxIYSTgP0bhdIJ+a2wLwjqW2Yvx6YHIdGv/xmq+RpjCD
b2wkt3/3x4H1Kv7mxLaiMpmYE+Uyha/xOX9s0t6P7B5tWrLsL8pLOWWsIy8dV6sT
BjRx4RC9QeJ43qYmgXlzPsqVA1le/3CvftPQStQVxLUe6buLj2WWIhRcwvDhSpcm
vDb7QpTI3dfTuD3A8mWlVVceMuXydsCBg97Ka1FI0+dkgft+wMxL1B6fP0ybnIbC
T3yXI+j4fUVAWF6JQpOaXso1FJm8q8hW0LS2k63b8nI3aQEFp6Ae4mS9tyKEU4Cr
OTyCsrmzmKLP9BG8ExCuhehcaETHojD2DLxqoKmpP1Qf7Ywjfh5Vom/+4WfZ2Ebi
QlbLDaPqJaXCazQcULB9swOG9T0IeNWnz9MEbAnbPk8bnx9Z8d4W7gW8Rimfvjtv
rpGhrZAFQZ0bCwZRcU0blgru7grZ2IJJS8D3rVs8DIFadybAmXRhsmnDMKxwtoWk
RjIoB19elHOJMgF9vFZTe+Va7NHWUK1FbIJ9ku0Fw174H/Y45q/t69yMbzYOH3bP
dGVFrcNPykAPT9/nHPkn7H52ciZFCZgisgeQheWQz//NQxicIKXdKBfzP8qGvRPC
axSWv50Pq6vVBzE68VnyImOrOP48xPGVtPYg98iXOHuNTruCjId7I6pb5DNapZom
ObDLJmXtD+EyOdkxQNayrOpCmZWWUA5q40SebgfbNE3FoceY3lEs8oUGeG0UbacH
OS5vGsO+5W5L0LL7MRAPs6Wc57M37dAXvGyXuCDm7Dr4qpI0K8plH+IDJRHqmkXL
J02fK13oMKi/S7oSZsMnhohrD0UkVmKtCFNyyx3J3T2m6lyRNg5860Hb5VUWd+vs
/f6I4KfdmUWwB3s4xuxWg6NRmRhGgZuambA4qSOgmeFGSDAIc25EK84l7aSDwQ6h
Ia6khIZ1IRg/A9wCc2x/wKKU3NblZ3ugbopV2e8TrvrX+XcllzRK1MFpXjpTrgCN
4EOSugq00nyH2OecDwqC5Zo4b/Zvh3cOB8THQW9GT6wVXNFBd3UGK4W84TWNyNl3
DK+jizTnqchFranDmVmayjnIvW9EQpocvhJhIb3vgFZ9BHyx0okDtxR5ZX+9diPP
zYbjuWn45lIiT3bdyh/ZXZ0STxb/BfuGYb0K6yEWcxqm18pjelkT8QDBWhATJ4Zd
olpdUKQCOZEIKqiLkzSNtqWu7iDMPWEhCOF9WCXAYsv4mqZxuUJhp1oF1tDUQv2U
p07opTlMpDZjCKFYybXmYeEM5XeMtyGPoBCk6vH2mzNkV4A3SJGV7CEn1yiwNvNU
rV/sqLNZhK+fJlaEZ7AF6xtzDpti55G2XPMfqdmou1teF63WeVAByZ6c0uy0Pl5w
q4N/YB7G4IO5ObtP/RlvS1Y14pfxJ4/U8C+l6597mgc97X3MhJFchgsr/JuMd4V4
Ugk7ol9W867AJ8Jp4GnFGFE0JW8wzxwmNXe1nq2MF3gucU7lgv0j+Bzw2bMlGIGK
th0GlE7fDvGi1tsdEv4tVyBgRtQob/DH/VRSrUSn/VZ57MbJgeBwXNgTzRBcKqEG
l5LFyyfaRyrs/loXADnjY/dd9tFOwz3Equ8iTUJQmlPSdxwcYX6j4m+ZLjFf4JJ8
DwruJ4PaZTw1OFqGdW4wo1MfaOmTG36yvDaYCzqnrzGULrf4EKRzKv1SvDvA2ri0
z1dKDDhUDMK9WN+b2QK/8xWBod6XaLGJ+ohElk2pET82FMWCWaRvjunvFeTTu4gf
bhd91csSa8elMwR45q8HFmfKhHc7wO4nnfa80QO06AsN7qb2IsPaUY5e5SqitKsT
oPCstXIQMnD05Krv2ekDG/rx8fRXgaCH36SgF+xFU9aXwOY+YA72bRcl5jGRl5Pn
cfBRPm5M5LfYmVy7M1hsTmVTA4HJRZKbzQUxI96+3l9XrMl5Tiokr76oTLUhIugc
OYmCKB1jD358etnC8dKQW37SkX3OsPI5Rn1JC1LdeRuXi1Lxmev9RuJz2+2Pk8Hb
Gi8qTw7g+CNxOvfla0utkf4jjooXmQjJF+kgdFNmUMBE4l+hlRdM5uUHcmCL1xs+
mlsnfZaE2DhbIyfv22TlYcDfl2NDpR7MgJAT52NEEgF7MItl2PSWB5LtMQLG3Avo
zHJErjcKdq/TLDtLGzQpzjo/MURad7FR0gZt8xFBtQptY5L5fVoqo6s40dNBOrDO
875r8dJhA86RVN98GRN8eMTHM276zbSzuV34bNA/UoZp4x0gQmeSlrEH1wB4c/gP
j5YFkuP80CpgnL2wYhyKQExvOHT1mIeOfYIJHUn4HY43XF3oB/ItYbWTtzyI/aRi
CZ6vTBGrWNE/bKLDqwO5FQUdqg6ih5lbZfxImAznHjzABcTEcVvvBvmreo00rONd
Ey/PbvQrN4Fbu69VxRPwVLT9Z/qnzOxYYCYtikgd7K4jUQFEJ9762/YfaTnmZWlA
Py2mOuu54B8lPMs4nHKxS+CzZrAl/6YE7XDYPYQi8Dta6qgOhrLg/L+ydkMGvsP3
SMmBTUvzzdGd/Cpz8BGeA99COiC3VAjkC76m6LchiQJTwONce8zBIZI4dKAfeYTU
N+wi3fyPst3BQF1/VJuvV816G3MkjDbxMHl50M8h/dRY0SqTrCsiBKim2PzS15/r
zpsXBWufmlWWI2di7qcP/8PgUPAjd4ZWClkby6qtzjkYO+f3+CBWO3TuSSYc/9E2
lY2wLHgn3ueTu8pXi4WtTtHqH5mhCMr1fr7Jjwq/oydINnG9xBexeDNqGOSw0vdy
I39M6mdWz8UTR1q0lIPFfkcd5oZPoGya0FdkOleZE17BkEj5+GYRyNrpiMc4CjDF
OYKOHxfA2uoqLRdrFFBkb5cjp6tJjEs0BikRoDjSgHn5wIUMFm6UlMM9p2kbCh2f
qxnAwxewvIr0Y6EWS4WM7gvdbm3cYKDP0zrsMeKCNhNp+bxvq8SVy49bm1mYyv5e
4+CfY//Okl09XYa12tX0KpZt1/LapRSooRzqShHzp7t4GLNS//crXCaI0ivCUGqZ
i5F8sXLSbqoEm3tHNUy6L+7H3hrexZHWrRnKsB0rXPQ1AKzNO0dbqWcNgkOBTWaK
Yb6G+yfWOUcksfg1xRF8J5OEv2y3rAIwnVxoLMMjGud+vs1QL4GzXW/pX1rauMFW
lR47GhJW5Cnh8/xkNFXnfBvygOmbqo3523XUmH7FUabjonFugchDfmNCdALna/zu
WSMMptX5zwt8zhlz3gTg06GzJoB+59DanmY4VLRRdS2ON/dX3DD0WIfvJYTMpjek
gaPC1yFr3jq6B5/ChY03BXjJ8eqk+RX46opLQwJbNrQ8s48RopeYLtonviTsv3YW
0C79KWJ4CtCDwVSJKIx+Rb3TIRcUCpjUsuBU0KB7C7eobBddGpyl2yPQi91UEwn3
uipK67KlqmsLH4d+8KRpP6IxHVcleLUMhEuTmod3iS+r4KMWj4blruB4X5a17pkY
bNjac3lJaLNOs7aV4YZHMvluW0oM+bmSM6rLthaN0h8rOsLlq7j/xA9VDqZoLLza
Hkhw0VziEN7PWSWZ1hdq8hVqzbL3EtuXklh8HP9O1f33Cf+WjeSohRo4dvjH3ECj
0QS/QTqod+yYbw31x84u3kORLb5IJeSP08GxxyTBum/TRp8T3CREUQo6KdqwVbsg
r3YhX3FaHFkKwE2cTh8uqHunjXdbIIp6B6Fupr++pTKcm5Ppp6q4PrEuC+bzIP+l
tMlMQ7CKnN0Vg0ERwNnK2fmyyC6sXfCThPj+vlHVa97MR9D910/g1oOJZkAurgqd
V7bjBm+IJLKa5q84F/trKKNLZTxKPc8p7g3Kalf5JLOC8j2flTn1d9v2iCFcR6Ye
pYD1E+qLzAjDGIozSgTIR6QUvMRouEu+R6tePikFaveD4l7B+fRHHN23ohINifv8
d7x94SLAIAXR0AVmDTX2ZxVJu0OYh1POgDbymDQXxW6sAvIC2deNUGXSvOqaPO3i
oa/237lF+Mv/I0IKi7P6KyPu4vkqv1PGm9KkLtQtaENch5R4XEv0KgA0JdZPiHlZ
4KVHFj2hv714wFdCbpJDJ4Cer08Zrpo9aKYx1NzHcO1dDffMB8nsmEQJC9WbnrG3
tV4FvlZbwPraKlkFmwZyDc3V5z4J2+o2xKh6L7yiqsyXus+VSgjZsYO7DVSegT7H
Q1yr7qAY8rHcRSswTOiCzb1Of5lf2VRa+gBd1I4TObWDlKbGjaWNYE6riPhQK6Bd
QJCMjv4EyIzck3v3B5Cs2CGZnYAkwoFxUDZ9MBwdM8G4OH0GpNbJeEeGamTdaSDs
ZALO4cM2SHq9RpcKAWfNml/0BvpObYnwTC6yS68GoRTSKLqrouuwUx7vz2RQGxb9
l9sPyWwIfm9/oBuWcySGrTOyFlJMffFnLMbd9utheQz2KNyUWW4zhTfaFW43ul0t
B/00muwEImrxRnNLSYhvN9ESoCFUu7I7EOK2zKO9sYUMfTJh0MHxiBjOkdJK9N6u
U+Ct+jD9wYlXn1lwK/HCunXEleHeTcYZdKQeVPUAKH4XspeCVQp2kL8z1eNJJLBJ
eCknjEIjNzA2o8jX2xDETHcCAlKAdNLQlxmrWYdhlLw3eYpcTvXnmYM8fEfNZ441
PfP5Wpd7QD8wYG+93NCltQkdG5OJ6h4JJfQBu+fvcvq6a81+LUQcKRQviabexu+z
ByzRn8RyTay+XypV4+7Qn3mC7kbW+tm3Wpw2tMHsia/K9Fr+yaXQwDB1Ubj6W0G+
xaJsa+Arhw5oWFhhufdi+FuJbxcvMCzbuZbD/5I76ppvbFXDODlfALRtXkN/NMVE
jMHBcuCm/mKjx4zKYxTuX/6wTr0R71XmY8r3eEYHGdldEHHW2+e3L0MBL2rVYh4l
yXiliDsTOEKH9AuwLaLPoh8P6wrcp33JwN98fY7hC8P2fOFUAnT8kdF5hkZ6KcG3
PPokqwv+glOBA7AxGmJctLwacPtKBP8/9KNqwkrU9m71JWlfnhp2FXPXIa5qfuUT
4b2HMyh+Sp7DAJ9uABp1QKHAqp5EkMA2GjcwQK1xbX9uRHfanaUfDeqqkAAYtsQA
a/yJGvtLC8e7FasWgV24hiXGuv61/Chtkmsnf9k+RBYBZIu8C9ri0coGVpf3XUPI
2sNBa0WXUIvmAM4cvO082ueytDUMiNBWJhf7WSsYZDy4X7VAHrhuwourWv8r4qFc
ufX4Q8P0ecRvHCLxGBbNksXe1kpcDjIet/bhu/oMIIDXMb0AdnaaLEg/pw9bmLqf
GnTgH55KOht5UTjOcI4eIOvUL/HjNtxZ9P8IX/3OYEww3zd/r6A3KQjp/mRn2ife
JTz/caFrIIRvSEgbx+TBZl9mDfxhuBs23r2GsEDkigvr0eqqffLlcYGP5VhRzi27
dOmemRYqce/3h7Q2k+YfuSTRUjvZDgCm+Psq2zTfTMbSmGSSEm9ipEPWIfS7XWBZ
RX3ExSxU970urJteSotsUMSYpnvwJcwopfcg/IB+UCDLfRW6NtAeF/avQs8d7cIG
o9eh3maP8Hsp6bExTLS+pHMnXTGZhXB4cENywo+tm2vqkWQN+mCw7m3mWZi2UjV3
6rkYqec+hWq9UXH5HA+i21/h1xH0TxqKo31TZJXNyuDvSgkL4TlAMPdCwbk4rH5w
dwnhdiz5Dz2AkM6tCGPe4Dql3+8rYg+HkOWPN8weB2/4Iei0HQSQ/QAkKSim6/Rm
rxoPBpYJwmXeBEH2vNCItJTzTHE8w0+DkLZzUZgnVYc30zbl1Of0xpuGdZr7apb5
unElE9hb/FzwySG64cHyour316ggQknfC5f1vNwgESQe+buscGLjI1HUS8fYzVL7
w9g7agpDe0A0jKU3OjiduUjTR9ar2iFN1CuiHuCZklZwIWrPnKqHWvREV+Ou3WgX
8tkEFD0zfBDGdJLnlYXEzCMlYMMRyORh4ZxzbhD5lMCQKLK6QUWnIuUiU3Xp4FFN
9KO+SuqPjmhwdf41jxOysxLVi4GBLVFp37R9gokkEpG6fGdE79B9TIZhOHtNZG/P
ddgAe8dqSVIC62Vg+avGQYsBH+u33q6c+ygB5tnVrVYGegIRJwhIsIkwSVJ1Vich
JE7UKQtkI0plKZKi23fhU8KC6GDk6SzT5XQfSxsTp3bbxLdmX+a7gO0gwNQV/F4v
S0fJEWlcG8OdoyKZod3WeMwt7jwyJ4kXlqXJibyWGHkomgz0A5YzxJO0WcNEzvWF
pRwtv1PiosjXPPfaDSsZm9nyLG621TNdyhWtT1M86aPODAX7t7KBnbJO3IyXJt/W
D9N9ODfooAW5Iv19l2f3f8XyvoBzR+hY41MC5AjEeJR34FqZduWBmbzA9XTmcfj4
MYoZ5JJjQZ+ZLPyQypo180uUrZ2aQvdcqHSnVcQai0kodSVuBhuGgMo91YhUWN+y
7yLxqb2XTnhN02QVYLOLikVgvqYnqdiUQhfY+nPrsAX8MSIN1TeSL0RxM/Mk4ZG9
u2KwkAIQEvZNw+qe+i+jw7SwKvASbe66Wx5HlmvL5NP+leu/6zPl4sB6vrk2FhqX
i5qAMfD5tQgE4lVo+zpssACt/kLncXf3rSgQ+TN3yQsRBynscQIUU/gF1KMAfnY3
ZhWLw4pLVacYEJ9MiMDdEuNRyJ11grVn1nD0ToU3flPquId8ZMEACsAWwSlXMFx3
VHXrV5UlLEFQsxvd5ehejHJdFz50Fh+d9IokVRaeId2a/FBI56BJdKcneStuYzam
LJAvWP0M/+oP4ehR+xU0QkJHD/ExpC3AA8+s7K1DkheBZoYZZyYWlGJx3Ygwdy+P
gVxIJaq4QNeU6IzEIaYhe788/Jw2u+0TPUmYbEvyNyrZIWtrPQZ3//QtNB3Vqgsf
rqhkLETpzaDginTnsczq58/CjSPe5zgT7lGXbAQwpLAdoonFEfNaHnW/OSl+EEpE
wxxYha3f9Mbnw8i+m1yaz/FDqQpTlo4YX1cDhPFLGpBZZC0gwTBn6gFjXrj6Yd3N
fzkfopWx7+VdCTpgzWN0k6GEZriXB08TPj/4Yb4m9RxkxskUipcxB9YznfCTqn7u
0P9scdHDqU7ay9TCXt5fUogIu7bK4Vt0oepmRcEPpACUXFoKtAw6Vdp+rpUcBw8X
uMEsZG5hZXnzx98SOj/hmfF+HZPMRv+J0t7vktJVH59EdADpWDuXJ1aFfDqF+Sk0
LcGGk/lD2sBpctsPNgfi8P0yiYVKMYkEocbE+1SadLi94/d8y7xobdBaKyT2Iohz
3QbK5XIhNO3ZK3jnlOJFwwqfr8cLGT34Lqfcm69vloYmHaKXJi/+0XOn0YXKUnOK
/fgJLn1RSOcFxnuhjTMANFYLY4R72N0jMSIFA0E95G+O5N2owLI0OrhlrbHfY6DN
DA1fG9MogGpR3a0DbfL7k2ptjR5GYiKd2ZsX+LO4Iwj/8urMkHtB0OGBIwokIjCy
lTSzNNZD/GAa5/R5dUpiN6imy+GW6601sOPhdzMzVhOBZH6Bv0tAh60USyDP7WYa
I07t1J/AFzy4a3olGp0Kw/95pZvfm7stkAV3D0+QpwFGEEEfVsz+Aue0eo4PgdBh
Tl3DEusUwhSjre9VdIJwdHkSyVk48Dl6UW/GEPKMKoGQSZOeEFj2Lak78vugl0W7
plhBczbxNAgvLbCuj8k86Szbz9zpKYUQmp8kPw1s45knisBWtXwot9kOUBfKZjgf
vwPfca0US8iKebM5h/fXXESZ3+Jb4UXacaqGxq7DXzoAVE9aayg81d+v7QaWWaQ1
dD4WX8wSEyfyXfFT3cM1uox3ZrRVB6gFEZTBGbEwXZtTeNeK+qAz2MFwGqlZUt1q
hG9Gg8Lty6Mlao8fN3iIF2hDL/5TGo9xxMLUcEE3Qor3OWo9ERzhLqCDU+/dqBdE
giBBWR27KjKgg/nPQZkfRK+WIlNrChmHNfkEuSWlnnrlCmWu7Q0V+LTnYElNj5RY
Al49nvp/RqbrpwQ8Qx4hee+cJnEyVE1uY1jptH4PWrtJbesv2GTQPlF/s8w0CUvl
nZAaKUixGsabzSf51YZXzoDE4ou/xmJXUgiqHD23djpRxS/m/0jtYyeNcTbGSXof
s2pNnCOQJtZyGU39jtWxUw4EqbOr16oscKdWaqKQNc/TnIdMbEBZLZ2EhLcJ9njm
Uud6v/7U3sy6b70KuuiCV71gQOVuwxuSaTckIHGo7CRMDkntX2+GmZEqJog9oQEx
sAhyNPjRYS32xcYzwyzNXujK8MxjbTpXNYKd3ATyu17qPcbkExDgCh8h46fXgBLE
Qg5h+jVEG2TlfEIoWmAR0D1hEgNzEX13Me9c+/l+e1lFcVjOVNW/nvTzKQPXS6tc
6aPOtD1NWBI8gH0wuSWfezP3epnL6kebBkmGzwRvh402iLpbA5oXmhCIAdpIBCpv
GUMm/NJdzyw8/osMtWuq7FP5LtJUMaEmHtlecUry8DCBDnrkZ4orvA337hX9TI4q
nGpsrAxlVbOL0zefeNkUV+jkL4kRsdNCUH2mKlCcTWt5wvxkM1wdV8b9VmR4I48M
B4aVJDy1m+BTFY6b4Ra0mvHRKHxjag+UF8YBYy1LIhZLyySdZ07cKbkFRh80aLks
J+e26953PdujxElIbzo09jpDrtYFHgM1O94XBBgB8sIjRYAcYu1BrUy9aUmf8X/i
Ps5ygTAcZVMJEWCcf7fFu3hKWxOEK6v2JmuJQujsbKRO1KYEizQJL73uMU2/UCKU
PeDK2jq9URGp0DGcevCFA+OhVEuRnLBDOCrsNXwgym5U618BFvFAYgcyxLR12EId
MJ+SLPHEGqiQSZzDbZ4P7FB5X2cOeZ/KHYdqmP3nmQl37VtGcLrVz8gYjSPW9Ad4
FZJzPrrcJaW/4uQ5yz16MSffK9/IY/gcR8s6O+KUtTJZGoij1TKErUXshVIEyhtY
g6fjsz0Ph83mrwdnrlM96owEgRtWYDOX2L64FHXyZ74WbRkDZ4aOGGgj39Yrq+jc
ObK5UZjQGrHDyHSyb49LPPa643e8VCHVTuw8pNBLNqLsmu1DruEtpqFPd/TDVZNd
hYLCnUWf+3r6KPzVRH6wOM5//vl+gmbRIAOTq3GN5Azv1Q1lifdukgzGooz3UdxQ
VLhVjcvyu6QdgTedokhE/MuhxES3DE+v6C1RhFMcj3nyeu0jMVL30LtaobBsoBEW
CGlBR91XuZw0aDiQ4gVzHGuJSGIN31ax+oIQYby5o7Vpzd5vq/2RLHZZgXhBxDep
Gtdr5tp6OR4cToT/pdoDVUP8Mr0Ut8n1w9sHbMx5jDIwbJi9PZmndNUND9dwUCU+
eeOpNiy+BM80kAIecalMITKhQXY4GsLK3OiuC80h87IOSWBfsGQ1yjTscSP468D/
Om2R0/6x79xkDb+/D49j9VTWZUA8tgGzgEwcqKccf2uYgJNs1XW9d8sBpwlzgMqn
S502ifzJCD1hj2INwD/nyWFnh5VcarYvJ2uDbM636RI9o9hkAihFhiJg9cXu7glF
3irVtnFyUXz16I57K+OQoVqqo9qfOieIuSicv2u33N58Gf3+eWjf6l7qFan07C0O
nXznoON+EcDV+YbQYOZclq+IrK4qgYCv/3Kr/JS8XQfqjOZL5NatP1RTCXC737bD
BiBLsOBPcbvxzL+PnUbclUHjrflPjwrAMPaJZA7247kt6kCM/8432usTNWyFv01F
9EmMnF4/dnA7NSF544nD4nNbNGTPrkthmqoM8M03lgdI99AlRE1lvsEYoF8nFMuj
fIZhA8b9ZBAa71TITH1FlprvknJ+t43CevDKgWH6bBBs7XdFCoQQTs4/bP8/X9CW
kUsw6Ir1CuLbNmTOYt4zWB7IocacJMGoFo32/+ODToxzB7WSo0g+ptxEQmBWgrGR
/59juKgtdmtEBHwEAZqjQZtRA0in2ZIJvcYP04o0Q4y7gNDLj+IeIoShumvrzXro
08sfn6EaqkV8mJflg9yAhw3tvJPBHgM0FkuhkC6UOKC+2cgr42cg2aMxF+oDy8T+
ZdDpYknLcwIC+YxMnKdrSxLRsXStnqU7MPmirgUvWQ3ts06oA8TcuGPKSMhfEXF2
XZimrUhfeC/epNn965NMA4mrBEOsoqYUTKMTOUv5YxYK5mi2w6qHh4Ynf0GqWsFC
czBJSyZJHNtbSxlEG43jhm8Tgw08xS2wJ4OVPz63VNm4SFAXREJqUTded8XIRN4X
v75OEydG3+wYc30LIxczCNMCjAHjU8b0PLpQ/BV0W+EojX7jS5mA06t9eNhrtI69
iY6yLKRdVRZF5GvF5i86yg5Wucb+h3BEqJsRX3jqMYMZXFH4RKIjsJoVskexGlId
VcThzuQM/f6l3SoFy+sY/Z7HxyftNSM84cFsqt1wC16pghPrjCMg+PJhdDxXXd0m
dpxBiXlYuuvFssu63cCNJnC6yQB12ineKZ8YMqwZx9CcnS20VzhBecASYsNSMC70
GhUUNi2pUlUXDZudbQtqf9fwjL3WkRNIfKsWJIG7xvr760aASA/6Yja0NzDntrd8
GoKN3J8CZfSCiAUVEZsILc5E1KOT7hG51y72fisaHpdIa/DMhqS8/elbPR95V73Q
qVSWXZ5cMg9+QRf4soLigC0c0YHvw9Oypg6aUy5YrAWsgsaI5EIJmpWBOpeYD88y
4DI1vf7lzId9cCw/yAFQRHGPRMUtCCqu8xC+OcCf7PFaHDtOBkrkHveI6SNzBz2B
Qrt1GiLqdNobzfIKmJK12wMoytyD1ZROWzvRQ5mOjEJXCig5VaSqSyAsPo2h5plJ
QVOl7rB6C2R2ISb0YikZUZOQOaO1fLAiD0fGHldupR+qhWoYemIAIQ/n0FM5WndC
fTnSMScSyviSRihYzfOLG8/2pO/nbuwmUUsVpWhw5C9P6B8HPGKdr1YuhlkdyE/y
nR8ey9e4hWk0rYAxYgs3wh8SNF+HAOjlNyqKPPZeWe49Oa4u+td3NNHnReslYxDc
ZMIxm7PAZyg129JdpV7ovIusVEk5rqJL4oWjoWb/OzObdBO+E1MWYWnIxFCN0j0w
t8XVAZdOLIRu3EMYggPdNfZ4EZzaZ0vD2hhzKl1yOJCuWXbtc/Zk4PkqITdCAEm6
xTE8uRHdYGkGKMqZCwBKYrE8MiNnMcCGgXmaVvdBhxrW4qsoboF7Nml3jClxdqGe
juG01ms8x97sw3+K5k/mjIcvg3CB20vhOHp9iB7eUwqBd+2WVsKMWpSyXAU5CKtm
ox4UpCGX+KJHLoPgCuXjinX0PKhbLoAtencaFp1EHuhnzHFSFuyeh76t0Ynyo7H7
s4oZBnK+iaZyamPzALDOtop5mrgPkchLrDlWekFRJljQc4ZYUPdvrOqoSn9f1cuR
JGT7xeJM4R5/vzJwak23VM0szc6De0ZkbVGbqM/79yNH6vQOTXkZInzt83jKgYID
AV19iqsvNCT3+uDLBXoE8R4brZuMPxHrbxDGV1MlkkkzixUYy5xtg4Yyp+bCMJr1
9oWj8EkTNg6Qr1Ibc3u1BmpE9W5XeNSQF/0aj5Xj9yewDkvMfCrBSC9rj7kNdfLZ
0gaqxnVaidwpMo2eUsBbQp5A43DNGQAnW+C3Syhz4OvZHjaaUtK4cpr3Kv5kpVo5
eanQZJfVwhhX5zEd/XbqLEsbFF0x6lBP+7QcEgeSMAOpBWsxYfTWoQM9D5kKuzwR
k54Tu+QdEYb6ZbH1vlLUhBgUSofbHX8a+TPUdZ2D6Zp9rkiKyny2TzXg8p4PLd4E
1MP2ezXkEusy/a0wJbopjs1AbVJ8R4RgQUIjLUHDGbBtR2BE9e9cxxtqntOUnKaG
bN/uZ8Q1zjt8jCwRKzNz70lxtQK/KkF8FHYIH/0bfwRBcMpth1vBqby2yh69I7rq
Gbmflr5KiVK/Lzny192ca21mzCfIeSDxS5dyFUpgnPj8uFomjHFdjrde/loecSRA
N4CQJ+NClXm8Nbr+zxn4r34efVolqa8cIFvf/C/R67S1UZElSpKS8aqFzoOpas52
CclYA+8pap8dvdJ20E7LGsvQc89HIkyQSEMlDzmqsr1JmLQCv5fDHrkmHnqXd9eh
TZGcIFEslDZRx1yj/Lum+arl7/1i6PDhuHpGE5IEvZ+Lt4IotqXpUfdcVfeHkMqB
NzqMKkx2ogsZ8d7fcNatzkPZV2kniIf5f6FoFdR4TbIJNa4hKrLvXcFf1YcBFX4a
4Z5ZTN3FO4sPvnf+Xo3TqTWn+P3nap3wzQrsWqyweoz4yyoVeRHXQbb9XWgIM8h+
27J25ZjJ48UVncAOCxPwJGjTq8p3sx6XGgwrzu0L7QYLQFYW46cTAlj9QqSP03+x
SH6Bgd9BSY2+9OlN4Yk48YBVAwLlsUPeMfKBhdTNGcJJ8iA44Frdu5lUGjKzjXFg
CTwia2iGoZnSNOD66Odwch8Nje7fYj3CyFC32vrZy2OEoqJttsOMjEKOGdSNHnJ2
aTE+RjkhssCxxjN/sxr769Cps1j/IlG3xQZC2H6m/i/p94qUPHzHVeRj8e/3uih8
BxtIs8Gr/xeODy7cHMUdYhV7PKoR0YNGd8T8QQUZuy8QHNbTVNTOnQjlu1fMINlf
mCjZgdjbI00M45HQh/CIwQZsGsnD1sgrty9jns4OYPNMUUXPDK3cfe2QWZ2Gx/2q
jaNgogIfYJPp210fHn3E/yBMRryScDQXLkyEYL2AlFqu+2CZM2SIor7/4/M6SoxY
kFS8QRF6IyRsGveH1Ic7mimsRnrND16ReHEcfnWPweldrXeTuiEnlAOJVEcVgKuS
dqQdVp2Fyp1m2xCW8i2n4MIhQLypfAm1bXoHaGOm2uqVY/1UZMOhOcWBXalKEvYJ
KyHwUfPAEmzaWB0fJTcXoSUqBWjK6hcNwkQ7Lquvo0gsy65/exkWkRZPybd1BA5j
9LURJAmybGCrt4xApgMUWlap0exqzxN+0fjz8liG5ctSyjWWBHQUAxqnBJ9cdL42
OjZ/LKkkzOIjLg4wMJBMjPOM+KJC9ImHEJYJcWDJEXdl8rabmzqaB1MeVj+vcay0
FBvp9A5gPSZycGtF0B+dRP8QRdWpfU4XVbW59rH9IvsPXihAYq7qbrJyMQSkZvC8
IJ6eoMF4VdmWkBC3d9fGnCdob1CrARVGlUx44HMe6BVV1h0sUbVw1sGXYaKRLIOV
juRoSBId/NMiaOQxWqyClxxO8TzjJ4qq4H0I+EaE95ztzRkCdLhVF0j70mqpR4/0
AWaaSsiWGXtZu8bGjtppp+yrVrlRnaXw0hA7+sp52WQPK7jn7yAOykldEp09jXFu
sC+LOR0KjRW7tKeAJ4kwP5UD8O6jvJSkKwC19A5ng0YCsqDYL7guTY86voWoYpOX
zNwXJLeE2BaZIZuHzGYXqLewy6Uq1Ns4ItjsQxSe2FulZiQINngdt67LbY6qVlDh
iU+vSb0vhmH1bO/IlnGcVyf/hS7spVSK7fg0BXCOYpivyhES8UL5RqXv6ujwQft1
leES75OGQJ+V0eQhbqb0cyvUccmYcu810AMZbW28S6JW3Xo/IcnYPcCCScpdn72A
plS8QhryggfSgJuBLAAZcqSDKAtzjVjY4xnx+cWPWA1cOgID5zERZ2PT3yGm0k1a
s0XoV35x5gSlBoT5Ej0vBwEQCzz138or62OZEuLiu6RDHYMos86603kqRGlFttSh
JR8ybrKBLTBDaYrO4uiNGRjLygfbpCbXFjprm7eQTLnRqkvJ8dthijZFzMErFlP/
6YPdFnMJOlOiErF14mpnblL2FKaDoCln525VVOuVn4PgkHNNWv0lTp6cfGD9cEtU
CvVG1u7dNl2yMbjiMBAoMb1am7GX0pOKjgHc6S7lV6YEFWRrH0MXsWbAKlJeiMOQ
MUsd+ddOaMYhMECgoU2ubdyAVjTKYpy3+QE1UO3ARWm8tzO5atoVhF1OTXNGVJe7
X+8oTpc9EQFk+MH1vBgPRFajpmOuzV3ZOv8WRrtuA+nITEqY41SZmMIuDgyt1+tI
2q9n3YR3hAvW1FRIMaEr2AeC9nxx/cC4Tx0ayTm8hbvxLwycPl/i9uiMnYploAiJ
HBUaw2inwLsVd28/dF3E3xDK9m+UNm20WNg4qr6dqKV7uISAu4Wxh7MugHqst+TF
eYVkrd5JRn/rUbshVNjey5Z+GbZDFuVKekXoX2oP8/k1OrmUFFko7K66DmIjR4Ud
5E6USB8Kk23XibTdFHbPR93goC/4v3MTo0MUsLaLZze+d1B4ZW8bDb8TVK0F77QO
0KXJPEzkC/fOdHEoRZoBEd/17lcIRv8F0E3CPAMWRHlTFxbaVk2x94RGNPR0gEY5
ixdJnVODYhuphBQcBCGAYXIQ3fpTJKtROx1MTXVXzNvB0OtctU1FwgyT/ep8lLUK
l5PEmf7lRKRLPN08kpTYHjLdsLCkYhxpB1h9uoKjZP0ZmGWpc166d9BnN9R3aCjq
kKKkFHRSvmvibf2vvf01mqR1TpA9L4v361fBc7yZl4jkkqQQSf9m+gocK36Q4gmy
ThahYG1mhopKS3BFnadGtnTzhwJ+xHmZCzuzXsBMQYprNHWaO/NJQsMfPpS8p1Cz
BqQjXokvjWP0EHibu+rzjRR8IndWo6KZZXdz/Y8DlF9ORRkqTVnTCjGAH4i3TWJ/
3lwA7wr8kGC0sQRhM2Y7zEUDQJCAlXk67LWAJETA/xm3Uv73zZ/ESXqM8lrL1a//
scuLsAZzlauZW8F9romsV/cz6ArwDqpF29mAH9I5GOZerla5N7d6rhuqyfJHAnzG
S6+iP1sTukT2ErLSBgT+D7luf2XXauAAWichgDxONqy4WrDBwX4J22eHfN/Cv+UI
EH5SBSg9rjPThjH9cEkwDmslOhDtO6J221LQNZ/ghwn1QreLwr4BSLbOFLoDRa1i
ChaNsDsRNP8CPhNhgvnnjlaLhFJtdFaAID5zDtzAg33VlrWsoYrRn3bbOGL5gi8g
H/Z6Orv21ff034aeTKAUAY2mVX4N1VwgEqFVwb85RPh/2CpbHOgdPzixIhWFJMRU
xiM9NkilzJaaVC6nWHuXeoGxF+DnlYpmaFt8Cj/qPqOl2/3Md5uU+YRMQHwRgVwD
sjDCdgPJRHyj5ScJMiZisaITRduNXHIWcNK5ryP3QCgwkORLCysEQ4v5vJSTCdvc
xUT/bSvqDRAvHt/+gss69lfk6jsUqasABhxvfUD+NBXi84toYyYoO1QW1nHkWmx8
4Oz4JUZDs2TPTKbS1Dn3Csy6Ii1jQLHFPjnPftohLK9xwEGHY6qA/aVSdX7IXhzG
Ie9ORdpAW3w2tAmD13VOtID9iKXpPS1BU8bbuMbeElqJApSyE+abhqJSnXYPcToy
DApVUXeTBhLomw4Nk+J6pe1f95Aztap2bIPNq/uOfGx/SDU1G/0I6QpaQMBna2xA
OZOqPPzIEuSkQMktkNcldfKtjEtbopDkPW6feYr2bv2/ggMYYSYnkbKD/NzkFebB
0poeBd4MoWn38r60PpAX0g3gd5n2yOodhT/0hjFOsgKvk3DNQB5vYTDxzm9L+kiz
avd+Gf04ORTwzuEi7jTif9O9yp7FI2BFZ0/oTMpTCBUgHa73bC6Xr3DbZ0ll3OSs
LGwpzQNcYSqj2IbmzySZ3IOF130E7CFF4Jj/SsTcLUh/iXD9eO3M1/k3LfpVkl8p
2BgqWJ4IzVvCT6Jlpt8wUQYby6U8W2gWkNNiSfQGbBB3dQEktdpB2FpFCU6FJepo
Yr+uauy5xB1u4G8aQvRI4NTa9B9Wu1e5PALSFLV59asAdTGPxSzrcxutFkbapcja
tg8jyEaEepgePlu3V9MQ1XSb3AStwQfF2NeNaZtL6VftrKWNTiM51FCiQOS5Lhap
VRv/klalS/uin6pqzwKTLTGxZB9+YdkwUlv9r1v/H9nqKZNx4xKiE3KmejoKHvHN
a99wFPxH023LrnHD11P03OS/xmbPZ/H4FuCCotUt7MK4Urda56YkRhxVAALPdLOb
onHm1KVp6GxJWhPsLupjXfuUxSLe+otKW6KKM0EW76PzXT/+QB1M0pvz+uUIzenD
J0uP2CgUgazjoZRhVcMRpMqwk8mMzDN+eGYQwvuVpZbs1k7GZgOhahd+NU0VSzD7
hCitOxgndK5GBa8ALNF0COEd4dk3dD006SKdAfdpYgUtYvEGDQ63nlhNDUBI3sg2
Pnt3M2guyF1Ei37h3yFfh6TjgeCvcETRPvqb/b6CvAX/TFLhgtGjKtHyaGnCdSK0
59zdWCPnPZ0Gu+OUqNnIU7E3J5FSZmdq2EX46Oy1ATEK9G41yPBShcrr2bFDjwtX
voATpvES8T3PyrhBgGWEUWtkbmGLKFCmRYlf+mzAzCifvhQpaA20F8JI5Gt7U+CH
y2eSYua9tZnkKhx7D1T1DsbQrG4jSMrZjzZHUHs3S7H/H8fD2NdGV8N9JFDvpzWf
+rwEDdyJt1x2Wrqp1tDw5a3QP292WBO33eXrL64vqAWZGBz+10PEHzQekTpWLOEN
i8Srwyo8/ENnMW5Zv3JkOSoW0LW42GS7ZMGK7sR6YVtjqKDwcibb/OuPfVCUxmQM
FEGVQgUz42YbyZIPEmpkQgZRGhNTdVo07WbE0W6KIhxBp9JImOA7ZE2rZ2kY37T5
fnOUTHAnsX3r27koMixZYSdx8Z6kY3DTbd7/ylE14rMrbAq6th1HiRbYMhd3O4GE
gbCkawPwYCE1j63qvMH5x+d6wudYyYSv89sVNH+I8zvafFhg2eI5hsiRAAUoOslK
U88rxyith94FX5wMbqbw8uXMJXzS247ZLIYzFx6WLGDNaeDnZ/ravoJ7ElIUS8E4
dbb9tJ6wUDBFteRKJr3lSLFqj1xMdd4j3LogZYjPfW1nZjyFs61CaNH51RE3XRcT
Nq6cbGckiI3lbnU2iy1VYwXQUgYrpuAoEAXjZ1hzbkGAiM9yckbRNd7RSaToZhEB
yY0Lu6ojlmgVwaEl9aG+yN4ahAmI3gqmX0rIURFhA7HrrNZ6DAbwGpLeMcmkC5AF
b9y7X81kfHMRPdmN/kFL0Wpgdh3ZJnyZrPplGfNcja5UzMbJChnlne5/2MH0Sc7G
4QLjaT7dfpQE/rA5Tks5+DKMr86dpHf+lzv4czwR7D2O8pEVYi9B+YSXb2HLwbZw
sDGK6rFOrII+xO4H2Ak/OnZqHjAty1F3QLdKVz9aEkvDyd4hRqrgUfEZxXxwuwi+
9SErQ/U+YUXhEBvIjP9GKYpRdDcCWHjfHe7ZyMUSlgYv4zTKgjMI+8iEgQRsABKB
ULZnelCEqE4P8v5Z7gEPS9wTbhzuPVI96mPB3A4Iero6FShlzG9zs42X1UjCtMNE
fq/THtGAXH2sJlI/0L49sHqzoH+0zjpQWrIoV5JRjJCk45EVeUoHsd23qkzQW+nE
CnXACSnuAoeMUYdBMsAT3C4W5Y3ilRvOIXXS0SHKNq2zOXr0OBCFrYt9OUlRIBdf
mQtv43eEG7kvADLxE4KS3elPhEPV9Ew/3IKBkaeYws0K9Z0WmcA9ost3hlQahHQh
fRAfA5+SkK+mc1vA727ei7QHCpLTlTwdAr5tjQxb3qB/CTZdKnbfp89SZsCOfoad
8uhiAZ9CkBEODCclUaI/pdmON3e0QAwc4B23YSkFStm6G7s8Vgx+hLv0h/O8yCF5
QyFkf46zbZc5aMxIsy3dXMmmeHjgpO72W93+1EInY8EFLoTCz6xitDWg+RIhIAjS
dCGJmvbgKB7faBCrT76t6yRz7zv0vE5pOqxvOpKqb931RP19e08oDxmL5z00SXGH
LctgI9FhpvEY65lqzNwhQbKBj0aJDesCwkvRvsEkzDjrfjlM11lV+/GIyozUVfUU
4tANdRxMp8bjIGqck5DRziVI6TKYZ+4BokbQ6vqxqb5qqQU49q8nlsnLWK8wfp+6
Zt83uxM+9ntsRklxz0tZ/W0G/Ucfbzo2x4V5mD3XtEBIhNCWHqMQ0SjYAYE29Tnh
YUlHi6PZ/vjrb/eAHaC8w1S+6ArA2bC8kuw0cDBYNOEX7Lr01KgNIkWBK1I4ulIw
9HJgVB/eaIM6VtBGowa/X/boSzmDyaZWHa1MNAaYwJz0SedrVC5v6KMOoyaeQLpU
KF380GIo3MX1HOBwlqDVXIajBQsVDyfrdv50tK52rILD7KBMkfZfUEOVV5zL9Lhj
eYZykdalzCYkASDXVdPn+Z9O7nScNs5dHi71k1mdiyX2JtgwhlC7q0hgLLwM1xT4
GxEkVD132QgacsVM4wK8OBLSYQjZWyVP0nNGTc0u6GR/lZ1HZ3cUCbMIuSWhw8ZC
G9J/lOYSfcgIfe6DRHI7v8g821aiSosopiU81EHrAMUiQcaA59PZGoBAvbA0xRcc
va4EAjjb5WlWfn1IRfbyMmy3yrGc2ZFZgygumeFd5jQOVFIxWGNYec6jCf6KDgPF
g+jaDzEJE3gnTQE1aZYJFGkR/DMM+pxyLogjckDynonvA++qyktyi4Fc3J4wjFk4
p6ychChP+7uRhyHiE3aOovyMhjpC1Ji3dhDioc4qTJvDyfcqgZHeJj1hive9922+
hDsDoKE0Ij9iN3szdU3S5VxsClP5gvuwV/zdn+8ldEWMh2lW3SaMk8xwYYSaVe/2
h5GdBgLexlRyinZh1ndjcG3Y1pEyp7i5kKC9GLm377O7jvzHu4baa/64Hd5t0BVE
pgLDzSgeRo4UAWcMtkrsbPioZkHsBq8+JI8cB0UsppS5RjKMGQLQqMfqGPuZ5Gpv
fpvA4wV8f46dhgIbfItJIDvZISHWECXVM8BXRsbbPev5QUqTtqeNSCWFVFSt050J
CfCO1L0saR9ThkuoGt2G9xHAQFKGCc+M57GVjo+zdL3OBgLC9cKEJkyFtodXPgZo
boKnkUaYnwsYbAig6eXrfcZiq4q/4mJCGRGa54PEex+B43d1fnSX++5LqxnUa7cp
2IQk1BJSoUtdivW1ekvTXoZvkdqpi1yf+ntNPGKwKCK8nrWwdpVbzfYy4avhEciK
A1APJ3HwgXknQXAbnWHDttuujst0LDHX2DFM5++GLbEHpjDKSL8GotDRxwATIeOX
dxf8nFqPYl72d9bCGsqkmMWbLewq/FXRewznTFVp3w6ILloBSXMotaJhNnpo8L75
k/WHTtKz/hu8xQfbQ/XqX2d0nMHhDWcTkDffwZeOqA/pDOL8s7OQF1SqgNHDUwkc
TFrjhy9R/2W7ayRBhkvz8wkuoFsF5r8dnzAp/M+vFyMB1c7wpwq/ID6payAf2T7k
orYSkTPEtvZlTS768dk3FXBMos2eAAkt5Hwoea1DyjnVK1TSB4iujz5krevYlE7p
Um55Qh89vj9o8GWTGRaF+8zaEfhQtTZgvEx+pCmWkQ5sUqDSgVF5gZRoqYkQize1
Ye79uoZaNlGkDGD9SuJMd5r9+ZIRunzPpWuf2+QveeF5pANRpKsBUEQPaCYxWtH5
rgA/3nSROK0jiGn/XIz7ZJT4J6WWA8R2p8OPgRH+q/hKX20TUQV9ULb/kdQlW+Ic
8JuFxP5b80QCSZbd8gqY2KY1ioAyrQ1An/mU8dShYpoqr9mb6YrCKEmKSac5uVVS
bv9JavjGATW6SnvNG+FImmPtU86+wPaJTELm5LEmsAZg9VH1GE9swkwW1K25Ag4D
wSQHAQQDKkPx/qwummtp8xZ+z+DUe1rM7WL6/23utSrEP/yAfujtuDu0fjbCMl9u
IhWSPiNCG7Yv7lUBwI0Glhzrj80jfvGf6+kpQL2KIgzoGT3gL9T2uOSEn1bUY8rf
ZsI3jp+GHstd3bWhY5eTJmNuSJg0xaIZGJYxP43WFGoqcTsi9sn+kYVtepVD5qZw
pbH3123R7/CZ+unQEwCJ8aOkvoDp2QnOSKwAbnzVrxYjP4mVUAqUaZF/EOGdfOio
a5vSNvUQA8G/B78Syn2uwbzqig1HXT+YzET0fIzUsRS73mT2MTkE9/ZsezMx9fBv
XNpb1sjme8RnwCCxhPEVHcaQHApOfXZAJimzeRsb6HM/LI6tv8DoLcCGLy2DrVDn
EIQavffLIeilqG9kI49er9hKbQ9kyP1IssC+IetDpBzZgXbCFrw/ojK20V5H1xed
RA2NB+wGAq0hHT+tLNh4GAZOUlZusfQQBn4mOj2DJ4qCJutwlPS6c3whMs+wXf/L
axaxsrhVjTMKC9UNeb4Rnk0Omah9UVNLxls9WoYUXAIWUEQZA13uJGgJ4sIcAK7W
wvK1QpScF+UwaGmUOnHjFzG6bP2VVY0/bq8WZ2NeSfrv0xTCNv183Ed8HU5sxCqT
XEdkhdxpyYsAuBoxBp3ALxM3Nh3o0Keqc1mGQGIRV3JF+X7olntxORIbbU3Rnnhb
Hx7jlURNoKNmwn1d1YU1aDnNBOGu7+9Q1qQcg33bYUK/oWhrS5owrhK0oECjb+B0
3FbL4Fxa6ksm/m6HEnnJCx0Qm5lHwRfty06p9dNDYs4P+5rSkh9IaLRA8FlrRQQa
myAiXW9nSv4xF1SXe48dMLKZnQH7EcLN7WYFlWTy3CUO08ZsUijYZCPmGSoXE//A
q9RPt4nkYAE6ohbNQrMl6bz1/sajG35P4Ofgm6GkJoqDmOMy61QrFMjgzfgPTh3H
2hPeYuhF2IfPM1Cq8FE2PoEBClkSYQpmXlZtXVXCRdfMdz2E6SlBv7U/eRuYtjl/
+mkBh0Y4/9WdN+aY7t1bMT8hqQtgCBsSW1uX1FYHsoY1uXZecWsVdcwblLyBfMNa
Ifzlpm8gJ14APglP5GkssEAkYfGYHl8vcFOi3gg0p9DNgA51wv0+5IGO/Y6g2vF7
X5QLN9XI9fF2QrPbMryKsedh3dSjoH3GtSLyJyeDpAGd0pec7oYlubkI0kCZr4hg
lwyBH+xy7no7gHNCYuZVUe59gNwEXx5ixHjUQrS0YB7vnvBrKQqcZ3UmZ0+gn1ze
d6w/14GUg7yp/w7KFTEo37sU+tfb/dhnONNkOHugTIDtKFQlF2dwDRyOaks9zJ6L
K57WFyG8DHqNfySKvQOkDCmWLbqJkHd4zg17O8HZfiIA6ApbztuLNz+2CtCg6G/o
ufnymLdqQ0WppSrlEPvbpQAQVsco9htot4ZddnnlDK2Ctx+Yl92+RWxLX9z4z+Gd
zL3RDsrc1nhPU7v7wmJEJ+XdeNccqtWmotdbCUm46IiOuwS5xuNf96pMhA3ueOoF
cSCiZUlp3AwjSHsXQ6CsCroqd/1q3ZaWfBs4j8U0yRIiLvkwhTHcW9wKEVhiPyKQ
ZJpGxKxhGtt5EdDd3qDgVdtmP3sQdISJSFPKEXSQ1iUHHzBw4L+iXfbIxCeTiuhT
HMagZzItqVJohQVl9EGJHKD5b9s7wWj7h4Mj5qMnl4XXk9bPsHlxPHt56eaI1euK
lB1vcsG4vWd8tyGyj85vMSHDWU7Z59OYb7WMecCbKvmrkplelOUa6CYwLgaZ1Dsj
jamOTCVoZy4FvZO8EDwgBsCDrwm6H057cEI/+45e2Pltwx91sWq7B22FHxrEHnLr
LTcXYECAUlZhXRdORqU7fCMjwyTptiGnZRrTBq0SjwGD1ita1C851aiWmEvGNTfd
BOOWCaUaEnZGa5XqT8FgxIUiUt0JE+EvPF1csXLGOTRHUAPTlQPm/48sqKhdzvEO
lWgCWZM6NhIbVO3LhLeX5bH8neWHkYJn0mNmKiqsxqBuPHbSJE5jJTiGqIQnN5gd
VOOb7NTNWBVpDI52yiYBS1ILmMHLj+/l44maWW/maEsfdo0aBuTIZ3aQJ0zSFP5g
fzE6KTqlwC5qTzmUOcnNeJRKDGk3WmSpdPyaD0yQLgFWG14XDkmXi4fhjfYa7YTz
Z/YpL1GWAeNc2FmT6GX3/15G8dhff3Ex9W+HBc0NGfGdZyqKCIau77Q6HgY9YMFB
LqVRE4y14etQ7l5A8LFXGua/wYofH/dxJcyGLKpQFQrWm5jUXzz+2/X7aL8gsFk1
iUXShw4F7NtjWSMqH6LkMks1R42yxUnqofo31s4Rv6Kc8m71/B9WU0D/Fa5Avgol
qV05g4wbKGJNXA2+iTrqB6oBIeANCTMydoFrOVkEf93FHTfATrqP6ZsOZNIaJrbT
Tj5YS7ibvg9gtrnHeicLebfS7kZfXhf3JcEF/gFp2Y2+C1VO+7Qthv8RUiWjYop/
ntxoOt9FuNqunY64OMKO/Pxhntm/pXxdQDahx2CMEOLTHJMewW4zArYFl8JUBier
dapoHcHgfvep+gsDxP/2on9t6G3DqjI/Ga1W3Z3cLIFODssqONLJ4Bn1yCS+H8o3
Yi6jMspF1QHr0r0d2KIhtvMSQL8jbej28Q6uzP0vD0vvhGefTx8IPX74g0USbE0a
rd/PV9PLDpro/HBu7VhVzwiVq+c4BlpayPW0+JdkGBxaobFOdMkP0jwND369Xs3H
cKxyzj4t0uRy/MasM2v4lIwlaZflu4dZYR5Ylk2lBHsputc/IczvmYTMM07/jTST
JhzC8FE1ILYq5S4DuBTsrpRBIQsfOuSln+sZ6qY3vjdIKxKr2JIPlFCMdOTiy3KS
iZqdUqsBIefO0ygAjCjYeF1k4PTSUtd21p4aAhIYITikcw/mb1JWQIUCYk8xsmjC
GMNQ8QpzQ+uHPaYR/ELIc2fe4tc85yMzar8XoWdakLZjQKm6ged8LOR077RTfIvT
sj48e2FD6aLOxgzoBEw7ouc3v+1Zuurrl6dCr6IYuE1IXBDKCQBvNi81MPRK5I7N
swgJhLLirTvOp/FtMTY0SdQGeY/M2ClxNISRlJCnfWYXGIbkw5Lm4FO67kNpqsas
UU86nlShUItN49BjZwzQzMivyxXo4xuK1QQ8F2hJqMNx2tAzeN0mUmeOoQqb2tUV
cQspqbIGVvOyWlO1HbeaHtIUCSnzXvbodzadJz+1E8W9fYHQTNAxyJMJccml9nP5
dklTcxmn420xe2NboxLSCNdKisnwDU2Kn29pnEN46cItdDIyP7tY0V28IFkll+vx
LKl6YCvWZjQJeEOlkuunoGNp0ioCFHXvDBERjEg7HwRnvSEBPWg4WrZqHSdOXgrq
lSrgyhIvqJ+lsRMWR4SAxkrwhnkDEmlOPZdW8574H8rZJdW1IYjtHAWa3yd6LNYP
F1kX8WEOZsortb7QcOHMAB7JqiMEdlQApCwWPeKboO+3jZtpUNmwlPB5gTuFxrpj
PJnfS2cSUvwH62ZzltJqmEkSDiZiUPAqN6j+79/AAVdjf543ZyRmS3bGZhN8EovE
MwUgf7wu5lrrmIi/Q3AT1THejVSsVcKkL3KSTrkYs8uIvxujn3Lt+9G0GR53bYPn
I1Q5tQjvhSXGtSHwa6RYAGIBuuQLFGyvNTpc364P6BFqU25yrn/7du0IM2VOBOMg
MnpCaII7E6yXYviK/PsHsOLuttre0RIXVAlCWJXAHCpX+2IjeSHx2r+uL1e35kIF
/aqSyIZI9dgrhfPNyoFreKpD/9BjFv40L1D+oHZz3z90R2DFYrdMqJ/LDJrultxh
9kmAuDxEmI3JObyk49qEbGDf8mGKEBDjdU2EsONmvCJOlOtEf1bGzwQQwLWDF2rc
fVgbNK0OkQniljhoXDsRnip7Vm+0EPVP4Kcc2h4xWoPkyC+Zh4Ej+QvFjHBoHTsq
JoGhuwCFO8vHKCS3cmdXDmML5CGSraUE8sz0z69D5mp1wRmOKrDqJfyD2Tqie4MQ
pwwmdX9FEZoCXXdurrNzDWP9OtNl0gIPESTka/783MbcfWXSCv5gImJWJ/5gAonT
Srmq7ll9EDxxjq/gQmp+DLu9DrUT/OE8Y3AIT8NOMcs/W+I2xdamEDzgYAeXgTtk
nfiixQeUG6JdxsmWNBf5a4YW3Jm7XG19TEEekIMfYbNmSvIAHN+l2k49CqP4eZBO
0uLsY5EhSQ354SybUAFh6n7mmOMd+hhOpnSiSsDs85wjh1kCzYN9sMq2mwnAjX9B
6BiiV5YRwFOv4Dhg5nlfxNvSjf6pI+T14ggw827heTRsdt1WQjcyYIxXGu6wXOs8
qlDEXS/fKG7q1oxPsobJeo3kc3X17Tjlr7FrSQzlQluIl6fg44FQ2cSQSudlivSG
QslaI2NMp4dyUQJHEIg5eKih31Xc4kBzo0v8VgpZ2hxrNuZPJ69FLZxiQF5EPKRR
VVGqu2z/gUqhLR/x3iGsSSwD3wqV4Ds4/oAB7J7hC5SIl2+FBqvyV4/NCRnv+/Zh
rK5+QYmyyYSFsm7R+vWQx7w9d8PC/OD1+VVQvHZXusZAz9L1ic6aUHwpgD5pnzmz
BpRI1oOPZrZTCWKEPOUM0J7kBeR8kBFTGavqFbKLhj4LiaJQzp4iu2l1j084Bo+8
w6ryN79Qev7H08FyaNXo6i+PqmPxQKF7DsQMoPJ/9oBlapua44PSCNJ0xtDzRb09
CtLofwY3kn3OsRV7q9X/ENqu44/4jlJkI3jPrWy2BlgiLlcFEIyvCJQA/Z9PJR0s
OeT5rXt+rkInVBGzeQq2DRcABI3pRp/vn3eXyS4stdJDbthRPjjMGEQXl5dJ8UF6
VQprQdnFYJX6uWZgQPSAiEszyEH8EHBdYfhnAK6cfkeUkJxK61roKJY9MTPgp8Q3
gONG3Uy9PboL7YVt/IScJE00KwGA3paojACDLKXjmS8bmytc9AKbggyF4qPoizbP
3noZbZWsfdJdqZdro5b0FmLF5jagkm7EHwoOYwULqmaJYxZr8DAGzdMM8+4mAGl8
UeUI1dvXu9aOuJeik8bjXEB3wIDQebz/ebikbSdeulW1eG/ERz+HBnOZXGFrzbnx
UziCZZVmq8aWkm7180edZoUGPgsatc0mYkssIaOBggeYC98LzXmHV7Uo71XH8Vh0
AWX0FQ/8FWWiDQzYGqmWcYlMzRkRKXXU+v4zsrjebHArQuEqG7LrLoKDJEvfiN1I
il9mjEvPox9bxvDdvqW4ohK8dlTwk2Rx7UezXAbsheuWiA9AeU5dcD9iCkN6wXem
iYpJPu2nCR1NclZuYYkDCf3KxYk7NqjAxtfLXAXbIwsp5E2cHpDA4lbkVE8H3O0F
L8hKuV5rknF0Nwj9jnRvxOngCat/5Uij5WA5brC/42EbVWUrGNbvFBeqS20NM694
EAOGSx+si3uMCUbRA+ZeTICksY6hEGhn/AxKo2/wRMtYY0wC8pCkTGJLn5R3mwnK
RLZHGZLjP/azt1La4LQ+5kMrvGEB0XXvETdcsyfEop4VTv+DbvlsZIz/NWNxnR/H
Rw5/0GvfM99+v4orgSdFhL3bQn0yR2CtxirEyHkzDNzLofV9UmKD9BCjUB9oxarS
NL16A3Z7PeplnDrlL/1ZkOxtYGmlIWqyLZ3/dlMa+WTy/krJmac9GvE2Vcmoz3TT
u5UjY9d8SKKdV9mqJniMwvYzuUh4wj7IoDe/tZYbzzEcztuZpozPtttI/fMFBTCk
MR4yrtwUGTl3HC1oBRdSabjHJDPc2r6hcv21i9Ijbg3LphHhCRxgzEUpu7W3Yo/A
CY1qIvsJDiv04lTv0gbprKvUhvOA0OHassjPUdWG8IGdMngp30mZceYJ5iBlBEbr
HlDYS0T2mHoMK+tjyzeLNDC0sczV2TZSkCPBZ8ksyN5RmrtmIZ8fC4gipdV5xRAD
Xk1ntvikeqyehSyX793zvctMjPcX/Bi+UbAfjoL6xwYLtHnexj5uCruAVk4MmqCQ
J7ZPhRQ/Ei9uNJCDz+tZJzMB4CquYVW0/i2aDWCMUTiOLiWzzUSh5f2K61VCwqAB
dAnytK49M7t4Q2G9V+KeyIJw+OkHtbGP15+ZaOsVRVb+OjXCQwtky1EPhxvUq+q5
Omgrs6CaxBssiy3++qU12lnwrzZ5ACjCP5W3elxmT7vH6510jV81U91b3F4jyn/U
3iavfCXHM62e5RaKsE/meC4xP3/QS5KFBwFuw23ijju2+BirqF+xzqlJ5XRKSR0m
W9RRbbCf3+ucwWtimSZVdsBu4wnqYa5PUnp+HjrXLL6P6MKspbBLeZm6dxk1d+ai
Dsfm7ldPdb2RxGQTPkNvPqwXWHiS9OLSJRzYYAu3Ixjpq2yDU2vvjRJBEmOJIz0C
7NtfwEujL6s9Itx0k3TQKCMKK+SAqLKhZyING+AHIIkF3P+VFt/quOyCcUPZbyjt
5GCFimLqSqUaS01IeWKNCspzoIiY7qIBzSeuYUC2hjw2BVLnoJIco9/MSq8+2+5t
A2MUUFCT1T7kmNvH8DYVzzGwF2DcN0Dw4G223vskA2GQFqPNLV4vFvZJg4ZIoxzO
osOhQ3JoX2VHOrzMCSOkPt26Lw44oqLj05iZpvo8NJlwkwBu2/R/5bZ+wWt++p0j
j1MYWaxz3UbzSKq2K7b7CcX9zvE14If3MjDnMoAVBOfBe6jZt8MTbo6P5tNaz8QA
RtzQMEhNNFYWkqU4SUCaiQDXRdI8t+YoUhGTvb2yKgbdIe6dvLQb0MusJtvW+3Sg
HieFuAoQyJazN27CnbZCePam9ohnr7UIfJg3buN/Z0dpW+pjcrENCZhNRb1BBJoQ
pYv/b3bGNB/9W0a4Eill0gF70htKF1fqeEhoUCcA8YRHvW1fFJBBlCgHS4YB5Ear
7XaWKK8THy4lMFkBryJO2UZuTtMyJ018oz1oOFtZClcO6FpbtEYel4zIrIc0OEDZ
PW/6hINo3g0O53iZlE7WUNsJq/6PuvEdYLvFtJL+rpjhX1zOjDjwcYbIcBAQDUhw
LnDnw9TBXmVmEn6bMME6rbdojHLuBg+o8BcEJ+sAww2Vey9+snjui7+Rsr+xghAF
BZH0TWLg4Yo1tW7xhLYz8uEiNi+4FXrelQzeh1VQn4/1b+bi1Rjw0oItmEBQKL6L
8JCF+v7OoURPyzv17gq+GbL9qDhKZv6+rPqdD8XP/56CmzYADRYHyOj+mE+3ZQu6
FbWAFy08aTy2qBw/2sdvwMh5xOlQsAIlDGgbmnblG+VdgamLa6YgGfisny0rT8ML
0iF/rSWkQTCbqM7dn6hMax8UOz0N46vIEPIwGvgqq/B9ErQ6T5/HNCbP151UnvpK
fsBGMAHSJuwKMo6Eu9y7OFzNJAPswqOZM5fKIANMCOPVcFGT84VjH7zwyKK9Av5s
etYFnH7TTlTuoBylyPgEDu3q81isEOsQn0GVRZDZgoZakSqfdZ1gSTAiB3M7f1H5
Ksa+6luX6/+M6Dv2bpQeH8Q2i61nCMLDqoIJm+IUIzUgda/FznBzymm8u/ZJ/9a3
L647L91IXV9FkI1AYcR+6mBWHS2gXvh70t/XUxWfW9U0ILk9xBBGymfGx0qHlL/A
MLz4E3GV0Q9F3FQ6yUa/AfhhY40FnJN4Z0nwrmaW1wB2q4HyjEJze0Gm2c4Tb1B5
YPJBQjUG0PAps2JVBcEOL9tocFytMXL0uRneLfd/bFot+iqlLmmdF/EItUs8o7mD
JGfE/BrBtR6AFB2G/KoWZL3Q2CqTDOotcL9XiVTszEelHthbOMzKkcjU/8o+cl04
CHKf7VTNxn03wS2fyx99fgx9gDP4pT1+rz7Ycw1sG9FWymJkJn312Y4C+ZkcgJq7
0+UJ1YIHfTEcgG4N/KshPQpSjWa01FE+dRjYQA09frcnpp1xyhWEhqltXGZe17iD
lZFqYby8KMbZBeHNnbmRDPA0HDQsp6Um75qiFQB4259brB1D7eumpcZ3bg+mAbiX
OfHPCMTY2epsqrq9b6o6rEpGdBRsP+q1OUTKuBB+l8sp2PnhMzpRcMDEirTnCadO
qIVwtvDz6u6mz8Snb20GP+yoSS4h188xbYRU7bGDt+8aZNcR5Nb3crdMN/mUmlGE
+WkgKejqREUVeEUaa7CnaaiCu0M0i0E4gYrbD30Oynx/ifHkDt55l8BnxV2DYLv7
/eObIt0qdLTjxWY2G/du3l8WZWdFYD2pmOtMqF8Ad1ZLFniQQGFaLqGk6+Ismozj
6GpkT+9BZ8bK6AmL1korpkWOzYG2QGIkyi/tywzr+jtLgLn8yJ4vSBU46uUwz/fp
XArv2diLyXz1r1IHz8GtjP0IUC4wTJVfjIcP2Yb9hrfT6Gv2k9GwnZ/dkPTdE2Kl
mTNFM7dq3bIpYx2lA0TVJ1/7NzI0144kZPO0LMeq6NUhizxuE9gKu1x88nzRjs9l
NLHT4YYMSc3Bb+vKv/zu4oBAzk0ugxHIp9eHtXbUIIsp9IWSm+NsGl154VuFhWTG
x49PtSzWfhecHl2sLIjIlQ49c8nm0sZYahFoO5LfKva/jQ0w/OqCvuPfVdBFTaYf
YA7+ZaiMZyDmHknszToMc48vfagUt1oJrktqrnOJsk0CPxNLMGewU7OTb0wSHhqH
HQVTSaJmq0fHyok6VO70UR00Cxt1meugXTVgSEqE15LuPuvwjAc35tKKMYvc9arU
Ktm0K12tkUDOnX64DMrk0oZHLfAOfCwU1k+F/oyZRFWbCijcl4WTbNx/hquns6JV
AkUGSqVqC04dynBQkC6UU6PsCHcJqPZKzTDn/BWdcJpbdRNIEYQWpIC+MvH4eLwr
e3F6Ltx6/gS+5iHQP92+VYyAD/JusvEhP63RkqOaLVKU06vPUIQiHY5Amo6lG/Xz
DYxUM17vAqUUoPFjH4b0zWNED74oy+UdUEmRp2zCNgfWmjK2tDgoEYPD/Y+yQQBp
vYJNArxSCgkEmoVeKkVZ8DpE+vXAG5zdpB8HFvxa7+Im2CP62BCOAYyjvBcmglsA
Pfpk8imJz7Nb9AYaKUEsKkYPUyXAr2p8miPL/wxnmoSh/LKUFH8MBFA26LHGtqJy
1v/qDGyvtmk+D54xK1jB0QIQPSUuuZFT4IMzdf+TAoQ9gj9Hlkgvt3v3yMgT0Olz
5ArWxVONUZy21008qTU8gsp06dP1LtGs4x0T4p8M+Vw3rddUYb6xuhnFm2K0ySZo
j6wIa97lV5sPMjmyY8pnyDO5jYwxfs25+67FVtD7G1fGBd8CYZ4eYTJrVl8cjq/H
jKBY6ksZ/OPcJmrcXn/Twnsdm1CJZFYXe3L8szo5ZNyGD9f1cvNZFgjZ/0/hosQL
+dVcYAOx0+HF7otlByF8kAFZuCyo53R6Pibmj2phnfeqFUlG7AL0fCNM+8GkRXZC
1UeOjEzqPXl8nydwh4A1KF2p1fxrEozabHzbTjCsMnyDIZx/iGMOUqmZLmlTxvpY
tDFMIxrIcJYC+t36eW0nHyt4UVFW71DkMBVsaDT7EHYuc0Q/Yki30dbxoskHI1I4
61JtXm0qOPFidal6DT+1Kz3+Cod+44jgtgMKhPmUCFq0rfYEecGU9BAfF8A1DlRn
Dije3H2R7y9ojxcwe3xPvd4z8PCfJ5UIWERvKNklk3FSf4zKmLkpjQaCXY3hMsyV
w09ypbYcx2i2+x05flcqWoT4FcJprVj7WjnmuQ/CFKKoj4fIbeciuI44qghmlm+I
HQ98sNvF2X+wvnfawXTIQDOw6IFKeBzbhOj75zGOnkhCV02hgnQ3LY7Wx1dqgdVW
fx3I0IAaDtoUGyDiEbf+zSEg0pnULXHxfMqb3gRAstvHWhYtovgnVhKmGxVTZV7r
OBuoLI7W0wktU8YNiGkyPtpSnrrF/fPMUni4anCK2+3TIEUWOIqTXsyQg6dyUouk
8n87ym7DzsLXqGCWXCOU6zqr/5z3hScW32iUeOYg4oZGTBDZM5EBMVrqkrXjIU2N
7CP83skEWFE28ZxYiXeKS20hzugqQMKb7f0M5ns3kUh5YU/Nb4b66m5Epn9sl1NQ
NVf64E7m6x9xbUguSAoM2UGYjGUwlkW7SYjqVnkE+6rJBaMEulHe6+y8JWY3QZOp
JsBOwBZWbSoi6hUKqqc1aRk5kfqKNlFK0THoSqKz2NlKI0brYg8U1GzrB5Swvvf7
xjrwmtgFCqLLRov+tdTZJVq9te23qQ+rY2reUJ2ULqcb7XCi0MZcRGXQmaO461J+
l9H8cD6H73uKY8xU5q8a3BWCy6jE/bZk51LvIfWwPPm8WjXEfjfEL3SzgBS5baRy
gFgc3iOz2UrqfiJ2srNECxHHOtoNytdLliMDyxAbjECe4a6cfL8hcFxusIknmy6p
kIhE6ZUJEHcNhYRqY++0NwE2D0JjUjaM8bEfXBfSk/P8gyRcm8mPHawOh0gsbUUI
EbUiYSkeTwScMoEbajydlv+a+pR/sMv1ev2AZHzpvBZ4oJpycBjZXECDQwwUrNgM
jCqMIdWWyM9SWEHFTKg+nVAFmR0FkTXthHXoQo06OSt6gSAE1ewTXYWJ6wTNqbLM
cfBuWlAI/bX7zHL3XL1z2fAvB1V6/X07XJ+VzOwAItj/600tPFHUxEqMNDX+3Gg0
jem7xi+hlX5opa+t6yJCtxZto7k1CgA2OmFKzXcpeMVNBWO9+36yl/NfGq3HzSCs
2pGiX0+HiiOacxUbxhsnxHPGYUCUw50XNjdTpdwlJeJ6N5UpcOg8I3zgVlheCXho
oxIROVKUklEElN6JkNnjXrXnwclfgryCgD7DiGxD/H6CSvSJVc1R2B2hYMnZw2pP
bIr08FAkwGzbkGiINuU0E7+8oWdsOxqr3KwUfmqoc8/FSQiLZ7WXnukWrOjHIXxw
EF3wednx0T7l7JSRXTFO7g10tOeieWZdwq859U7S1xwkYsZlvMht4TAaGClqtOve
4y5X86CIL5EregB26yZJOKUNbqA/XwvxFiadW3K06ILPmdXSHr0Gzt/59q4IJ0sS
w2HYvMPn9SPdo9vVkmv5lU47NgV+kZAri3gjXJSwSQtKy3tAcXGmdlWkKxZyreTr
0bRVSWXxQH1DUGQtAdNFoj3Nwxo/X1D+PNqmHruVF5Gh9y3vgzvVMrCL3UXrMs8h
4ZEDa6XFhp6PCgdlmLMje7fFVaRoa1w5l6bcY9IgFbW3ZUqfoONY1gn483nUTCmh
brM76/6cm2/mCFT9/Ob9Kg8bhCVLaR2LtZOj29+S/xAz3KoiZktVXy8ZKEQIaLGc
aKQSEyWaK1CcI/F6i5g5IuhF+mjbWGzLNJqPGiawpuO9NsRiPV94b0cBuUprjYJg
7d3cJHgmY02hfzOlvkGpBl/O5mtv1ELUzSSK8qMByU6CBfH99LyHOhTK0aBfPXDi
FYYKM5cGSAPSGcs7Gqrs7EUHlEgVY7QN+4hH3qIYtcaswkssh1C5mAxmV8bWLyME
VqJK34ufHjJ+9X919MH2VvyPn20Y4gtNhD0Byvomlof3Yu7TS+K57TtOeWGexbnu
pAdjpBWw92oIeOl5oa5yzCZYS9Vjg1VMd3dfMwcJuhdd44Wrc/0BLR7fL2kNjx2b
rGHM5rH0/h5gAO0MxiIzPIHCig81TnKd+DYEFvRNEewVe2UmbIadw0Na0eBOJ8NG
/IcGKLIlKuFIzpLKCv1aQODf3RNiYgcvzmbRrn35+UiZsDo4GutBtGzOfeN4J0RB
8dbg1qag/nU5jKiL7w4r4WposdLbidOdU66UQXlnJwwz+vMJB27vIzQlurGub0nK
FMRJOVy6TESQNqnYeIJapYOyHwSypdXIZSuYhpVEYvt3qz8joP5LbJMjeWxQGnUo
VbuaMnezNkQK7YWrbuL9PPFxYvme5oMlM9q5rX1LsRi0SrPD530g4tMUeR3ChlLB
yLWoM2Q/ewzkKOB3OztkvQs4p4b29wsWwRhjRZ8S0BRIeinXC9xv+nDmmLQ104Fk
ZDE7VrE8pREAEHPMTeYL8arwwn5GPPu70yPKGIXozA5mSXMm4D8mMIDAtKnhj8Tv
VNtakRlrIYKLIg/CX+yU3sdKU5sl2b+8b6rqvAF6BiCZPhsy49TyvRLSLXR38xEm
Ng7iRw+PI0UgjrtF5Zf7s4ZWGLsBQGBiJ+SbCXr0mrXIAlx4d6TBoWQZ2NzAjERL
Xxepi07JUBxXH3aTxTdHgGWaP0TBj6loMAaCkTU/VHEw3zB8QR3CP47pvQ8sCZfo
AgbqsQqHteMX8Qhu94lC2k6dqv3146pEwUYU8YM6L80GXkHFJ0yMJvpO+3MmQhSd
myYGdn3PfxKriyhaHLMvhe+Bxcff5gotLDn2wWQf4+gWfAEPVhcr19yLzGaoiCts
rvEfJxze+P+szxHH+9CFVJaECJHF5cMth7jQtKpLrw+Xcd0nqYuRCdiykJKn6D5J
AvP+GKRc5eavSS6lFsQXeOznRTZH5zA5KdUfHeal1KpV3r7j70ly3JjDj5minQJY
ZVfK+pvB4VNTyJfT68WFeWUC/Huvw2eoyI/TZw+2gT5o6JaeXxhECieeAP00qGY2
HVqS9r0EC/ezU87r+kF2+hmYCD98ajzi3kaD9osbxUBaUTvP2gxQU6XGCBuUcXTM
3Rnwr7xN+Btzci/XYGNa4jgfgq1/uowJwVoCT599fT6M3J/lIkZf1xaZV6Y1jtC6
9YJNWRna0sOejtJJ+R133JuyE6njFhhPPPW86ocqbksxrSbXBnDIgXA1+c9WbaY1
ECrtBv/8THk8EAthR1f9m7CwrY31K3KUEt1iNAyQDAexomB2NQ8ArDEfCPMDLQi+
XJKWojBZTA5P30n2qx2kV4Ct4K8uzCzrwbIokgJ0/3sFzPwS7Vxj+fjjkZYsg0Vk
4AgMAhp7K+Q2iSECflUrplNwQUN4OaU1jcPorcE4XDWh/Vtm/+Nh7lXhcRsyep1n
5mSMvxt9kysgE1nqB+M/9+T633xpptmpYfo7Xn1oR/a8EBgls1EG/SBdySJuCL5G
YG+TfsBdfMY0gRAwWJtR4hw4WFKbDhIQrpEJ4DX2vxTC3m1NbFWhrFejtGWa8G8b
AjvhegqVmBPp0AupKen0Ss5qvxH35jAfC8YQEXRods41qPdQj9tQ30yUn0xLJCHF
eANGKoQ5YR4+9xemo8ph9bxtZ3ZVcHVRV1l8Q2uInQWPkwNmFkcAzcsAyeFUZjmM
/1z4JWLk8yNjuygsO5GOGtBr47HozXE63Ut3ATZfU/CJYxXWa5BTYT8jPyBF5Inc
bID0DZEvZ69z1VQuuXlGsREIxpSrvvAL60hEzBJrZaFZs0VCktL7XDPV1784VHnw
u8ufjnaHGGTLuLPB4TunPRPcWpkejE45FW+wkhwslNgw1YV0K+Fxy+MMAa4PeMZ6
5eWHu9tYNMrQp/1s/zOiUSWpKvJaVWzVK7mpsTIM/Lmo0hlmLY7Yv3IjwiLZGh+9
fj4XuS5NaULqYjtd+mDCxuErZGukGUHq6xuQylSlt+VNMC7sVCTd06FhoYGSj6un
wz03458W6bKmuY0kwwpUZUp4br2/Hpqw6s3fhk1NlVKi49+iu05v3LsHr/5Z12Et
oEj9GeyJ4aPYXRSM5MtYd1/DiV2lQlRE+0Wv008fn9Xw7i75yHxsu8kvmwVUxfE6
EoEGuUv+XCnh4ZjTSt1wzROL6ji+lMttz7xG0CpsbaNtqSx+Xo9nAPXYyiTKhp5+
Gd7zenCQ7ScCBq6U3e3RihGuRQALMhMX2lOrrZTFYUuIxZ03/FM6byExsnMRt4YT
WlI9hjMNo6f7xDQtiiiKKobOZlnARHiQSU7tRXdTdnI1f2nbE/0RRuf+6yiv4HDq
KGuDkfYp9wi4Z0vqTB3yigE7ggc0QZ3cP+YYbQxZkhw5/9nCsvfZ+6oPkS3z5+cx
Dkl3dqbJzN0KMqBEFeSUVSZSA74AIqoB6Xc2xU9L/e4OeIHR9skbdZQr/jghXjba
amLTmNVMm+gYy5LsV5+3YV0vFGmgYxcVjFtNRLCK4HtqhhuxNNWyucwUcP0WGs6T
cjjEtbF7g0qFQa6h5sJ6eRwBGBRwYJBAqF14SEBkMGMfgjZDu02YbBJew+5bo2tm
+h0Xb4xWGejnKHLZMC1p5ExdkR4b83m08uuj9RewQo0akpsrzznV8UWzzjtjxsoO
AioYbWCNhLVCMlludOURR/fKSthyL67EE4WckaX1XqZ1oIDqgqj5yR3DXoB5T2MB
24MLI8nkbR1RSLfWna0w0dB+MegrOsnrDYu0Hweie/Gb0Mz1iM2mM8obQBwKUiMv
F6Dkt3P7H+QJ75IhOLD8HxRqobhWTB8WA1G0iV5p2ujaL9Ezj6Mj7y9+8tWRZycS
+BsW+hApQG5rO12gCeDRDxX592kT5AuC6r5x9rA0k0uuyYEfprxW8sNcCVLPN/Ji
j5z6RYwX2ia429oMPuc1kZ8G4b9T4id9qmgwBdKURtg2622BfxuoCYcHL5POyz0m
Valgj34TcKrnpmxyKtWjwyYzw54MhrNl1ipieqk25fvzUIdJobSLiUu+2A/EET7C
aSHqbBR0QIoS+ZL2fhPQUCejQW4FDu+0XTnWmfiTaUpGJjYX9zLuFpwa1qZpOGS/
7VoCFzNRXqzKzCyYBB1iLDe7tilKu8DRBkeXo3K/1IR23mAkqRqcjFoDA9I8G3Tl
ic7QrbRFvBTvHpb+cdirvuUb1uyTEW6qn3zxkVtMTDkIFKUaY16u0N6uG9walDgY
HLjmYsH8gBtktNQOzoEhmNaiOqSz7D+apCfIRiQkZtqUL4C9kx/6ofCG3Iy2lkck
pxOo0ZYtD5thkyltMttyPS31ryAO+OECNjaZAaL4JqCoMfjNsCOAVJ3RM2YWaqAC
jznDLLeHye+0c7EAwzFweRX6Sa3HgdeuAsEyOwrwowh2y0FILUFd48x5QHqWjd1E
AA068ui9jQYIPhctHB7v6jv6Kg6jmCDtjZIUho+oKyFAndh2DzELC11G1SorNtVs
YzZXRly0kvWoOEbehNXd0NJEvXQ8+DsInIGy5hKJwB9Yr2cbrybYpU+YGKmCvBzZ
F7mVSDzUy7dvo/mnrgNRBDst9LK3oZiLL7JA2iZAj0ce43sEYnMPPflQGMLdeI1L
sXWXHZn+lN05zjtcPxbpP6YqA3bjv6sPq7vyGJ1McBTbIFkah8AOQWzU9vGBxdRy
o4e+Tw6laZoyqT58IezBc+2g1ERUGTFLTwf1fCUur3TDBJ+BKqxIp79w2OmCEAt6
KLBZSZwJD2XZswbslyE/JX28WVjj0GpMifKIbyACKNehXP6rAzZFoM75VxjNNKF7
ZpCJdCD5FXrGXvfExJ99bis+g4goU9c9PKwoNO7P1jYG/ZENjvplwUesuGeiYLl2
XYKt2a1APPkBkVpfzL6hhqV1dHvnNRXcHZmA9AWpYwPnMxtTc7r1A5a4fAoApln9
CEXVywAKQbrpKltfpH3gSSWlqppkID+7KGJVI4NNGIFfEmnrBdk2Ut6e9rIBhKpk
0NP9Iz/qa37pidVuS8XfaBlbfhSo8uqsOWkSPpiJsrJXXtap+SN4WUtbMnl9MucT
NNAIzc5UZCRjZ/SS2cPRrfeELYKIb9Fu1ERa4U3ebuJQBQdIvu3zH7EMg00G7fHZ
ErKLUqsPRsds8NE09iCAoFPYrS79KhECxcbEBFqGmF8/qYEpFTpft5GbJsXi48DD
uzEqDotnLMCFmu4cONKbF/wKLon/Lb+HU0Fy2KTp+4nJ5qklaCEY9Leb1XkjEkNi
uWowgEtecl/9jWb3yzBcpjM/5cODynJL0hZ09v5fQGiB/vRQOaKTZPWK4D424f85
jz8O6/UYrncrauNOlrE2ziDElmZumuamYK7PSQrx3PQJiajaEhZ1Yyaxdyjrfp0X
VaWpTfhxjn+6xi0YtoP+FWBGClIVvs5ZcHCqBlQ0JReJOFRIVJcCwxlsHyZrzTlq
TK/dEHbPyA/ZQ/91vBarNpRP2YXx6S0IuEGAA+53uYcbeo1Q9WzLq+OHoux7MpA7
UMW00D+RItQBxLoROESy+Uu1YLBceqUxbqT7g/fkWPZqRqa2gJPrl6LQkfsPTM3T
xBF5v99NhbYv8vVf/Jd7Gs/8RxAfdlhg5ktUrHVp7mCc0jyrUsuaGTZlCmLBttTI
JXXY3Twg3eSSDsNABe+Uw14Jh1bSYMlia/dA932jxN64You4nhdmXZQNvAPWBXYC
PwvbqVfNAiUgvuouKCttInHHvnmS/xRrpxKJuhP+Vewu4M8o8CO+jfwxvrl6JPVi
UkUxKtTWMzICvAAlVqsJIWuE1pMwWioWEYbOt1WeDfgl+nCFGofsx7vwNpGRolFi
tpXutSahYAdNWCw1D6hXzxt7t7zr5WFGkK8Ci1xT0m6X0rS+6nmEVNhP19sC/fZv
A83pbaUkCihavQ+B6/UKu3Yr4GNKFjMTFh32Gu/rKmgvaCL+8LdaZ0S+Tq9m0oux
WzuF/cl94n6MewLYigamALn/FM9ai/EeuX9WH5RCcsBNJ2DeGcq4DcSB/P45lFIq
1lEP6X33X7nC+0WWyICe+u6CHZxwvzWQnnjoY09ZLPP6+tMFuBhl+EqLleRkP2IU
Ub5ChU6SJLG2ANXk9Bv2vUrOlVJynBwU6Wg5XbboBb5D21AvpBayYxdnJtSfwEx9
KpE12eSbx+k+Vws2BimqUgpzu0GA8+JfZKYnk/aZfO53CA9S0E/5jeIIFyyksVUx
Islo+i6qMloPDUbmTQyJab6RC3BdF6kjIXhGdP8TmlKBNfh+1brC6ckE6yVQwU5w
Z63hg/Qdu3j3b7o61LvSECZYDhAitW5RmEVv3yBsWmkR45ZSAtZWkn5pvqbjKydl
CrJyEw9y4VlAmJ7R/KW4WIM3Ysb9hyc655lvZlDyPelnGAe/+4lCLv/GZXNcEghl
ulrXwGw+FrRDyWG6X8GN8OcGwaz0zKsqRvC/ZVRrFVo6WBscj/Zz4imueRNYvyeO
NZ/Jl5P8qxj+YEOkF3I7VLZvW3cZNv2Jz5Ck/uEBKuPe0pnaKLGOmxQnN4IkOulJ
Eq58IDzA+gRmoR2uDYgi4OM/e6Ieu48SNYUW3LMmFoJDOjs6mn9F8Fla2x2zzWRz
cAn9qUOcyGl/pMYPAs7Q5TL5CHwEKfpLWMaFgI9nMQydUBJ0m1k1Ow07VOHQ+yOw
DGsIdhtZ/rZUw28LpcG0v8bo//Wk/9uI8GEpgE772yGjDCRCz38N8KXTgkDQmQKS
UdhFvyf5A4HDlzFTn14+tTPtP4VZPcEnD3lTTQId7Q22UU0k1yJw7FAyVXCTkAFV
A2kuCPtIQIb9lL7p09XFTfLVnGhKK63RPmH+JZEn/6dxmoqpyz9ip00JBRe6s29K
ZOQr45nmMT6Wj6fw1KV5pmBt/1GJKdQTAY+GMJrg2cG30iqDBtFTB96X6YcIvyLp
/TYItZ5TMOJvna8sYTocWmjPLf/IaY3YQunCmCgzR/1zCGVcAsrU1W2HHZ8lNxll
Mi5Q2NAL5oS+1MtyG0yXlYH+DL7lLsYB6+CfFA7EAvJ/CLk57qAQSQmBgoC2WbKD
M679d4VQbJVRuv8R8qsAVf0N2MCzI5y+OoRwwCE8WkzyxziICVhyX031ry2LgTwG
/JOQugrXYms6ByDoep8h48UAbB/VRZ2U650B//oQ9zoezFylq2fgJMd1/QZ4fbzB
AaVZREtFC6dBFiqqbq2bQ8AK3+RdFuwaFOlgvWDVgaGJtPoMkEfsWjIdNL/uu9R8
3cK8h2Obw0O/OB51ATdi+jiUISeSbgw7YJmMZKnQRHRJIlUsz8dh0nwwWclu19Q2
v3r8L36kiiRFxXD/jNdSlACVxiEwmoeEKvcLJJRCKiKNQGo6U5MVRa4TjCCecycq
eT6j59cws+4aDmo0R3sgiBGKlnRgKKj093bBjLZlkdOStMx2o+DmxFAwFJEJMQAS
lGnqhLd9IJ/a+Oeb51Ez2FXt2n8T0lGywX/9SnnTYKKro8UkB9p416pjqx0ZU8gB
w9CBekVDAUSnKOHntAOtLfHQ9d3WGOTQxHjYj/KrAlff4C34yqRG+CYmnVylnu/V
gTp1Z5FSI2NAEzR7afMK6vnue+5oEZHofdmF+y7LIO55Y38/7ZmkPZFd8kFfmAP+
QupV37sCqtZtZx9JcFtIG/OdM0hsaSumSZ5gh1kIN/ve/YFPIuCsM37UX+mVOgMW
qqEYi/wfimX8QWrBwV54m32NCWyQbjYUa+eyxjN5QrNxUFmADDKbcIzawmrI9iO5
XmTsV4nEc/v11YRqnDeWdnZQ/w2SDV3xYfkPv3QVg3sHFQDdbypjBfZYymsJOv1q
zcVxNnPWcsxw6EWPcrDwSXF8ZawzoE8lTHDf0DYitq7bvCHdgIwUQ3MJtAb+r/3f
l6Py2P1bU9Hgu6PVEfoIny8vdTQqHSBqR5nXDt6lCoN6oOUiDZHWVYpvpSdXUiye
gpR4VddAof435XAgjcFGSwpOXkKKpIP8OP/F6+9Rwxn/HYTl2M+P6ckiqhSFWJY/
qwvHmdOZlLh1b0A4HrXjySL4XVsXSaSvdseggohHQtQmIeGasB8J6kEcMPfLQSMd
G+Ki0ZNT2gVCrjBCB1m3L9zPdffxEoklmXDcwwvi5Dld60nZ0s72HEX+bQ39fGbw
dE1PncvYDvAXW2/ImpfxtmG6JYSjj9Bar8SWAJcQIXw2GhMjBLy2pjNWoJUN9mj2
wxBggKRgFSm0VRLI2afT4BikgIpLIZdeVrMQ44yLKZ3MUAqs249NhHQzFt586mqU
a0RQZmbRd+jsNLPzT6UdplFqT39wC4BliSgWu61HDWa0zSYSQDClE4rYRVAlqE9e
Eimifa+X9Y9zlHuOb3H+5nBa/4RL+YGtaWtWVTO63xL6uyUQ3+AuqOzB9tMInxya
lii2T+U3ESgJ8SPte4fmbS60na1RUMhL7jtna36mf6VorJeVHKJwx/mmTKtxC/So
khEyN8Z6dtKuHOAzD/1zLIE5r9OolqMlJ+5m2QoaKERbY+b0CdFhEOMgtOwmOi/t
lmeNE2JVIbnjugEWPNxdMzIeIWlfMduPkdfLvmOMynWol3hXZ6wPnYXsjKH3Cgt0
Gx7ElusbbEPebIkZKP2NsdrTcD8PKlrU6+3t856mDBsfCBl+PIz4rhtPbviyZwwQ
Rttsp9HNHX9q1wdE6bP2NjFkTCUc8MWTy+KoKzjAi5GhLzYREKmhr/OlUsyo4TrI
jK8AG0Bl/4wAq5C/gVj3vgX5lW4IgqxEUni2GYcAlLPZ3cynauepGI6Ol0nMaTwa
u+waQYmimW2DgkP6RQcsy8u+5Qe1o5sDD6huWAYbDSW+6sBS5Jmaqgq59y1naGKo
pI6gaEiJ4gBIcjqDhjtOBBCDYYkI11pBUXb5QpCNPSjfkppXrxvzZ/9LphtRT1V+
fvBrQ+Xf10B1z7BFhGi3Rf44GMtKUiGNWwJgxqtqAmH91IoGCdCKAiwP3SmPODYU
h5hqmQV2z3hbfX4al37eEWK4GVal4RaF6fL88354pzdCjCBRgTRArsmsrIjJhyMR
ViYYJfWVOyYM+++g3b7ZI3zk2iHy81OV4RS6z3Cr9tOmbQGkYhmbVQS/LmNqSdOZ
zucqBBQSoHPtjE61AhaFW5oytVWYMuPDy0BgU8rpeIkYLRtS/vnOJf9L1cRTDjGh
xqKQK56q1p/iQQHdOyt1Z+u8X08uwIlNnyG3/ZLM66C5KDcu6F48TWKQYhKVoZz4
f4VvIlrHM10wbgVsDj7eACLW4DORlsalj1ZZOcNMy3TSu7VxnqJ0Jp1z20GcGfFG
kWFzQzDlFJtANKci5jmcm6LZUEKd2tDl6asd14buFWVShL783znem8u9iHv7EJl2
ahZWDIYGtYfeJ6VkKw4PBxdisF4L/dumcXCD4c9gV+hxKASrdYK9Au1ed++QNvV0
rfqn1ZrtnGMo8UYCkrBnGco4rBJpxxnIQBIEknPVmYOrwskG6j7j5TPbAVIPRhqc
IOKbH03f2SFXg0mEj0Wh/o+Re4l1LoclyUNgHeTDm7wuMf7Wvnoy/xARbM3Rwt7k
dfSMmM6W48iSUwUOOALGiwsRI800AYPvnymhl8/v8JxrzDMoNM2stktRHB9LXWev
Wlj3QtWqEGoaczuTDPZBMtGfd/+/A5kImx2d6Aw4SeKhAlcdCtAYfKndb6G7r3TV
GbPewzJEqlSEDnCwK9bmdRyVDBLG8fV/43azkE+Sh/R59HCGrV1Id/Zo7gjrTz5q
HKs5Muct3dRkfRF6aUtaiYLeu4uXkRObKzR+sj4rvaQgWm8rndlzFL0ryKTwIMbh
XFDaEHa8nt0Iw5CwLcDaH/GpvbSxr+8Q7sOSRD9G8OvO6wN6Vie3RcJnCyYk6wQZ
nXeyMK1PxBaRIMjyJA8P0HYv2rsRFJHTlBAq06RX7WOQTjXODL1PSwbWcNEWvdNR
uLKGw2ZC5BZskvDLsvKiMf5ln7mNm612Pw/IttrG4fJfFK1x7e+HqJKjzG8b2M8j
fb9TS/ne5d7b2/s3lS/DFHJS7rrQ8SXLXvYmx5Su+yHvO8wII9tR81crO80LbJB0
f0vBync0q4T+rEnS1yz1GbRJnqZhNbiIV3zM3pTn2Hl4LSI/2pAsG8J3emZFx8s1
hVNxBREyCwhNVt8JechC4+G6/xdxvhSRFfEjtH2bgMmKnOBU4WMfHVLkIEI3c3ow
DJy0EMa7M+qQJ2ocsZnpLvKumDgUL0trRfOas1RLf11Ix1mtAziooBwaM7B8q8f1
db82CmiZRrEGKbwgUwHFuNBtJVXzWB5UMHdXhQnpSkmtaj+wKGi334bTjs5meT9p
TlgIs3FtyX4duoTKnVdzyAQgZaYLsjHWdus+kyZpjnLmJkQ8ujDCjiHFwU94MIwJ
DfZfWcJ6pst6z8UgMhFyfAVzZBaM/dhRSEa65XkLrPUJQQD6RS3RxrsMCkqiI7cf
MA12DhtTrY14LtqhKbnTZQBB0NU0C6fFCJEQBZ2FgdNlHwBfl+ajsXQihllvoauL
AnwHjNONLGYAuzmxvNfBeYwmSlIDjyP8oNBguBOIP2uWzAAN2MKVAzmgGaVOwZjT
8gaS50WQj3pqwfv+9IqgMLSoZ/qJlelzu9x+s6MEvRxYy0e3AlGtTi8Ywl0uU3lT
BVDMLQOnnWnj34SK8B/HnAPrF3WGDWm/nCeaK/AZAPqhAQtGqe5jVxJy5Z2SywEl
JWbBFm5xVcLi4RZ4H2ds04uWFrRS5grRdlas9rNK3OfAbMOpvurneMO1QKsd/BcY
Lpv72r30ZrpZaJbXt9h1/ZZdQTp1/vt2a9+G5Jh+EhPa4nZ6R4g75EEUUnvwOYM8
6Eog3vW23PZ1taj72QIBX7Oo06ZRO2dL+BFm4kjXk4Xsgl/vVH1xROuVa0HBHS9V
xGN3ke//gHuHuVuTXEWiQ99vq+NaLd3oGiSsPI8LnZ4zDS3wd958UlhUekRLIS2R
sk53sBEST/ZQyPdtuSC4z5Egu0vsy4mw9na6GJusyTSN793WuQu1FWSVdPImGtlD
0v4PhCISHZ4YqICSPr0RZCRc/NkrIWDeXLuDIZe6Q1gNBg5wOfkVgsVV1d6uMlqK
6ETyapbVxXk1tjGY7a4RQhzcjyKI+JqqheWec8XAXoToq6GEimGbCGyt9/MsLU5E
gjo0/V8KHHBHX9BRrHnfdvW2Z6KQgvlnQY6wbwWiTtMq2wQg92NHWg1cnD/of0xi
K9OVur3CzTCzvVgOvL9Z0LBAY5CQ/l+5gdL8t5dh93IRx7SZRETBCg6jCHewNoSA
K3vnfVMyKsl5TRmTXEVRiyWaUR2R+S/MY1wMurwb/wOnTn1JnFFAF6NmjJf37BCv
mIu+c5wNlEH54tunYijpXPH/E6rCdNVZy5JzbYXGj5WRRiuiRvs0aA76V7emwqz3
QgMBb6XJ85SjpF4LY3gc/XBdu0GChh5rHenXd/tFtoMVk3dBB0Qtq4riis/yYQFr
Srnvj5+dFAFk8Xxuq8u3kyFHCaQNnKHGu83kDmYDJOm/Ci2p8BocrlR3pINvhmka
xZOj+4kyo6SPpZrX75Td5hlvamfsDyTt8/u0aOSMTmZjgZjyg5Ly8Et36nwxM7eP
GLSVGBQOtMnyw8tvrSY4jfWwx1Aoc5fmFshj6X+8jhZ21cqD5qYz+nQuZi0ltxv3
oWpEIiDB3w2jnEeQ6krb7jYTyUv4tqitrU3wMmEYSgWJrhP2Rmt9QuMwwPko7nTF
5LlMAnFztHWQdiGOerCcRsxuRJDR66eW0v6WzdtxYPTn1maG5HziWsuqqCtHeyTE
W/mNnhdSqIIXtqHvRP883exwVGpO+PC7o5u7L4F8pfybIyp4f73PLN1obxnnCdIC
ZUOnooj7aDEUF+uYfDWLas22WGvN2/TXf+inHOTL2i2vs/korRD1HPZFuu1LbvZO
wze5glI1OTUNaWInDup6GBAAKcNdz5gboTnF0ae/H0e+dKs/5DbgRqpdpjYtD3y2
niUEvX/sJuw0PqVfDiUCCcrVFZBXmzsEMewOLyg7fXSpito3kvE88vC/19KqMt1q
6dN7lCJR3n04v0HDx/KCXW0T6Qiyqgar8k1dNexHG4KHMKrtFuif7kWVKPwW5GLy
k7dDjWKEUCJsL6GtN2k+tXpxvlXzkBwmd24c+1WYNCY9f08QZf+sBIjNDxGrWEzl
lTxw28mGY9LYAH6DQNRjYiiLy5bOKq/irlaNqT2pgcdCfpyGKfs7/gswuLTcvCbw
9/h8l57N55uUz3WEa+/Jr2LDyzJEFSDEtjnCJcPz4TTbaMFqgsvya1HRdPdc07XU
61nvrYgyUfSMcrchcLxLgdVIlWFz09y/WRhmjCF1ZaI9TNJCJSHkGEV6qqLaB2FZ
V+WxRgk5wsbG/eYE9Cn4qJF3d/Sbu3TDA8tXwCbeR68EVxk4FTwxv/xLYMxcYmld
1ssgUE7GUUX1WAIE4bQ1ZqJ9JAZMKtGg9AnzGCIHhNA9i42cUZ1fHc9mQswqvaKC
sU5h3GHICLffyLDDtzNhO7ObZhHKcxUwJetAWAU9yooWEayKUB0X5zzkzNoYy7Fz
VI7veTuNf8+5bRagicrxUwcrCufABJz+NflfOe6Q1VC70j6twesGUTdbBAZxjG90
v0ze0VOvDSfTIBmNGSTrM5ssMLMRrozbMWhGisiaun1AwZS2lyPr0nAALG5yud2/
N8AbkOEbafdWNHsxOSDAwS7IX1bW9bQSVOuwuwmT4vjfR0FqPtViHW3uCOhvvC1v
8O6AVBZwUxzll+xpmyl6CbZAgNIztSDSQHXZUB3P0FsoQ2CUvQvigfRkskMRTRN+
rySMnNJ/ddefWaGaAbTc4VxibEgMDIKWM4bSmgmquszp3pRk5zGVY8CM5W2sEeqn
2jVj/9yEyFFYHX9Rl58HHqCBCKKmTZplfDm3XWRYgAE09S5yxy3JLuQtBuYzXDGZ
DHQ0ZKKr5+OAWcTq4ZantCxcr4bwSDNDoUxbxpm3mhmrg/tHfgG5mNrvJtcgdxxv
YnnPZNPnT1yTW/sSLq9yJQrD6bukrfL+8YEJvgWndgHkvBtXxfelXx6mMIC7C652
4ec0K9XID+T/jhlQcVjV8BOi3ISVhvO1Z9lCPeOZP+knAsa3u7GojpHU6ROKkuk5
WmS84vXWU6+YpuO1e6dvYGv8+8GUnJDW6EOSYF6NcRPW1Mlxah+wi7cvL1641j22
Rnd4WIRWbwdp+OYt5CRqdwbg3k8MSbE/qWzludsKLi4fDcC2X4wshPn1jrSSTuNb
982FC0z9qDm1ObCccsF/3fzxXAdEAps/6C5qJrf9awcZnAX2FMJq0d+EKT0HTeWm
7rXcvMH9iBTOKFkfsKf02a+489H3qm+E0YAQN/8IjinTtafMF6kg1kwvLaFAdgYO
vQJuu3hwIlt3tlBl6I9glsWtxpvC6jYf+6ADFcykFV3XUvW9E4crKSmTdz7+d8aO
7+/DRzRwF7HSX8IH5WdKSeySqjjgoni901PlLUB7JqiaO86Sbdb4tf65ZS1gttxd
y6jegcgVqdyEVFvEp6JFInxiWCn1KTyk/WbQUHJ1Biz+Wu7kCHprPzYHsPTqlV3T
g9zK1TjVXA8Dt2cGbzW63TPN37XW7G8NnDmoqP1leDf2Moy6a/pJVu2s1F9KVzX8
jC8N1yPCJtc+t8dJZ0OvcchlbUwwbgWdjz6ETS+whTlv/L8wqpedMU4beNtwI4Fy
0ZyY0AXoj105fs2H8HDYV/xbUJ3JladEs1/+aQMHfgEpIlR5dVfNNw0QJjRsIJn4
qIezMaU36wBOxVOGaKTReaKcIVKwcbqNqC6ItZxUE5OqVWa7izMPC1vjalpIrgLi
Is75YHWrspZ7BwmI/iZ2cRUCq3lE9FOzHIAkdAe33oZ63mVuVAhNpuPkGXwDzJeg
/GzXgfEN/xg8gcKcEnzCSCSI8Yudk6YFMmQbdRB1oc6BJFiB11HI4xFLlcp7a6lx
FjXN1YJXhu4dMOTiN/BT3ZySprUdOMSHmYAyzoBtkyAJXoDKvcpUN4jyNYN+Iy9Q
TQx6Kqa8CqPaczCMcuJJFkQUWFdTza9en54dAXtmul3npbwGUW/U7JD3PEJpAtbN
OpEIEdSdP2ZcOXPpH0/tCtHmdoIjmRXcFlXDvKh8tbO84FhsFvhbB+Sy+uFi9zpG
JJsSja6cDiRaswkH7XHG20hHoawQAlQsDR2Ps8jpl/1YCrXoMQu59ZyckCdngE7n
qbbZGeuzGPcH844sc27NuQnCPi+/0XP9b76p6CwbUk4EsyHFCVwAyP54m2KmOVw1
GGjDtGD3YRDtzGshFALHnV/HPcfSVhcNWKojV0ZlnMRdl/c3fWeWRkcDwGGUShLN
9BiDe2OfnDSuyNJJJd5+SjGbSNoMp69xG+Jy1EDvls7J9hmlaDE/CD+yx4lEAXLN
CVAQuSI9hLptKycE0/XSrXlEeFAj+iIPbmROGOZowrLukZOw6prksAKBDV/uID5p
REkGD/4QQpZ6rJJhQqztDhUU4lA4zPlX5rIG0mx2tg/r5MXqsdNwqdmP9/ewkmGX
5GDZstT2efTdHreca4oUY45N1A5L4jIdFEINz0nJ9tI7Kle5NxLdrsplLu/PwL41
TLkOu7Vn+TTt5Ylsied2EERjNBRErIRVTzf/fpqU4qHQZBXtEHsiOspaGA77fSqB
jhylM7uyojLKQvlNi9WHSnpO2llr4WSY7wo/dWbF7hOWxbqYyp6o2rxiwtI6rqaJ
Drnin1b7OEmr+x0dr4YMuryaW/FlkaIw+TlGyn4u9LlMe6xS+2tEcobKN/ZjbKYy
A7ODZXMSV1ERZ4iGZ+tzcPyp9j5r67ovOMWg9bwKju1UxqEiVGgg672V5rJ339dp
ucxqwNEI5kMaZedvpP6jhI6WQ9j68Su5+eCW3R1/4N8lEUukuDTYzQxK2oYsEHRf
OP1xvUN42/NC6gtXeYH4SIbHjBpJaUT75tI+ZP5FZ90IXbe/SkIwutlXtYoH5HAl
eHLpuSns92P82Nd5VYIYeOqzZarIAjmTpymdN9IVz9Tjdb3MGVamIdtE/6WwHNTP
ruAAwzWTkelxCvwswhKGYUVWbToAxfHoVIGIyjL+8Xvnt/kAWkvLspSfwATwBBI/
5VD9/XGkB80zspWtR7klhFb+I0laLGs6yZGNc3Lbl+rIPkzf+77Ksozj8NBgxPSK
R4TXiEJTcEghXYKhRmQqex2IL3uL5nQKSbCOhYL9PyHer25mykLR8dYMP/NLeOk4
TP3omAvC3S9xHyvwlerOU+NOCEEMxoVeEVI98VzMptfEP+bndnEGcQPFi89xrfCG
1dVf8Xbh5OAMlQ/+rBl9Z2+OnEXxwO2N+j0YQwHyK8uJeDG4m/2EDdg7aPBL9IbN
BDxd8+IF9bgSywMIvMw0f6XHuOKzIuMGSX0KzAnGBtpMAlsIJUrHQeac12q4uA18
LaMxdqkWJN5zOKnvkejHA9jHnlQAbCyGRnQYP9nZFqyoFOVwQl8+01x0I7BEJmzE
bOmBXBXa+Kv5pNy3tminkHGhUfJ7aZxxc2JCtkMtHdznKwFRblqABMFSz4gqd3HK
cGCUbCGZgzEDVXNMoZ5jAez30Y2jdWWEZeC0CoqiXTnAmXNwp1Rp+TtTgtNyg+hk
F8Li8bEynl0JDbBRvCyyyyKYV0lRbakuhjP3xrbYYotW8m69fbbn+B5bC5ktcj0p
mcPB0oD/1v4YkbXUPKXtveaxwyBwbvtaxNCOPTGWmcB5fT/DfobyFIvdkAVq/e4S
E1NMOflvFgWd9vJGk3pAhX5eZbnlA1EVVd0S78miTN/xZ/djzMXtCFu3BhCpMnh/
FklUktN5D5KDDzzcZSnnkfuDa5kXqO/0d7tZoV/0uGaA2Ll7CBfy6zTEr9EqhdNo
ZZMWTOVoCDmDoD64pCbu+JRGO7AOA+vyf7yu57TAPSGqb5lAXyHQcO7snr3EGmVM
hOo6u0frMVIH0Epqq1I023Zz/eKymNFvfU+qKk9U5iuQaz4liM2x/Q5/4qV/DdRf
4MwGlhfWN1vXAnex3aSWnAQj98cDcVh+gFXZnKlTjk1VrILSBa+kdOg0OFcXv7ji
fB+ft3WrUaaFjVL4Nd0OGemgM3TFRg0+lOptxFrCfmf/+za2lX1BtFqoqvuX4LHh
JQRSVsKN3DApTp1PJP1YMN+z2B5fkS/1PguqygRQBTyri8hDa7pU785MctsrDKB2
7hZksd+MLwEIxVjMpWbHd5WES7CPqUBXJsYCjhXYMUjrSQZNLoJH9B3v/2SQtroI
RfPz4iJZjsC2j2HVRf9okbAsqSQQnqxwf0b4XCIeGvv9G0e29fZbcIRT3TlEKCE0
jjThor3FEDCo6QEl3tb5Df67+iuriQ4gbuGeY+VsYFglceZZElkeaOAZq4kPXDrf
49olpwye8XCkKtGLcM2I0eHU4TdbFm9tnpCXjHFmBmooI9W/V8bRUVaLcB/XH5Sk
jSaI5ZWs8efxa4dolIruf0hrG5SAGpRJ0oHMJZIy6O2BXcPfFNt/OQkGYnwgPCvj
ezJhCsi0tjJ4ximkgi+B+AOImlyO5x306nWp9QNJnQHRacB0dcKtEwSfBTfoBJut
OTGKGpY7FxG/WisXv0mcBMoF7A40YAkZwAnspIT1DTiUE9G+VC42xRqQz2a1NheH
2rjHwGEFGsjPKMs/BHPRWnF5XbU6u2jXunUhVr3A9kTmr7e4YAsXOiX1J6IB+55L
eP+Azn+McazwXI8RAWYCAx4uS+Ye9aMqghc+z09euAXywFIamXYmT2XbcfA6tC9n
jjiUB0b9fICH9dDQ6NaQalqKRJ+w/U6qOqnVXKSu6zNkA4dzTtLab4fwBedjQYhR
B6HBzJdKQjQxx+5tlieOGR14lvhhOiJGblolS2ow8hSBupXZ7KbUK/1nW+R8xMaV
pFxM4Fac5Lx8uSkNU5rpTtFaOGQicKG3MDvgYyIGTG+oVfkl0Tb/LujPZQq3sDRZ
B2s0eDriHzTVwMQ2un0AmfiSpaP3FGQH93ZAJUMFvIpXMvojG7+bL33eV8OQXoxs
pn1UddJcCnoeWuPdJf0CspxSjzmaAHYBFdk3Fgo6htIcKhk+MRXJxi+DKbwwqubX
1i0xS32i17GfX3yoKY/zupCtpt727nYXYsjwc1aO0eQuLvlj/1Axsib/TvLOtiHJ
d+mi70a6kQQtZUqYZMbsl9Tn0Vq2hV+w8Qo0h+MxqJ3hKUlrzrd8ZngzEx3OhqwB
3NpGXBVQIwdAX9Oq3MPqRRVJtAZ3yMjdtTJhoC6/rS/8MUgghAL+cTPNIWu3oHHK
daNNn03yx+kt+E0xJNh0TfIfrRessxdE3sk0CfSXtj0iNMYUKRZ1sKY/Fz5A90nR
pxww0eDNbpg4xSOdXpEOB1xobzM2hNdUMC2konf8qWl6gOcM5uJIxKeJTkOJ2Njt
qYN++rSIqUQ3kWcrvPT+ykXdsOB8JbceNI5lCfmx66U27iQHecTw7Mz0bRGZ8p6r
NP4LTnFwXwb3D/VlCWb9VNBncDAsMk8AUx9T32H4JeGIgJw43BJ/2I3JNAAN0B0u
6+t7WMM0J6pSm5PkcPrwU1WvGQz/Qoi7qgUMcDHYPWopT9p9uTynRGC/p1RQyrJc
tGbsjVzCQRQuwt0WLl8n5g1TSaw0a/H9BWkmq4va4qwd99Nt1Zf855CYsg/H1Kee
iE+i1js5iyO2tT7KbbY8VaqnOSePonZxnki4duMr2yJt5cxlBf/48EL8QOI5IwfW
SmkfFFwpW6z231fAoM2o5r9LrwyzhXm6sTNHLPVwH/MbQxdR+mluhV3GF0RbTqOt
c6J5qsFfewjq7HILQYSc95rkKzXYIrNzTG14PtDabSn6Z2kmebDCVaCKmNUJajUB
PdHIGG2KGiEl4L6P12MJPdSN1CrnlrAaI0gqtNHpf4HkjbceyVGEKrskXWyr4Wmj
CmH3E8YqyC2l5Heuu2EzpzMCJehuG/a0jJK6pfPFzl11VjlylkukKH2bOS/FhKmA
5QHtf72lC3KpaIx4uJFpCZg6Il+KvnlHB6LWiYo4RbqLZvI53+J7naibQn/qj4fG
wTRNgi2MuyrEOwgsUZdz00Snc8WOgNor5ch1LMRo8wxj+Vc1MMqACVYFJaSnlK2V
GnMsyt3sS34t1GDhqyINoRMf2vOtpd8TyT2T30DE+BTW3+zSFexbd7HukE86a35N
KsaurYXO7dOMM0XpYw2Ze9EYP0fmnPDiG5HKPKgUg0ACOT1C2MaTFo3LbxVmGa10
x4Are4ZXFVe+Pg6uebyVuEqa6i57FYbFT8XGtdrZV6CidER1p43wF2oqJpGIiSbW
d5Gw5d4omnzj/m6yOjgG6wr7XYvJhWeHIncZV13KeZiRFe3WdhAd58QY4JWa7vCw
jdbLXH/+k5AjahcZR3K761TKxVQuz4jKJzeAgKuIcUOkW2qTxG+6sbtmqGqH1t1x
Cs9EN22aCv1XzaPiGtJb/0xV3q+RhLMhkq+cb/OhuoQKOjKKm3y59qmzlwXCTMil
cCSsSRpK6nu0EK9qpRwUE1V3FYlbBzVBJVDA/HrjO6kyNZk00HqJofScGkgHS6Q9
15HtPVpbL8l/5ul1OVtN5+ApLyG3syF3MdvniikZDcjlRbEsaGkSf1/5ssNHYXR3
0K2VTpybW9YMR1S4U5uPG1ym379yBZ23zj72ES66V4w/b7JXLsmhS0w8hMbv8wnH
wJ+m8THRyEcUKVlpO6VP8gbyVgXLbyfxLQ5RnwTGVNXO5URbUvi6HLYMrIxzV5xD
K1tx8Epr+JS+ft3EaC+boL1cAnMaK303pM+ZiQyyPIRsMeXMWjXxOwJWZSol9eRE
w+9E6qOjIZIAP0Xg3vqedtieH5gQHsQsCu3rxKCMzIWq0msusnv7MD0ewMWP0J1j
Zjp2YFFz7b+hsx2c8vz0OGQYNK2/DNlYfawo2rNr4wy1CrCP40Hgp45WvrCv+e+n
Kal8Fe54ZgZBB4Grkv0/35QeNQX4BMwhMMq3Ob3WPQKBmg/0dvNVoTtCXgWkFA3R
JpCPtTp1IhOBvHQ5b0L6c0s9b8rjzj033c2zDNfIbel9/AHulv/yOUEfcMLqtJbL
ljrWJzuEb8BLhWC0PDCqkiNVdcuTShkExiS8KP0P2ONPghBMZFUZ4L1LwbEjU/SA
WdExmyfropFo0HTVJaJRLTqwpkUYPwjrAufzsGdMr2jSNLjhISbs3skcVCuQFZUy
tTqzrZcIUh+WfdvcxP1KbeXmVkNrGBgbN03j29xkJerso9mvxzf+ZRx9rYV/rJDY
rkm/pO9kB1L8impr8e38MXQueUtMmxWyj78NYt6dYGmUHVuDJXwZ1S5FNKr7YH3i
64XSkg3/RhthUzyDojH6PyGD+lLHbUXQo+ntHFsyfjcZ5xNzkNWmA2riwmRKoTPR
btSkxjNPIY2iDd0bPmjWvrjwH5gcxjjZrgjKxZ18V+aaEZQnIEV1dt5MS1IAyKkf
2uqkMz4vM04w4vZPgCctOSIfs5sAyPH67OZ2l6EVLXSZpicbVS868o/ZwpV2SroB
pJ9e3iS8Skd4rtNG9GHKU4Kic1p2/M/tdqAupUeEfwSrv1gnVC2n/kBu8fTLCcwy
nGTZsLm8VAzwKzl+bbjaDFSL3woOwwamRIflsSnW6xBVReZ2Uvc5CUPlexFj6qwk
MYx3WaiRYo9GzxJTM14+ff9JDC2ctOlY43znoTlyNpV6hWvKKKZq8YaT4U9nIjDA
qwm8nRRjdOOf3Q8lachmY8rovVp4NctcoNI8oruRnyvgoq+1YarTI/S7UDnoGBqu
B3aVPLraRQFIuXPr8QCz4CK87jj/Du6CPkxJ3s1beRbcyAiLlYmf6uplT+fzQWhp
RGxnzhOLNVEY/uGJInM0I1NSDBgqkN61ck3DBZeE1SUHCxQgJSl484CNgtsHabad
7FnxDnW580QZeiattvIO8aTeMKsG+4qogmk/TfBMxMeIIzjmYJYT85O8Etx3rgna
O4aCSj6O2O6koUhOCKu7RmEnZ1UeMeWqlnT0Lw3aIwEMY6s8sYkwp+hL1xZm0uuV
0NYcU1mBd/6uZOBWhuxsTy5PpNLLL3gm6fMBvH+H4Ah3IFmqeOKDVBpLMUy7iN4k
mgjqgKY85vw4EgpxVzaY3WpG59QlyneJ+wAcyKOucItMRr0+9YoQvp6J4FrEePSa
W9ZDJiZvJEl/jbQucY4/PxvL8csuvfhuV0bT/6r9JteQ4pOyyIwtRM8mycED4EQM
t1KIsPJgZPWI/a+39sQyMe/FWIJkcPkhpA2anPCcsx8BBTEWDVBLsAzeL7tt5rHt
ZGdUL7Ge/3uktFHnBIRW1njzHkXEByrxs5nkeZU5ZQJ/iGHxm5G4LowItg5qzSit
2FI/1ruZC0AsP3yEcGDS8u+mmPThg2Vt0BzR6IOtrMe0CsAqCkasZmC+2cWNlAjI
4+bE+e5XBIVHtC8UK28vdSKVTNb2nrbPviYwu20TtTwEtbTyBU9XDiZ2f/GN6qHd
j9scPlnky0FEKTXN3r/avDtvMnvMFD7XIcOBX5oJyoGbQuvfb6Ee+8sQEDWYnGpk
U/bD3ia8CI3PQHLagRIso2GyoT1RIeMhSaCrO4CVKCODO3AFm8+nEMD2B81lcz5l
/knoDyKm1mJYZ8lAEJPnJtlGz5VO26mskN5zj4odbauNfA7PLgt09IwRETkklqtP
7aT16sNsL1iI1RYlKoG4az5si/P4dg2NvWBObnr/OP8AKY4qPGvDGNwECaO8jawU
tW+jJA8o36fB04hvWPTKFnY5yXVGcruIIrXMi3MvCYQ2pFPG4drTUw1QvcSCpMvg
FgUCw7nk6PHzet4Qdr4IOmxe6Gj9U9+lI9/NxvZdBXzVIkRZop+gqkeWc/iIppo1
eyvpV+9oQ/KI7N/0fH2nI0l/ViYYFwJr1lw6QZECCwHJzSIwnFzoqKoMGglnnnZX
6ltm9kPcpPD2rHtdaXVWEPmm9+C1x5UkwM80xgjpksGqyf1K2EG5q6rC+bG1CtZn
8JQbdgHM3NpN0YwiCyVrD+LgpIBpOeDnc9LBY/pgeA0uDRNmUQA5GTA5ZW7sE8i4
pxRThChedcp5Kmjx3CfMijT7dx61D0iFTRy1YgXw4fuYPvdC35cmd8M3lA5mYUs0
xX+JgGPVxStr4qtei7WPUJib6NXRcN2PImZRtwpykKSt3dHuYpSt8UWy7AJaGgZA
Dq7H5eafcoIjL4lHqFZM+XA2XCxjahIi65KjxNyOK978Cv6t+kESJ6/Bbe3lU77U
mCxSZN+ijccAPSHvjBfIi3xpST1KmCnVpdA0TKFUmcJ9Y3YLmepbwy9b7uoRJ1ku
mLsgxrXnbIHG2cdc4dhrRdBPMqFpN+ZM62eOzRWuwnq/ehw+DhDw5zHYjj7CzjbV
pT8C/evYMEr06VNG7aGGHiNVC4b3t/GJ3TT9BRLpJw9OJ8Wj8eHJWzZFQGFMJstP
52CXvjFs992JFV5gBXYEW/Ma36GZ11iKFoMWcTuP8tTXU3MhmfBHo+wkzdolzMCH
gK10tAVP+pvkT57kXuqHIFpjlYRExl4SdWj9ZCt30AodmaHmpKNLMrqM/ZxpxtiX
P9louPeWPGVB2dbQc4YkyFrKE4HdEyrTor6eN6zKoY2asSYA3EKGY9IaBe851/vu
0JMtAzFGyjQj6U7ak3xiZcvdZtTBgddnHf8vjpXjif3DIKKsz4/Wwc7ABiMN0YhP
TVwW0veYqfQXeFDeI//NUAweH0QmzRx4pMVBE4LRj9Uyj7lXK0BvfE4G08EGAizY
0cAmKPQUOvIFWSEK5DRe4s7zoO98U9tYcZq6XrHVXPKi18fGNn1O43QUQbqT+kJp
ReDUW6Ai43aWa2F5vCTwBccKem7+EDi0Gd3o+s3j4EZMjcQe0/Eysfk0++FmMHO5
vLA3h7s8kl9EKmQDWwet6HIgbxZKYLgFcj3qmA7KCGq+ud6HMUQwKGt6QIHDRgcZ
hWoIJLb1yKW5ZW3kZB2s2m7sE+9NPnfq+hTA+4JB5IgY5lrqh6E+5cpXLYLjjKLp
AFsea4KdRoHstoXBeditnp7cnUlZj618LAY6ZvjMUfrdMhH2GcHF2O3f3AiFWEm5
aJAUzWAg5vEuFyahelN7eZj8FCxD1hBnm9wOpEPJCR8hD16XIuyqCF78RkCVRvSG
AAfOQhZNZbNXSU7oFNjY4MSozohlVDbadyf2NJ402JME4qgXblNe8AHbYamXxk0+
oYn+n6ycqgQzXDpedX8fBK6NvEYPKAxhhUPUwfBJtOtjmBF2s1oVDu9uISVTqlkI
502XQ1URzcG2trhX7rsnYtK87XKtY2/CF0RRYouirS9yrm7d61nX4JJhaNaP/tU9
rI6U7yCls1r8ERvZBOrQO0uTW+DBMgY/w4XPt6WIIe3mZTuVx1lYEJwdyBm2s4Aq
SPn+x+vzHc6HvUoHR6CIOwNuGnrdIIMGdupW5lYMbDTJSucSUPahC+h4oUTWTIYl
WNpWzdJmcVZCfG+CSwFdyUJCC/LFkcYLgYyl8w8YtuhCZZwQiPmcOSrBheLE733o
fbDQg9FYylSuSEe/L+LTr1ImZWpbluoe3x6TNmcN9prex4l1Pfets74AQpVJeZnZ
oA+Zllgs9IWA9BCYfrKjC56bRrCBlr+WQOLEeqH0Y2dDyuLi8AxGkMT1WaTM0f/q
eB2tk2o1XVwUeHFWkxEKTQ9YYPR8W63o0WazDfyOwP1/xu+3rRkJM7j1PZPaR0bx
AsccaDDAQJjKf+V1K/W9UNoRuRcuYhGAY1BRiAuNNx2AhLYsiHWr+kWarl+qf2ik
CJ9/j+ixqoN8AoXlkTLoTcjHLV4tvkUpg96wgTOPwiQJ2w8TAsM9PCfPSCuQ/Tko
sTJBT3FJ3+9IPBA9S+6xScQbbEeruWw15do/T7wTRAajmHt/mzER5/DM7Md34j+3
NZ5aPjirUbKXTUyzLOoFvGmZnszAXqDybKt3m68ML38l3KO0d98pEjeMF8ayjyS7
kQG9Ajd+uWkofY8O6sEYTfuu83aAr7Y7MaLNez/RURuCK6oelccd8vi+mKKuSMSL
w+81bVFCS40WYvytbC0g9D9n6eocJ1/yhCx/+4iXANCy1JKgcD05Q8RdyA0qX5p4
GmaH3tHEHA8AaFWT/CzALtd3l7kx7cNHGJlTMtCD7REMUadELVmidkOFEdlZQLcV
rUnSaQzBYSfZw2rdgnwhgP+Wpdzc7rfdcfmDlb5IWsIeV9eYPwbkPLhS2wwpgt1p
WPWsTR5O8hgKqGzXbuAGMaNvnEqa684ohBADbcX+r9rxLvv2YE5UlboOni7GenaT
YumBKSdpUXODh0a+JEG2QapiZ1EzVTWGHSV63mgoBgcv15uGwtV+NYCXKpXypmwi
wNQi7LyBFbEPHqEiKh13Go0r0iAUBzsDQdK174eFJlnBSdfv3rbW54rxaOIYYz5a
WHs8+xgosIxE1H/gNk4qgugaRdiQ2RVzevUnlWhw/YztnxncenplWBl1Ep5gQCbL
g/i51kbeqm3r/CMFLu9RWMzK8l3VMW+XAw+ZvhBwtUGRAZAfBOVe3DqXtbc+ho8m
p6v5SxNQraWwzK849aMZt0mqC2Xz35VsqmRnZcz/Aj3dxe4jiyt7gPdPtWtpAQnv
xH12/1vNzj1DrD5YBkEi9a/spLhDn59FIy1BiRxrFRkojU3tnEj+mbRWVq+rKurS
58yXy/0ZZpRP2kV5jNHLm4897Z7bQh4b4K8dxR06xY71+2Anw9QPQML5ssQp4vgh
undL2tIsPH1dcXuWxv7FbRx1stFTzoFjNgwelrlD45QHWjapzLgH5MFe2X2JnDgv
ytnV0R/vOgMmtmFvQTE5nvXu6m+tgxYC6rGmIAUB+9iisa5cfQ4y1j3VqfdSH66O
1nwyQOiPjOJ7Lsgwe2jIwG6xi5zs5t3A7O5P0NW+u1SUxeMvRo10Y4PTdvMhgDIX
KD26UfIUhQ35fyDke+orPx73lCNrq3hdAn8whXv22vrryEAofaB15UAaqrF0EXUB
d6U8kcUCNZRlBOH4T6/tvbfCnwHAhGDc/04eaGmpyvGncq5XjOuoxrh0FXpVIyUJ
c+kMtocS5pic3XD0Oc5xFDqujtiaf69y63DYmwlNzd0Z2Y36FuCQeXECOxG8/ChA
p+aoA01plo6QN46KuOqJogfU0v31qmhvITVHReU+mvBcoNm+SP0pLNR1i18gsNLw
CAy0y3uXlxDVzPja8ZrDgIqBR3SuRVQn6oPHPCGtoZ8J5eAKx/Lg6Eq9LWzdNC4Q
M3bbtc7CCvDScIWSA9SCIZjTWubbs4w2NMcP8X0c5Tv7Us+bayXk6lKoa17APnQn
ewzVMqBkNCcSXRXL/F9IGI9RaAFWU25UMXuv1AP2tJX/uE+2X8t+aQ1TWwdzjSyI
pVuo8rnEyb7zuceJq22z1/IQXXPAHiCbjFcEdZ81CaGS8REikV2gy8GPKyphFVDh
kDpqMDyvNPHdW0YdYrrZsX1seWDeaGuplmRO3U2B/tDooYdyz+qfKEJ1IMd+0ywK
IXgLfoytBn/xtz95IvvXxI0yDdBpri43e/SVxR+otMAKU3QNBCTjtGV7UiUba/la
L9zXBWs/0/QgIPG/r8BExLmmN4EC6mykz5l0EjOkUum54PpJjaCofio/2W2XamPj
ErJlMZpMGvFQlJVR9F6bEKRWqnrGT9yUNZEF2D2cq3pVpmltqfWUrSNm76lWxXso
KTLOVxDQJhDszbpf0hX7VOKi6u8pcmNpvRQwJ16/tUpiO5aYq4zEr/vZq81fZBuI
tZ0+glUD4xjcpI7qixfH3J5NM05xHyzt1s6t/vpbIO7Ay/wZZtlb6il6HqiP28vR
fJN2XYjz/EU1m6epUj4g2wXrI45/vjWmurTmonRxb454JqVc4W3ZGZs8Y7v/ysip
palkpMVWQWVnIt5smx1HuLne7LWzTtTZruDIpCjYmDTp1OIGVp8l0UzpmQp/qmb6
II0ekl8Fi17myZafnM07v+0M/LefeNEOs597iNOCtHNxufDqgufNvjyLD0J9D5Jz
Agj78uEfLYBMZ7vwtefnho2q/3qBJKEwIbVjbY4831Sh+196WRpRqvs6VEb8XuJ6
UTEN5urOz8AjnKi5depQmpzRH3G3bLAHb0hqHrJQCBnCurh4A3/FgY0OrsN3LxsA
7wMf4DCGp3CAW+6CaQfVrY5QdECFJXmrpkAA0wcoxdxsSEt2aWxH8lV9nCEh8QOv
G8Ua5zmJnn8FTbz3S+1fiE+fGMUjsJrbiPmc6pnbbXDiMTfDPdDNa4QVxQtaC8PH
9Q0G0uomozsi1fd9mkrEgaiXCwVmS5UBILsttp3HxQEvjIltygOd2xCKwCe2yfmq
OjlwKqllUEgoO4RnLbBgPOqzH4Kb+9ImKv5IpUoirTxHfFeyra/r5HPfLSiq6K9+
lmXBSseFuRmJ6yrnSN9XY7Y9dx9K6UqEIRA4za/iGGutjyg+VTx+aVVmjipPwYe5
kumRGwx+BB4TZymTiVtEzxQ0GLI5R01idIFmdCyuRz21V5pl7WuA58IhIX/AQfq8
e/hpB7MJM0k106LwIdlaDM1or8jpjoUT8DV4yrcYIjHvUtlYGGau14Otanbbi5Nf
H1deKEj5OUbKWt7th/hRA7aQsWAzWOBAELi9TTiU2yE3IIZh7Vw4XvS5EEhSIzIK
ms547e22grM+N0D4kPPvIXYgksuilyhOqHyL/sHfblKbQpTo9AwOTQUbT7eI0Pam
XoStr1S2xxvupO3sYK6XGa5HXrADC3q+OwM0kRfKSPfFCh3qUds8cDaNlxF2+09N
qUUZvZLdGdiYZFeRLIogjHHwyjBh1yIdjGqlKi5cePvOqU+uILn0A21WHfTE18vc
aquKiwAC8k0wEq3htQyJPX9KI74hJ/1qBtFdkTK+A7mzzA4+FcVe6kBM6/JLxUJz
3eC2CdEzemaNlYfCfZQhozTF0yST5wnDh4jm5PL0Sm0lGnjNIvorVcQPM2uG4KmT
+/kaM3QyYWlyKZgf0fd0Aa7FdmpQ8c3l4eODmD2yJVlZDP28W2iXV6+zM2YsYL2y
P/6BovvLehNgc0hQtyJKOGCduReiNzoDQalK0mbXnmrjpjFpefAgghuvhGdHLrSL
sjHJakGRBc0kn5yKpiLEZUVOEalhpbD9GCRfCIHIUABW/PRHJx7VBkBgqllsnknt
jYjW5MndKp/6Hr982vytipD7N2+PwMpW5S4t7JEcdXbuAlAMIopJKMpgrBhAkhwC
XYSMhCWB+JbGd1HrTeoCxG8B7kYd21QG3xhR5DMAlFeqfLlVBFWkNZJYD+i0pLAk
8oW6yrQ/jVaZtdmqhRTNIMFlz4cJYGFiIRw5aES+90/RpFo0Wdb7aMw4vhrI7u9q
esx1sMFJkPfos2ld4wap27opy7I70M+/9zTmD+Ksd3ntWLsz3O5CaYn5MjZQcMRi
hz0x/4SN94owGfTrfDqqp0BZ70lOqiN1yS8mH/1rBEbKEhgQobhaHXvZ6kq+GcAW
MGn0uNjR6bxbRcyqJ1wIgUIZHbHOjGizYVfnlvYmL7sRQ7su2a7zKzmsXN9E4Hgy
wz+xYASOIQgWinLYEvpXHvpARbf1u6aJr22Xdc+BYkOkhqEjTA7MST+vedEPuT/J
01f+MViRBY0sN8Om86mGgvxM9pz/OfDZpBZ0BU+LeyiB3EZm7cgMdzbxHcoHKiP0
9cFeCtuqfaYY+1oxFh8RYmph+ZMdyC5Q4sFVWd8kU5IJtm8YnLzyL5n4lKZSFIWH
wtHyuGx8XXS9kFZ1iCRfVYmd/iS94Nx/DFGLe2DiPQzuIys2ybKdBwp8Bw6ImYzs
rXKc3e89mVlodZKxp5/bF56DubWlRkriSgl50aF6utSdqqkTUmpb4oPWYzh/U4DW
+nMtVfvYM/EQJhPPAMw2Y/e70/xRBKtm2vfTQadF6wm/3l+5G2vrvaMvfNUoIHDR
SlZcO16EuzOTZW2zifaVgVr7xbLkSjicsn7i3xg6wdCsMdWNfM1GFi0p502Z2FL1
SkkN2TpcSYa7GadXtXOuDPqOCOLuqQxgwqYy5sdZdi0CrbmpFlhGbqQYYHEU3nHT
TK2WzamCk1T482eoDqqyEEKCGhE2fR/UOIWL3kccRw8NON/Hvaid1COR3Vp7C4de
WRwQzGN9KEQFttCrNy+TTffL9uh9JW5cytwY/ImUT0ZzH0dKhDBEt+vXMzQvjYhk
eH7pTQGo6HRNGTRn2eAFBMfKHZP4fldzIOm2uXGYXAYLLQm5ngmdfY/8ZNysWnTz
rVZQSBaTxO/0ZOLBGGBVXvcTbcXS+a/YMaSc3xVaNp9dDrfwXyyiTAFT+IejPEJg
T5dXIZsymUG/4iYWJ8sCpi/z3NSa2I+A0EjV00+k8gpKM7EiPpaDogqtlXudFTfv
rTylcuGQ854OPVbO3HdnwgY4Zn3YG+hmmhiXHRttdUF8sMGmdV9NDHL0ZrGPfEro
q3ecs2QT3dpoYJzH9aCG2So1tLf755U40AY/IW3tQcfZ4ArPxpsgO9PnH6CYFAEj
BvTwo9zIAIMUjb8WI8wM+HIq0QnQJkoIin3/36KeB9c7wuxoH8SEagPdIOPsueWx
poIiOltabknnZzI45c1EnOWH8YSw//7XMrWP4I6TOaAxIOShxlyCsXoAs4v7aQES
D3DdHCzwQNeubEFR8QaL3LagLA1tiB7yrxSM2UDmMKJ2e6t22g/esF3JSFt5tOMU
/UWg7/jxBTtg0fuos3b82/u5oCobpK0YfYYSrsZaBamLaDbFJuTLyu9u1zmAavQa
rW4Pieepb17eiMH17t1AYIRCiISmyqQXhNjJY6OTHBTocDvNt4MzNwVxFWCNA/Oz
reiJYhST49P6xbn7p09YGfKDmgSaI6oJtA+I57HW2ZWCn5TbKyAiwsvtmX/U4MGs
g6hB9Xn7Ylg1z4giCDOWbJsjFCIbaRexgZViJVfZ3D+4fUrbg71X6HqCDn6AoPsY
EmeEnFBgVzk+icCI7UwvYGoD6tBRH0CyF3+UiFHvbCsUmU+bd1PSxt2z7vGmThk+
dT/yqlnLglWKVD0qSJIyUqug1JE5tfvzsqaUgeR0UT17HM2wq39cODcrcQUeN8sU
AsD/CGchvLEk/En4zGx0UXkAE4NT7S+UOgAWhw7FgbouRWrLZ4v7gapM/EZNMuHY
NMJyh697JuasomkWE8/Bq481JbPFtQFiPiF5ETF2iMWlK3hhd9UMde1CKJ2pLUNm
Tl/rY5zttkxPYrGg8/O7hjFHYcBP1ycF4f0FwRRH3f5gj8+FVTqzrP9Mw2yqAPwu
iRZQeKCjlvRDNrTjRvwP7vZeKf7t9i+HifpQT4nVK433Pn8Uqpbft8aANHqoFsrS
JwBQ+/4JAA1mqb0MKUv3zoUWhXZ58UVCG48C6fdvOXnQX1Jxlua+pmoBLxTnt5nF
2MDDgVviA6c+uqrINTFeptiD7kIQ0Vc60xTPs22tefBUP3AaT4XAgvhUqFsriro4
1MVrTm4DZV9prtsASREzpy2VOKJckshhOVcoGChEbKeXokd6iZl/hVV1saBdyBXY
+TCxQimvA8KQ17fXEHpguDJgyi902xcQrsT5U21wx38AkS77XUix3miDVkMymWYV
G5TDXxA4+JbFfGjrKIuLBPxKP9phKPnwotLznv/JtsLhj8VKpvq+a2+4jgXesLRO
f2ggJKlf8y9ZMQVBikABs4M0+sDggedr2S9yk/sZ54hSPPOazrfoRETvGjUIVbZi
Mx+rTnRQgeou2jggFc2xxgUv6NN90dWKe8W+2Q6G8pl9d31z4wnNZGt3I7XyW4B4
pMCokBypF12GqYKBOolnjtCKGLlNL2+pPvpi4O65X6fnzRV8tU8CQUFWEXX2q4zH
EfzdftUjr19DzV1lDat5CbuQbWLZxKF5wl0YQ1fT0RCcfVby1tXopGkHkeD0d3OT
gSWvuYSsGHjxto8wMI8r9ES84Vde0keNwkbDN05LlkagTp+VpE7IQzCvSDz5S0jX
DeMeSLUTWylYPonIHUbagFhTLOp2iEW/5L4wbvsJALG92/HkYzZG8QPSJWR0waFs
lRu/BmeUi7+CxOKWZY47uGBfu0SP/6G2spAvL66sq0b5WQzBGcys6R6MgARzkLUG
yzwGo7Ny3Lzt1h3A7x+6cZlntn9XHvIR6FnKSLfehlJfMPGD61ptx9SWWGtpykDc
VgB/0IXcQMTlWdHtzH1ZJne/Q5zxGkbB8hn5Um9V/h1aAlGXg46WZZtl6BpetEaY
esH2ZUn8NUHBHPTU+cMy1WcuBh0i/WKQskua/yYV0G7S7dL8dzKAmMNTJ0plAbvH
hygyxO3TUTmnSL+U4YtNoMkfsVEStB2cWn8X7LeHEFznNjTsYQ5QJE65aK8rxxYN
wOR5dxUhSl5ALWrYT1VwSdcGHZzth0Nw1BvPXd8c2asNBFo2aa2+bMHJTWuP9ylL
pAMJ63oWKX1TBZY6S0wI3ahUmZUBwzCEqUqvQjEQT91RaAr6uW3xhRMLOc9UlRAs
pdGU0wUXCrFb/dMYYFUidvFoNMCCjWMmlMxHAbl3V6T4c/DrIALHjbBWx31wwwcZ
ZQwcb7vuD8i8Se7tWGwzVJNqTaoAFDVRZApnv4BNejysE/oOq4ziwnz9AdmSc8/a
teRV1KZwmyvsWRnlHPpOxSRgHZAIxuuryTHSsJAT7OLYQiUlgM0EiVduBCiqh3AV
nraVnm48Sk5BkMIfZrqQg0oWB6sUao38ef/qBW7yKkQ6B8ghGNqo1Fyo/G18FE/t
BlCZWlO2iwjnbw6sO8i2L0v5q8wqnG3/v+XWXq+5+W9QrzG2jD46pBtO27GfN+ZW
WiS/D8s80jIdy7D92zQOtBNdMxWDfRLq+Hz36rsARspy+3zLgkf6njUiJujmHPX7
MpODvDwEG5DYnNcQWPv3RSWvz20sTX9m0W+t2HfbeDd3lNfxloMSnlcZyChCFXZz
ERcTG7d7Ze4dxxctSsmnnVgBOMEgZ+d+SraNTCHfFK054/6sAQ1UGF3ci0vI31AI
HfYyt3URhQVSrYFzAi5YITtpkpcD+p+RGgVYV7vV9Gi6SIH5UfptArhd35vO+Z7F
Rh6Ldd8lpmgkThTk/dq2Yu6gfa3j2avIkBunLaWkFrUx+Y1BUj5CvS+RAoggnFbR
frJAohVG1/tVAhvWT/Q7NMPjieyba1IHVYQxUsTGQvSQbw4sb81RUtRELR+0G15I
iFxXbsmLm3VtHLtJIrVDr5uTLYLcwOQyrEy5ea0QD952/tsUSmyK5JXx3LcUsKuy
fga7YUvXQAiEZW3GpJh5oKfY0NB3aDdQ6gZ5CYHgtFLsBZeQ38OJjf3LNddS4gPh
4UF3DddCNHuH4Z7o0wG0KgpgyQbqBTz7yf8wsqacwajNmiVqlJDeft3PJEMBx6mw
HmdUcHR9bmAub8IqWIhG9cTqQ8m84BvYv14om9mrHZPdq+52b//vyzn9m35Emp1A
duma46xeyCvilIhUl6luCDyoLxdOIMAulCQoUE6dymP+ozTxFGLaDRVwfl6tKE3I
UX49MYT4hgOQP1VEOVcrmidikL9t3PYlun3ugDdFus5JGq3WkmuVILplgOv3bz5Y
9JhtKfbvLL371aAmc+DypNnUmjR5zRYwucjJqScE11R56bF/WHI+JvtD9OmVUpTh
MrOQABl8n1gSuyT8xNpJFj3dmpFrKmPIPpZsDEZvhZYEpJakBUedBw8aHszguhPT
rGON4pIsWNrpSvPzu6BYN1xyUPDsFp8fD0M3TZA0Cmcfm3ujMm+lRzKzbd/kRPdr
SHzKW1b4HDiA9kN1f3b+YcNK4tv7KgOSEKupTaO635JSbNAKQO1GWpwDO2BiGQo9
SC8nI6c6rtDnnUskhsmCqhg0VzoiUQ+O6WmfRIFCJBE5mPLAUfS2aK8hrSfu+dR9
G/+xG1CM59f2Tms4mbFQEVSW+jlQCVNhcukFibNvuDd6Isgttol9gtJniGrKsihF
UUkmcFeQCzioFTO1H3n6aWagINyfpnZibxA4wS5sI3MRz709vCBVgVbD1G60JyLp
AjLs0SodarCULkOBmO9WTgfCOniOPMwTU88TXlcac8FjgOEvVs/dDZs5BH8xVOEh
ZXPDyBz86jDhX/buV262j+tp28DcIRBJ6asGRhsw+w+nNX3fxgmMmdU8Bhv8YJ3g
NcRV5nNI8Tj9l39GeGtboE6KLfcTo5tp6a0xA5z+8BISzEK7bwI7zof++puD4PTD
Iq96yO88+c2+Jl7SIADIAlhos2P6XLA6Po+R/5sbKKRhN70Iyne+uhLqM6BLJWE2
Z7qH3N2scw0R7KEXCawfCcBnZQiSJN88e21wam8mVwxoUOenm6OGeab/3CaZN/Ae
V9TG43zqtL3Hvspy6BrU5ge55Ey9Zx7XwlChAK+2G+LuTWQLSkQPYnmAJAaTGwIt
dKokbaVlkYQLr7BR+PnqA5jM492/2abbLF0bkqyn2WmQdxljhRbKMHffQ9gKfNO0
lNH3bReJ4flWMSPupOUIV/5Wrm1wHcbJOkbXkFJBh4twIt6wFz2i/0eaA62dHmK9
ZSQVtVb/wzR7Eipb+F/x/Ybw+QeqCEPrFF7sFUllIUgjKsoQHVjrzEmDttAfKSq9
dVBx/O1TvcKrb7HTjtyn3RJWikU7bTqIsX/Ur/fx1mfmuMX9Obra6F1FP4jwSbVf
3kHtv5O2jJ5+/hxlnwDgcMtN5fO/pR5NPAyyIrOrRzqRc7BAScRYpI8OxeSnKz2g
NiLwnvJLUDOklklfOkCR33Ytg76fQ6uIKxzyyUrUgA/VMzfrAhQjCXzpfFFycP9Z
48gh934MTZYWutHzaxM0kMCBSOpcSAEsSKDjRKNwzUnolx7FSr6IXErTozjoTXwr
gzlZVTsUQjMY0rpml/82ganD/AYj0f37F4aXoi/0GfS7sIC2TFHrdwWYyA0wvXeW
jozLCZvTFUeJdAMB4TBTYxLJLbgU74o6dMYQ/hpUZB0+XunfmHRD5M5xKMGQvLiO
fl10H4hlOy/N4z5Fm5h9rrsg1ZTS/Sijge8hwHmLS7vLN+TakAqnEY0A4pOeSsds
+vbK7oxG18gG/GJ7fd7DzqyS29N5D4Fz6cmlELFX6Ym8O1eBPGS+sztaBPYsgHmW
RYY/jL9deRljdnLKW6imOP78st37UVvaM/H9RlYQw26e0JCtccX3+CinFbSE1o/h
3GRsJgsS0PJRAcseDkfn2NQ6DOmoW07Q6U6/hdSnBZn9peS+jSbYpU4T5Wchspka
jv3X0F1EPStY4cGLnsOfIMKjLo9GY4cKrwwxH71NANqnEFEHpHNvqDRVymZlpyEE
KuBrjRsz9f4vFu+sefnNrj4Nv8eiMTU75lGXoeISGEzmEViwbQnLw3oBevXFC9j2
ozsDau5znFVA1F7Yp0qS13ZsW7vcHVR+6as8dUJlt+Ilyd3fk7F92wvDZwDmIoTV
Px55iquGzKv7YIo+CRHQKQTl7Z6LWb3k4aK0xrLX5Iy7SRorI/cA5aVFCK8nq6lM
An28xdNskzzwQci4+bASOy7AOiBKWPf8O25KijaNFRaEdVSY+KV0SMXA4+QW0u7e
xq3Q4fwRz5OgnK1AmZoSvPQGEiOl+9QDXTpGZLbCz8K4C61gnCwY65SS37oauVCs
2GT9RMJvNjOiwqa9lbIBPcDD63QbmqJf0fsyXFPdRIPakp1yJdIUO92ylUlbAd2F
pwljk632WejC49wW/ggo5xLl2YNrtznDzqZjjkkPG/wdE9WsEZa4/UAr7n8EaSa4
HKuml62t/XgnJYzt6xLlg6N5nv8TiTHoLdrX/y4ij7tWAGxU530sBjL0SPcaN2Md
eEXtGhiNWJBk/2ajhrPkYtmidHLsZcN3lJxDMzKtfouv3tZUYu3n+1sJ7LJklBE/
fwf94MX3uDiiS5el9w73ga1cZU7+2KuwzbxVuBCgcldv30p+ogOgojcgkGPIVyNt
bmK6pHHZML+ciQEk6FqY67Y7AXWlv2+QfJEFsIsdQg1wtZdsQXTxcJtaORUQkY66
vIKRnVVR0m/0s5vdylsi+oMhElW/Xo6yDnA8a87v1Pw6F2SXyf+ijGHvayMoXb+Z
964CQvy6ZAkD0l4l8oj5YI8kXUIMWWDQpqbM5DBAoZtI3wpfD3qTTrpY30sX8rao
7gHTfLw4xN4eXvjtKKkTK54e8kJIawNcMIOYaJMibIRcY3x8oZeBJFInRyMKe0eh
Rj4TEStwNB65D5tvfmT5EtNC55rdtQFaAPGVF7BnqAdxQ0FPZvbZuHA8UpKD2VhI
Ro44k4CCTUVoU+tS/ZsJ/ijy81sAleMr5ma4BFon1IffgNCWLxTTjkQT8Vy2RW1j
Is+0hFtfKD/sduthYlujnSaMtsKe/mIV2JXoKe2eZZkxTlo4Na46VVgod+g4m1VA
ee01dmpXW/yGHl/tM9h+J+SqIX9/6YEBgdYrng5UY8dF41v15xBp05pyWued9pra
MeWqPY8O8JpZ5T1G7tFa+jb9Erv79ae5frvl24JaiXFGkf4pyBUWzGrcEMh4ewW0
hwQqkZPlRSiELv9SKQG3iMhefTQLQky8plMcH0nyt7cw7U5IeLKWTeqnWnrR/DVF
i0pKiQYfhC6K3sdMzik/M1lYkU0Gqb6u+2Jv4lftiY9xW4BmGcVgYjNcI5XT0Lbm
8TAd2WvhAEkv7e2fqQ5k1Jxe4g0LNOJoO2GlYn2VmonRrgN4LjeRrIXdoDWnOpL3
F2ZSNeMfQ56QSsiC6x03blm6MVBNRNSciG8FyWkIrHEBniMu1tpijRFAH60y7USQ
Xwts2oFSMiQ5D+chSg7Q/eArtXtv6xnXetYhj+gYYdcEZzW+MH3J1xN5dAxkFhp9
Tv5rvsDN1JxJBoOft17xc10cqjOEl9hWyrI9dSX/fG/Lr6oK0jhakWncxXy6gf4p
YDx+1zlhZrOMmmauTx0zmt5SUq23rYqsUKVnFd4UTiuFLhG9bjTnw30qZ11WIFcG
aYNqSfbfWEgq0i6/mzdv4tMUhDQJCLKQuK06WRSyCWLDFVE2qaEUtfjYsRxpqpEP
0+Gv1m2koR9VhjJMeVJGvYbIU+9I2EBP1rrFvZBd7Bvby6AXfXtlNSX/FiLL7jSz
jvEzBeT9/iOnmJ8Wmeyik0Z+Ltm4XntL32BiNg0jPPHD3tpIvqaU7mCbhvbWSx8e
7lbm2/E/4isQmh48tcIjGloDW81NxMKJ1WevAThbe8iXiOkKMOFTObIgHJq5/YAb
V9DLGWyM5It8w4B3Yv3OaMZr/E/53tThRq79KUSjpJUDW8ICzqZa56HbKhgQeUsw
hEYwl9Ljn9uJkb0IOut/9OduJNGX5RK1fAIomFp8Dd0EGgzqGhPeTbiIQGTBOaxV
FWLjmJu944trNCfRUwZzO58ARCWf6GmvB42oqj7KzwJf6+bIt9EqFLjN5RuBUBEc
mRbnK87cQI2FWNI5PKMU5v1dZ7TDasW2GQmvmGBou9Sx4GUseNBzg/QYXRBmeMo2
xuvPOL4/4f8CG9Z5r/3UnF577+lwWHpVbifJAMbAf6BBkv957Y+Fcmn39BG2/xHZ
Nbabeos8CxRes+szO1q799Wwws55ZdqeaXP/RAv/9o3vNpQmsEE+NwE/V1odaj4D
sgJk4nasaTgbekUi0H5jAyFO3EhnAR3DxFNdJzAHNNMpullskX3RBCrjnlY2whJt
HIYg9Ba1K2bn6h93eHzyWCyPZ49ax234oHY3e28wnBdLC61Az1ywV3vX3Hv5GdxZ
mGnzF+wsCVp0f0LAvmlRLfgSnTxnC0nhR9wOMg06ehnSWoRbkTxQtnYm7vgHzOt2
tp8m5cJA2f/0tETibz6g2LzQBuV2pB1dnOi5seRLdWAq43rM56VU4wA5fuv9vqbK
aaddydRjGB+x4y59r6DTJxPLbfqiozhuAUH11b7e/VDhb7AKng+8lfxXLAz3MXEA
QyoR/X7z58XqSV+ysBdasNEmSKriKSr/5I+WKG7vGFefLP/7YBAyrbivPMQp/j6j
Q67rci9MKrXanjrCJf0/st9GycvA9y0EIrxi4tMrrcIWAhmjsHoNJ0rBCbtZhebI
EPxeGggpzY72ssy0u8gz/fEKTpxNEUNqbeAa2muoX7fECqoL1j+o6vfbjefMCgpJ
VoBhTehoN7OEmgxUc0Y7T+qGOL6CIqBG3ECLYOPAqFiKkKpA4biXFtC6z+5uBJFn
F89+IZYToYVLeHZ9jaaj7/lLmYIsHVJSu8uQfHL6ftBirrDeLWhZMAnpIsD58Jcg
oOJK4dW5/ngELR7XjazksZpIMiNUj3Skx4r2hekNxyqJNWspnmrLg6i2AAqWJsId
iKdGPWOXdMhggGiboxIE4SuUPJ7yaItOik5e/obA5IIRbrvetzO5oOJ1LAxJpk8I
QPFZrghCF+VANRQMUGYfAlwwSdsnjieiDoWLFG+Es/c/Qw33KKw6RDm2HwP3457m
EdTozk6QaITGDYhlt4l+NwWwAGqFeZXTN/7jrJt6mnSz0cN/Ogp1j3+m8eHjM7VG
NlbTqKaU+28EKPvXkVE8KeNZXvOqlPQlHSL7xyzyS/mypFruhcQNVE5BTT9Q76re
XbFXJO4oc06an07deS+JEni3InrxxQHxJPf4CKuuPY5rrlvYNAeIBu1/H8dwpzAa
zwBCUp93IUvR5ayq/q88CG9K9C0sL0Eo3hNMciAJrl8iE1LoMMGIruR3bWnaBPG7
iB5Xl5Y6aLE9ZP/JJSo9AxAUuE3FlRvk7HA7ixJV7FMepj1dD1hZev1hT/UrQBW9
SEIDBJ5yFQciv21ZS/IxbZwTVIC9SEjNthNl5h912UROaf8/MmDhm2HiQb/MUB5y
JZlolo265hx2ph4uTIE9dXk+TAd4Oqtwwokg1f3YUHKl5/cLh5/i8efbUzWnffL3
mMiekJSO9ZtVGkZzkvubgH5RnhnIDBSESQh+sh60lGfpcfFd37zcbzVla8sMm2Jo
LE74c3Edmm5YS8uCsxPI4n9ksQADaqq5/wTvGNzOHElYljptfwj16XtYqSu+JS1O
gxQVBgXB1Y2g07rwJSKhGY+1MCPxDDEObSXjet8cuv0nWSEDh6+w20bxfIbkPc4I
gENLJa/guqUaATaCzrvsKC1w90KG4nBAgVs1tCmWtXRImnShc8ssOjTq2WZAAD9u
6Um/E1chH3PDDEaBOJY8aAjuW59QlFrgGLorYqZR8ypculksV4xCca13efSomlFz
TZPecQEYMHoBkEJseZ0aZOV4Z3IFY8j3Gleni/xNWDyPKQ4HO9PAD6MUEDSz/poK
Gle1d+E0MKO89JDQUwxyUBHKP38yg7+D/HsrhnTr/T2P5SdNRdxZWBpucg9kz5u5
GW5pkUjFzUgEv09UbOztJw2Soxntbbn1KVH9jp5ZSaEOrPJJXm8l987Gk7Ks9Gad
2iXgx3ymBKvy5KmFRGEtu5Csrcw26bJm2RxTnNNLeFnemHdUsuhkP423boCxp9p5
A1QuiKfs4c/UYZ9AIIUOocN/tC0T9VtkH9aTERvTPqpiIS37vIz6tB1OmF7+t40L
GwmGgOsNUHyY5lVi2uFk9mLnXq8Mgp1N2eOMzqd+6YmVIvndantilW6TtTXJT89Y
/m2UJ4JcW5mDNgEhBBehEHd7+YiOhKY/pjkyYolF/iP8IFfS7f5SJtpb8IOBQ9JH
TgDBMGNsD9FT/o5XtOmSwbSz87cHh5iL6Qg0Yb2YE628zpz4gPK+Jaw1+zzQh0MD
u3hhlcUzrq+GxmgQrf9eonMWFWqO0l3mu6CjC5C6JuOyCc72pqGAWaiVAPwy+1o2
qp+jpnep1Uvo+KpGRE6dQl2pSXvRQTOR0Yanv4mmf1d/cxN+0DABnJ0BeKI+TT87
7oyUwShg/DNeHNVoSZ7WVrj08r5NzelcBGjA/ydt73B2UvhWuJRmpY/TMflqw4X6
vsP0I3i6SSVsBsxVfyntwy9MkwRvQLVlD5jyN9yhXi5PrbhAlXJhk7NvuSn7X6hR
st4uIRgguQJBKeVFgSuk4ILNXaJDuYOowPZThspjKhQIIXAFo7dp2MZW4ynpGKmd
8Zis8qqFT8yQ2tRucWuBVsVJRjVaMoeVz3Gv0NL+HZRnn/BJldeuMt2D14kqys3v
VNOZ9IbWB0Wz3D4o328n3ZAAAo7123sWraDrJ+eqMrOq7MBbvlhNjDLMrYfZVyeK
VI/J4t9fZJ/T5J1zZKOQmLEjW384RilesFfjNaTwAREfSEbCPi6dH7aI5gazIMyc
q9iZY+9MEhpJEqLuVsW5IuhmwbVRQCMtt52zdZ3kyhOZ7XiFDcJQgrFOThG5iMsJ
uhNFtHkC4hKDDa+2OFNN5HegIzTd060Rbh3fzuRxcoRbYKIifeVuMTLpu7OtLmya
apECk5Xuh8hyMY526GcjhB4u/p5R9pmSZaD4YFTkL6oldTLc0FnabQ7xz6SEMnHk
oN+3w3z47h5gkHwmYIGp6V2qRz0aKUU9i4TrTewuYFIE+7re/A6GBmjXzikdJ5W5
HaDoWwq526oxoBBx/rAIOBs3PYqdkiy9ssVuraF8oh1subZzta6gk4cNGerka/Fp
sDPpo0Is3X+sXAUa5zWCpMV/zmcJZ6mbxocbqmFFXndpMnO4uDT8+frrYUBaKHRV
HiRrHwlTF/l9se7I9TxOB3dmeru6TFIJWQflwxOvNeGm8DefSRhjhbQGZLtfhRHd
fRcD75qVu/6qS7oYxMV0a6+z0jbJryqCEaOtUlTM4BaHGs+RnxyBHD/4io/zYisj
AuW6lkSuvu69RqLZUW0OnqSAeGDOeGwCGl7rr/l73ec+5DeAFaQ1qG7E1n5hu+zr
Vxe2Fnh0gG3mwwx0NCKhjYuzRfQJzsvzqgKtbdXhiTEg8lXfx5f6vdGedM8lirkB
qStqhRfbr7GBFIOoW5DP2fYnFRenRha32Oj/peT8rNIBwNVw8hrU5v+TjqPnY1Vi
VB3viM4CqCheJCv60zMkE8w+x3zPMKD7ie/mA2gu5kZEwmkVp0dvjvgDl8yQP+i/
toBPThnBBmuPe5QKyqWpo95TfdCqI+qBgRvvZoq8JdPdYKPtkpFK5aym95F3kgoS
+RUrqwkAsxuPrVSVErbB2xGSAlezQXSaPpufVwukP+4YcuRabVREkyeCKgxKsjwW
F4QjpO4hk+xRe0cjxyW74PkxKmEEDw313DeLKP/oKjYJoQHssCyZnHmrQt4HAAk6
I4wAPbknIawrZ7twpxASG2LJoyN1PnxwOyJ9F/ky4ZXQ0eLqHM78IXY2/83aDSo5
brhM9kPy4zbKqoOXgknN2orfTO2JedWSXQwsMrlv/kmb2SR6aK3GjqRIOexBKjIS
pvBKUYWGNo/pCKA6V68pvx9/1oaELwjcghdqlkgsZNsxzAGadmrClu2jugim4fhR
77Y/1F9DTdHwU4AdA06Za7flNUoBBSjkXEceZ3Bg14SANhV9wW7Taemy9WDPakRh
u5RhxPH4D6Qo4A58K3oijqrkNi+zHiSfzrlSioCbYOd9qvOxhg/09Swr3Z+vXuYR
k0JUJnk47PXlH+8M55Qy4Z2rIBNcRZxYcyMt1KkqhWB45Glq3uD1boCzXtfy8uJO
DozMvdGxJik+unNav169OQvCMuCI0UaoZYCW8cAlnFdN/ou08LZVErGh32+Hev0/
rY8O5s/GH8MQtWnAN9B5sVia/4BVnTI/gIBw14UWN+srXrMBRdEW4Jd2rfYy9aFM
5eklPh2/WmXoS9C2c0WRz1tBvUXxcFonKHAYkPQQrFW/svWBbK+oqmy1Qdq78XDP
s5pMuLQ13qXcVJZkMcRI09sjgYhTjLkLrms3EgFQDea4hjoDWxqJbwYFFt7GDeyC
HHSWa9pAUzG+d3oSyp/s/jFMDKmaCvdlwD17oDRt0zwAUaXYmO25fLwW/eX7h0Jx
yzJZtAxWf49uU1JgWXQzBYGL7v8jC5FGyeHmBkQh7kfGokZ+dpqgbU6d5Unl8e+4
smJOpoAsRI4hKiGZ8uy8e5yDhHb7rxqUKHzLf29nQUBdu+RmTqfTw7bJiYBgVnCW
meUj/YdRd3LpCf8sPzKae+qQp2wNn25lNf3F7DTRR99Y5L1oNVcYOx4KF7z0+29Q
WkvaPG6irSgyzCojb9Kqp0ebYLzWjpQ4d1pMyHFT9LdfhzlG71N0OCFvmG3eCZ/c
mgPYFjCmT3jbETcCJ6EtrmEnJgS2FG4ivZNpbI+KbV6dxsXNLoRG54j3JFJmHAj8
HuZeFACzz3ymGsyWCtFtrA+e8IkxtJYWC143ZlnVsh+1X2Rax9Ecj84/Q9utvZdu
vgvK9tI/0wj+jhS9nHM9oeP0qcGXN4hHRF22dDVf4ltRAgD8wRPOUp+Q1fpF/Vxa
R6UVR7lKGpHu3l9+2d/I/Q97lVUAM45UGxBUYZPw5kb8laaLnwg98Hf9xAaeh6DQ
CLggb/ZFCztTU0SBPwz77CxZyMeBD1cfyZ8bBD4a9s1M+4sf8aFP9ooM4kwl/p3j
f95pJO8tee0vYLJK0k0L+7L3xDa9wWkLFtnF36t2jaXd5ppt+rXLJb3wqme0XV5u
Ub3jmMbKazFUOJ96N4wqBdiC/aY5yfYXkdxQl/5D2N+YHZZ+F3qFQ7fK9SafiQNt
t6ElY0Wp8KqfAG3pQt7TrRls5HxcWRijCqpX0ACzctS0hnBpajXAlGgdXFIKW50d
606HdwNACJNYwwdFGvzdZYAp4vu00HYucALWFHfsRPDF9Iwr4mcL2PhuvLnybGgT
ZQOihyBPhOr/xFyATX+YKPG9NOI/GL/KvNOoNBCgoMLCWN2X78bDLllkhDCwLxHv
trKQieeCGbKk3lRD58NRbXPSFbm0ss/hDFrnDFWs4XG/vMmNDOsNU5msqgYBJqZr
TxZ6Y28o4QC4wDCzH2m01uRjAuRjpxPoJQClWaNyO03ASUwGi2g4fqTUbBv6O+09
PwPO1QQeD2NT2gEARdnz2jxnroPeFriSCAX7oW3fECObKoH5+GVmgDJPX4MSPo7n
CCRtLN1lLN55zkknheMvWGFJqwN7git5HxJW3kSQDTrMDcXbkjLHoDUiSF6Zrm4V
e3YW3UKyoxdYKQgNdn0pfKTwOl6GUN5ejI2wFlU3JP3jeTMrfJxl6Pn5VPNaibFG
ez7z7yXIK3/9gfUGpm+LyvSvk1oqmBmB9sUdGWKSq/or30b1lYSu/AJ3OYbkQFHr
vWyb0qovnQW/OsxkIo8kHhR7+ALWpT0oRkFJxARtbbBrvHUNNNv/osZJepVZH6lT
S7qehAA0BxyloIjYh+X8qsYithOZCSH4r1lVuoEvNr+v4JM/VRGUWTULP4oH+zOA
T+wY2wwShHC1QhK3wrIwAHhjmae+Ys5nrKg1iBj7pd3O64XLaU9OJ7O3NeSLEsqj
lUS4iB9AiRFWxaOOWGZePCxZdr1pasgH0B5U5U9J3Y1OTZ5yGhj335l8/mQO9/p9
/qU0vHmQX3MO08Euh5hKKuCfLgSQAvXJOtB1zuzMguAOcC6nkItjnDTDuwtnaIRE
2wm89qIrWSSWJ+6+RdKiMdG50wbdGt/2Z8zgmxHV9DlZxec5dve2aNX8WsEms7go
kst69yB0VqqFfBEwS+A99po3p4Ya6IdqDq9mzgqLTsS0sJY9w/PKYfF/YHDQfxY2
x/HsqlWuZUkj6D/bC+gmxMk3+4N2jsv4MHyVcHKuuY5zStBF3B+yux29C8IAkuQx
MMojxKay69aHRBnD8du+SuA1ZSwldYaqJ5xsrui2Evkley+/Tn4hCG2CdkYrHScW
Gpdf7ubQdYD11x4YnfMaR/SbZfWc8rsw+sVQKI+Eq8/6aS79lPpHf3FBa8Ndi6RD
nIsK2xDf7EK9jJA6KPT2eYZOVgy9EXVDa0P0OcYyM7iLf+ZlLu8izkmFTxXuEnvg
yACnxbP+rAM/YbMh6lbJH0tWjI3l1qF7NEqvmBmWTIdJAGYywIHDf/TOTiz5Qrwk
eAMlm/dbNOl6n4HoGPy3OJvF05wUhhjxAApYIfZRC/0mxdjDKRMoPg8d2k6ZX49Q
WJGeiQmD6xHM8aVmvUxK63qsVl6c5/hSM0AXOPxiYaxjMyXIm2BIJJmVufyWNbxN
f06nOvZN+gSZa+MV6X3H75RV9OfiLJ+jKswL5W7Nu371glAzuZxJhkdF2MxDfyRl
VA1LNcTtovGFxNM5E3h0Xhn3Hih4ErcebMSPmv1mJb/S57qt0VsNAwyOmi+3eboP
38xJJj9matuK1q6Nbw6ZPwEtKUkXQXriBguz5yWzRGTPLQz3kDbesq+RPLrLLcHE
KPhIKBdIUnvWOK+jZtMIf+MZz8IxsLJkRFaOVbsSEXEflu/d6SjUZvRbB/Aw+4RT
a/HLPX6z8eIJPL04IzL5s4mZbfEj9ByvEBlxfJNuwIfRkIY0z3UAJcYsmaTrlKVy
AAVz1NpbSAzlOwlP+l2NWJzwkfLOOOhDuJGTxNohS6vyu5NheiVAY4dN9PQkSmKx
txOpEkZTCbKQirpmGpMQImmV4bLJAhk3dyZ4EQHNUE64TpIvqAE8N7gaFmngSIHf
1/guMLHlzgzCukrg8VG0AkT2LNn6ehy226W3yeHLP+6sJmGeVeNcqw5c8xRIj78S
BJRztdJ4O8nUCzH1eXwXdxVPHrvy4kHJPZC/i/XJ6TqC32pODzi9aX/fXl3DLrqL
DGS3jrx8IsTLFNmHC8ALogDvv3gqPc0TWltjlaJXI+pfQwNFqp7svqLk6EjJrHEq
k++cOy0I1y3GemvZK9FBU5MMOOQdrLjderx/yd58HoylQEA9YcGbI/k5iFndGqEs
fiIRDXr4s7yV8YlRPgIfhccmJTBUbh09j9ihMtfJDgzVAKypjnPNPmCuHZ9etUku
JAg2+JPOoQ6jzXpxPkrKjesXWy//IJKS9jE52dgdSpdKoGQrlISJ74bnxWXU51am
Jae3nhIDc+SyuC0SkjbEnzS22tOXOiXYtDiHPGNT+lZXEZfrmFfHTSeMS2dr+x9s
9EdZ+upMls7TWM2QbqP8a+QsGwUZcm4neVkdM8XIAydhKPF1vxNgA7lczeGClqcn
1TVv+VE22bG2b/PEhQGZI0rg8677ave9uhPiARhEnpNvMriFXcDTjFYAnSg4ptj5
tL1ahSGa6nCGbS8NZ8IKxaMF70boclNkxOltyRdqhbD7tAxrwjKtY0uJWlFumNOX
GtpipxlE0cXRqi5oFgrXUKnhDnHNinBo3vQHnBBdlyN27Mqudw1ZyT9o0HOk30fx
rzo52y78jMLcfobFvonWOGU5NtfTkjhjbX2a1f01JqnhdxGOapKNrAHuUnj5prml
SsxP0z5Dcwb/klS5ovMq2GnPAyYc50n28fK4pWkMzKvTbgOQ3jLljObW/k8eZHDT
EaV0QYBI64Un3Ac6z8vPbUKAlhKsJ1eKTJUNlclwNhkvC9AhF+irm4V1owqTsfut
trHwZxNnYn3QrOOYkKPyGI5cAU5yvXcNx1+TOUpVgx9pXMGX6VAOw93hJnbgo1Yx
8XvZd1/h+SOdzhtV/RcAv18uPZ3c6cbwgf0RWwTsr5mCTcu03/ubWAp0ku96W4mb
P1R9ogTVAM+peo/oPAAgf9nAQi6XvlA0INER1hnGHtCyrPnoxoryE2dOt4HUiLrn
xKz7/MTpTAjjaj6LYdA38xtIMTdE5gzvVOzEaHOp2Ocs1t0RX8JO8TKDInd63k7+
4xduUBFlxJbuHEK9R4zwrRdLsaP42KLLEx5HgfzOsBgXQguAmxn95pOm0ucjatP1
pQ1yMGkIpV+DnPXlWjled2jjUWdcnS4xI/swkKVRglbUzWa+34xm3LxE+vrKq+/E
JGM6Cw6lE4x77FCj+yH4ZXUhkQys9K9cydN2vmT5V7niEApHbNKNd3YIJZ8Pfrp0
9OtAJPny71JBWWW0DC0ZSZZZycJLj2toZhsGkZiRNoxh54iYoMhZCn1ID9elQj7E
qagTVoGoE7NZwLNfiwm8mk/7WtrNJ6qOZ7XLn/v/rjcufKLOZaa+SD/0EDANM0rY
yReFYQpnPFGTHs3CfRi7ZjrV9gTZdkMbgtb445VgVflK+udHUy3XxFtxhFyoZ9lQ
ZNvHFhEUSDag3QsZO9r7Ye8D5bPrh5z7+oPeIKNJGcyjtdS9gFaQ7DtD8pjzh1Gy
56pMUZhDlHqwJckzkvKpBMSDQ6hBpa0uTzZyLnR7fVyeSGU3A6d/t9bnHiuJwERU
KrB3Vkq0kXRxdu95MosRPos2dxf9kJ6z1GnjPufqqPQXE7pZra1Qqb42LkO1JsID
5tDTlc7h2J8l28tUZhw0qQ2nAAN5oOwCssaxtKIjoUEE3QoQ9BzTdPbOBEC5J4Eu
YIOHXkX8z7T4ZI+IGKBMGqWuF/TQAnOkIbk/Anyvbvv1yLYjkDOzgJGREQPPrvO1
oiUiqSIykliv/wZaVRoM82rwdKJk8xAMUNOFmm00VPgSTNjE32qUo/A06QSAiKav
uUWvFM9jEFRLH+Px+P0MsOABFOApMO5yWOMec/22BAa7NmFCSVDP5zChfXnAOqV4
h499oeqZc6SudBBex0Y26WsrfiAzPuoa21RAR0MVO8VvvWzxPnAnVFetU3dT3Tnc
4+veEYp6SnguWHXaX2BazyGdJjft1JHSbwzrcoQlIvW4Xwxghly5o/GtJgWYNnaX
QnEoN2l6YKCxuXqyuLTOMT9lwS5Kvvfykt1R6SiNEhQWBgFIfTO9TXCtmOwPoSej
Sz8sXQDrRP+4m9Fv3vIxmADIZwAtCHpTH1UcZaGSfPs4cbAIL3MZv5DCeUp+psTb
22qwoG/onzyBiHm0yuDLqj2p9BUjwz+VufLD8EPlMnEtvpHsUriZeP1ClGlXDbVI
kfB+4P8nVmYke6/YnskkMehcFpEpTgYLZgZhGRvBvYDFIaJ/2QQGUCeudo0PxJ/p
UJgdwrEXk0uQU2JHdVSM+ZFbonOOXuaNEdaHTUTdSg+f11iBLTp2xItPcATJE1IZ
llJsaVYjhiJ41nApnP/lsnfK/lZvF4qIPYBiF/QhVzRf9aguH7sR+5xmLcxG24yu
0RKQ6+mGpHqes+2UYPoYToCU0Es9JOovYcgTxYr50sSYds+m7lQmAx1gmLj2aUqn
hmjF4JkYmO+TgK8hRflYkqW+zjMKy5MAAQp1jRX5Z6pgeGlvbt0I9pEVuyjlT6UM
3TB9s7725zujFIDpep+zLXyLo1+tcE1ghhqbnRzRLIMTPE/dJUG2+lHEaXepfOF4
tz8sY7gw/y10C2b9SA/bgExZ3WiBGm97+yWhLl+4oAbZlkLW5qaXXIahDL6KMirn
9Lp6wvjuupDSJjOgINP41liSiboXRpzWMZ6wS4y+3HdI7f18v1qVeohXRIMIwHyc
AmE+ZS3O/bOixsGkhpf58Zk13s8qRrt/IHhyMqF7ORdPgmfKquuTxRCXMPtuoyRt
qVnhrcUAZ7X4PWy8jZn3YC6kPDDJ17t2nEMVIFfxO97B16XBGKwAGYSNOrGSSC1h
zC3KGhlepRAPjqUApWvz5d0j5sppwA5kfLvYlwLUJPVjNbaJgqe7cVumqYLcdp6F
2PXD6uoAG3Vr4e3GliOBedMdenR8pl3YSI4/QbDbzAg+0qn1PxHmXHG5MIX/szEo
mOOvaYlNN1Kly1QSBIyckGEC4w3vgpNkOY0xHbsgyTOTmeLvEFQSJaLNVjA4n5DF
M4/Zk2tMwgpfCAVnpEg4i8cBZaCDshDpshLZkrL+dDYGW3ZpECgC/XWsscyWCzDA
CKkefQoYQ9fZBKmJZ65yl4/daXvmAdSy2WAEd1p0Ry/DIYzLZpkyAF2k09Gd50C7
aApmiS/GvQYWmr+cgyrv/3qHjR8ShE6Et+Vnk21sMphcWgQ2Nqeu2e4DYwRs+nyh
QCo+IRnKbMR4RbklUUFQfKfQt2rWMXpl/buAqpg3GNGu4Pac/VCF3JSVsaOX3FDa
PkYhsuJUsT67BX3tmcNngj86q7qZO0hMSTZqvMr6zcKUKLJVjzUgMvaAvtHvxNR7
WNDLNvYeAIIEry9T49MZrcXxmlkRH1LL4m1af9rBBpg7A37ItaHj/6nXyGJ0hK6O
HY2TR4hnyHPNHqxG41DKB3UeLoCrnkmtDoMFuukSS8hi7f1GOUbBY0KK4ryJdXVS
ZvQuLInpEu2ahZ11/XUQp2cDrGHJ5Ji/2k5EfJGuG7o9+qdns/dr+BsvgooZIf06
9wMgwgPBX7OElygquXr55QjTq+YHdwVPWWHA08L3PifPOQ7YDWPlGv8RuSERz8FT
tm3g7Au5e5gGPM9jEvxnhusPyPC5Ej9m2Ax+cDERJAMBagHddrKNmPhGTJv0HqC8
V9ZmksNrLmI8KWBvBLbqi/AmvOENySMKvEhQZMXBm9Lhq3UfGt642bfRJbPmMOgR
2ec1GzkjT3Q90hzj7CL/jpk8NJQdsDTcr8veuVlpOuJOGMxu+o2GCPUM8msQG43W
aEzzB85IO34ZYsgtyI7b+nEkk5bc3VA11i0mPlkYWIwvYbXI18AKt0fF7p3RxCpI
OHOjKia5/UWCfMbdQJopBgOPsFFQ1s4f8SwY04xZqaf3hdz4p6AUnXVV/76x67i8
dDNxnRsDSp0pqKAkMAbKx10CmUNm3MTW9l6fgbQ/M3eT4nx6Qeyw8fAaqEscyw7/
SKlFohiDTDTccuZtDUPHuCu73L4HNwGdW0DNarOE+/FKbNcyWBUJYFrLW6NBueSS
H8cPOx1Q8ZSCdLsl5pbQ9EmoCn9YjpCtjaI+ANN7vE5KLNRsVumBghHF0TTo1uoo
pRATvldTvH0a3hQWzx3nQNjXIuFtw6GE3Q9h2z4yscu/DUIspzZx7Pp2Cd3Md3aj
DGdqMd/IVeAd0UhxYClDdgoayqvUww2BOxuhn0jvFq/Lyo2FBE3laQOSCH9ySY4l
aTmsSZLQhEeKMzf3v1JV/79/gMKa7cqLwzvUAWv9BlEYjw8+An4cOiFBvVlvwy6b
jg0uDrPIm2KDUp5lTLgl3RtLy4ycJ1wkBxvUoNQbrGZ+o6urEw9pB73/M8OhDu87
wNCbsE+SdHZLHdWg6V13NpXvFoPWwFFAcRbB/4ZSa9dXobMTj0dQKcWz++ZyYZqW
9bV0+RK5fFKgA9or/rWOHOG+8acw7ETNhCFtEZzp3z1knZDMGmDFrtgJtvpq9mKD
a2rfEFN7ivylf3Me6cPfLTdBAFOsuKEGVFLljd7knP6tbaG7S0U1oHw2hofpVFDB
MSiCwuEvhOf2LeXQ1Lku1d2YUZyb/xjzaL3aGz4af/bBJYITMdcPXQlBO6W7RS3J
ETqMLHRLDVT8PSeS94NgC+1shOcXxtRYbG6Tmt28FAwKFK5T0UIeQdKkaxv2btMz
YEcYhXDLGFjYFmQdkomynDZYr/pWnqPxxv4mwnN5xr/TwDqBHOP0ex73P6aood31
t5N+c8Kjqlk5ZDU+OwomWmhbpdIFtBlAXtIlfz50McQqhRRtoW051zqyh0ZIkfQX
grcuXzGfP1kUY/Uyo9i1ywW4cIxDdAqt+30UAyMYV6WPSmXDCMDj8U+ECXq00m3b
NVYUPUr0FYXh8GRK2HqlMSzousiQNE7rlRIIzVv48YVpvRXBtk1RpVBCXbZFjuNR
HpE0mtRoYbmFCbN/8QwXhVi9E7SumXPRXnCJh0T74bgZGtbNt3RToqwhjfivkK6b
b9B0iyT2CsEs8JkAgz6fUyOWjQ5st0WaVmxk45EjZsEI90CDmh3S/TvB4ThqAK15
d3es6EspOkFbv2RwfaxqaGFyzFd1x1b/99mv734NZGwvZBwqS8Da2XzX3LbLyEku
kRH1t1+J5UChKeJ7AHuIL8Q3m7yBRArCXNzN5NPlo9RHXxs/Bf3m7Km1siiVKiKO
lEL5aLuSbtVmWfT8dKjHx4g+p5qDcTSlPozcE0QRjHe7R+eaA+USwC4J+llEy6Te
Fmmzw5r9HUxJ6FeMDFKjYGCy2vGYS6VkU+WO6nn4/kOzKw37hMvhZNosjX6RKH60
pd7K7w6eZm6g9r/qjDEPSypQrDv5u6bZoCAgmnOVihs5lusg5jJm+i0XI4UoqxCu
DOgPynk+pnybmqTnBpkfNqNXcHhPD7Pe0QhJ0KmVwG3sh3TQzb2w9jnjGw2TU6RI
PRBVeM8cKXOPLkCPRS5Pc+F9Bc2vKhHtYihVLfK8qY2CQwJQr0MqRCGJJTRpPGtG
XC9pfTTMWdmaRc2e+3aD6lGNdx0BXyL0rpAwP9UfKTirwT90neTVcbnLuMeKBGew
1WvJXPAZi6PpYk7fj5RNQhEkSjrmv2IP3/6JxntcWSs/OPLnRItiWt30H4kCZjWq
WoyUSwTlo50kxZeZWJkckZTpW6c6iWSGGeJ3GZLiyDFOUCPJHNr7LCXZwDiclyRs
7mC09KpKN7GHKJ2V33jfTAgDZJ9FqjVkGdEWvg2z4sOTHX5knCvmeGEwwLLhYG6I
kK8dCwCHLCbGCgN3DU7uH6NZcHse9Z1XC+LdU97cJxjqywnQte7Om7CuLTVGfrBp
eMricEpBV9FwQwzjmkQTFGetJSEAzmTJabV+nsVl12vSYzt64vlx26O/Tb1yKw6x
eG4ptlkfQT67bqCGxHtX5PVNKqqE2FNdJYKfXEKWKvNB8PGUWvXAnXHZLhiPbNhc
+k9X1anweI2bIMK/Bxlzpe27gogrLjd2n87HxtXaLPGcpc8SwlnC/UgiycpBNFHp
OU0ctbZe3MyR/iO8DpE1QbdLmSXL1VsQvPUTFlSHWkEQhb+25ZLA33cdZzdslgwD
VlY1bAbSLDzOXAac1hY9N+ogVoeu1zshkaTcIusSXqGF8EhvRCdJZ64tXb5KjE91
d/qZMVm9jc+WmG1OCe0u5IDWA/V4gXws52e2qLn/JW8=
`pragma protect end_protected
