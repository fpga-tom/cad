// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:46 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RACq0RJxvffKrMIvyagVG68lpaGskvs5ySwOvV4LcptuFVJ9bHYf/wG9okMbgXkI
T3hgG5C7DSdqpkvl/DeoHUZs0xZ8yOwWFGQJBqQisi1El5MO47viJcd4aREazdxZ
MesR/ZZmlAJcEHSjJJbxOM8/4dSO1mY4lMte/QWEEx4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12448)
/w5i5iCjLyAp4K8uLWv4K604bMFch/coidqNpFORrjguJs2TIYoFSP+objiuSTU2
OjMGhZPpWkHOXuwly6E10HkfKpEQOEQDcXbW07ZHBx+Wp8Xo6MyOF3jBvddFrLxa
PdIeqXVScQj2L1euqdsSup/FcGrLlvoWPozHgEihkH2mk/5kzEusE3LqNB/tCH13
DSii/rMJ+S1HOHQO1SjYCaYkuuLTTEsP3/9H024LJSK+BpJKi1hlvDGlC/BW6yOd
QKQTbvAkN4KzxbUUhzcjy0vxHUodP3TcVFlfcZpLjAvDTFNsx9sa4A6YBWlI+EeC
6BRv3nht9iytUuwQwV2bbNgupan3EQFeKHcWDlCWyjgefVswy7S5xLqLOZoEVTcL
4rax/bFiMgUpV8SxTKa1aCIpXeifi67I9tVABVYiyikkVS7Blji0C0Smf69kCaZM
zUCxIu+4jXk4NyeKN+UYrQ4GK0TMVjQAl0wxf/PAYKKodqNH6kVjhguzpR68Z49N
vR7qS5972lBGYs24avpxmek9Xbo8yWX//uznvI3uz7+enPg9TPhBjSKBSD4nPxZN
TlXBKp1VRPio1YejHP2WFHm7yKpdCiVPMIx1LvAeojic81v4Uoc5NvXOiyNCBErx
pibjVGtO00SlXxuW3pMLkjiieIQaJl2rX16lHEI/qUO/kUSgnXpQPyeKQlHvKVOv
sXV4C7etETqzHPbu+szCPgrG1utv1/Lz5y7HlcooXILUhyrOWCWea196wYP6GZaV
vfxjIidCyuXLFRXaRL0+IcvTb6CdUXDyY9kWZykvD90llRaveCGqwDEDNZwsb7Xb
Es+dAYDwpE3FPwe8N2xhWQAavc7aXys+vQru23K+i5sT3FyKpAQ8lvp6H62INE62
P8Gt87rAsZKqEnWSod+k1sOPoH2xPQJQEZLQg46xX52s+0cXjLcQmL+npTxNYuTx
TsDXvCTSduxoP9lHfyPLXWIZsp7xkRSyg+YAXHpACajHMJgLG4V0gBEw3wpsGiAn
YxY4+rCJ0DBwrLlWgd4gr8fsT4DeyYBX9dJhyaONT+qnJdfLWxridSgh2AbQLGVu
BoTipRn12K9jK1i/9pcl8W1dmSLeXHFL4DYJP3G7pwO44gAw6tliAvWrnn4Qc45x
PGTDeyW0y94AG01fdD+FsZGNUJa1dQiel2gQZmebWpF0SFjwHt9qsrms83A0Gafh
dpKtgizRoDtOzvVhFSi1dLhgEurTJtCFNu93CYkMp2TTe3ixn620RWhTso3CWc7C
oUYNmc+esyu8LkKJshH+hLmBXWPXm/aAEJ7y3X0cUVBEk7IdssSUBJCQoqSaOs4W
QoQUbRCVW65v2OjuROoM1qZvlSI7KUik/TPNN0airyVZjtGezSsu2OICH9xINehb
zKmboDp1JXIu3ieCKXdNw4xcTNTmceHEpMF2+tF0/Fkyrfuk32h3P3NhNeiM4Dwc
nqdiWc/zNcdbhsz7rPq5ZrWb8ZLT13b/Zf8GXWl6suRfuIlfj+Y8DabodgmtMHRl
giiKo9x5wg0HKMBsZZk7QsC8vSbAXOrFaVU43yBlqJnptvekJIv3VU1DZujrmOIk
yEXSWNnKptjXqYTL/0V2do44gAOnpjJcdFYfya3biUp039YZL1imwI+RCykGb8TI
qPQ2RuZnRlw2sOsHga4fy2S2h7ZVENGkKZqz5u4HabjAq2MioRaKqw66/vE1pHIu
upKEfGXV277KJAbaDvaoxIuNrfarNW4pYsK1ygXZQ7ChCrvlLJFCYQ4kqz4WU3UA
n56R4fRJAQ8TfHOKApWQ7hcwrx1LBOZMYCESQGd9r3aXPysc3MHr5t154lZz/vnU
wYJX3LuBshWnMheqPzDpucEHApTzL5oOzT6HLdLAbuv2K7U2q3P3qdT12pV8d+MK
qH+MR5eV0q/69EHM8CqiL+BTiYjphvcIR8K3DqsQBKO3tvZVO53OHYYuNNYOTPa6
q3apm+GV9NiTQTfCr0grfGKZfmzMOEgeUb4wErccc6jc0lK8AqmXmjXdDD4dIRDd
KUi1BzLeookCpMsQ1/h7YdC9ufx1qwLHrT38ZtGO8ytLkRmVe7w+QL1j4RoDthxg
Sz8b89tiwg7EItYO6xnXFblchq7+dBg6+vDclw/seMZnHKxs0SCZEcN4hsbTYBoH
yt9WHEG48GgGnA6/kZjpvu6z3LUzoP5YFRw5teENybCqLEKfvjkgEa44iMcRB7uI
bH7fZG5B2d3Odxz7ecgPxle9mp2nKIgfv+6krVuiUJJUqRsjllhIldFc86h4PtUS
CRT3oiaMOpRgqTPnw0ISmbI2vIQ6OsqUaCtxk/Sc3WEcOtCDjx8Nk25JHJhMQ1GT
C99GYdDt5+J5l/ap1oQepP8Ox6+J6S5woN4Wuc/9leqZ+rZdYF2wGNFRtsmDYl3j
tfPtmwruCjOEyK9XvY7eQoo1+gNxwnj6rqL3/CCJdNA7Mlar7/BpXY/vBJMCu7mp
OpC9EbRUJ0x6vay0k8QdUuGXKhogjNsylR9trMfdAp0nL5r54kLKZo6ZwgTfp7yQ
qmiG6aAnftG/S+gSFnLBoEk17RArTKTGFrrpE93HY5k+6Bvlu7ipBc6Edm3vGOEt
ViOOSQQbd/w7QINOYORhWGZL6Eyu709kogWbZ1xUrN1mn6x8MKvj3Mzt25KcxkXw
GzQ33ydDB6LRr2gGg2+5fuSX6uEDe7eeBKjmOsKpVLThEooCBvMjgCvGlO3/gu/8
ylKmDfUBK2PWGlUntGsi/UK9DJd2bHZcXplV41tTzgf3R0JVaPrzhAlRHjuUbm73
eWYewSs7wvT3g/tIk3XMknwP/cZUT2ni6mt0cs5ucVNT2FbYezzHT3qF7vVb65zH
uGjLiuCazBAYNqdp0/OHJss5leMPchEajRWdXJdmKO1+MA6N3dEGuUC5Fn2vlBBw
xgWKW3IfTwDOBtEL43G4zla2/oNvwXUWG6WZiBQHTnVpdLWOPsQik6cdBjPMHhcw
V15oBYvNREsEMkLyRrtsFBeY5EWH9KWxGRoiexTQJ53MyV0sAS1LnW32AoApVqEk
bFS6ku+6nDFm3u+EPOdfi4I6C5qNewvi+JpyH9S4SYk+kujzVWgkbZP4Avk07jZd
uSkuEGNW/Cx7TOK/bUhpBjA+s3THwp9abbtIvEEJ0YCVn2yk4V3stK6yEWN36UtH
sc/utLAq+CsFtPRAlw9kLiYTMWC8C2sP2eKXSJezYQKnOYhtZGI8Ae6XwqtijaqN
CIut4aX78CRMgi1QD8MnFhC3vqtz1VvHbGPcfeIBJ6E4fRhPkTrZLn0R4RocTEf5
6qYdyZUO3BWFy53GHoLKOiSZLkecawS/fBm95TGz+71oCmWHRxXt8X9U9Z+K24o/
t9cEB+TrLcvCmSnV052AssTonM8PgzslZGlOtiQK6jUwvO5a9QlQ+NeD6qfiJ5Vu
YsvEHKCFYh2SnW0oLO0yxVPencXytzA3kQ7CGxcyPGi6aoV/lhSSxH4nfBOKqTPb
60bQAX8MMh/WcDDtJ5F45RR4QDPASqQZsjDGyigzXX2kg7xd3pwtgpe46plW4uFw
VJ6G3ZVu1Tlwe24jn8BJk73H2XX1DoBoDi4+3flFh8Ni9/W/gt5doK3DlZONWBPt
5/QOobGo7/sAAYiBw+VUHaRX9mnDOaw+zWVOiK0yHFkNIyoriWI0un205DLkg5F2
oJhxmwGZoRPztaQauFFFzwXmdfpdrn2PnP9VM1t9UuFazd7b7a0RXRkeYv7Gk0WH
VKdR4WZu0L0+/d7SWDSrpCuORjbMyArENgmHXLukbhDgwJhJs4cGOgq37oeWHMJ8
nxvC+SICIxqZxjf0yDStGkRGRbuVfWkIVfl00UTsBG1jgO8kShDkNxtEo5Zndp7Q
Kkgm15nyHacTgtuxF0CtEeS9Lu1Qne2w4qh5+zGTnXksdJc61+BMbQMQFDbe9vWN
PxPc6ah50rNVvgU/JilxoynK0wCg+oo/fIVYPsnovN9if41DxAHotgzFkLYHEYwb
3wKV0vePNeNf63ATMx6qkIaSzj2omYZlD8/GARD4HHCgcfQ9crb+0xvfRTptbDqL
m18n/KHdntjg+jQxuwH3syPuj+PNLiWQqYRnkx1ZJPwo0LlrNUnnPyfrl3Gtlt1O
GWry5Wv3AUkZsgXUKiL1R0ZsDNvJCvjciL7zBW5jMZHETRdaxRH4Ezn02ceBHI6F
UAdlO6U0YStQUOhCzqA74E+0lXaYm548ms9EomR7IZu2/0TVzlHksONE0bkUXzEf
J3eC+vndWeHy1UR6KuS0B7Dy/NvYhL4d3wLe7DjtaEhMtkfyORZMZwmBgHaEnXKe
CVRYG8A+oY1v11f98cLg2YnjS7j9p9jevxU/vOUMv9+0y1IuXr+VFFazT6K+KAY+
BtSFF0Z2cgUQ5btwLOGfXAxLMSVnGGm6OReEnh7NclcCfIIXJprdUWvJk8ZSsczs
ISNQHzcEFmsvOKQFjzc6LygxXH+zilHuUkPNo+dLbyvfvqskEFSTEsQgbqyryXDN
hsQb+KjSLZ2qZifA8LodGAL18du+vi4rR3z6/7pPzBoomA2Y4vvoT4ud9W/sF7Hi
KFoEXkx1s/8syIL6yXJrwLgxOY7h8mT7veU4+DGzh8McsS6YN0PgsbXS8Cwva2cA
KLC5Es6ONNuOUlyonYOYUNczDXcmSUT757BJbN7izd1zYOC4PlVqBuqfcM4SsfOC
t/y0PznvAmyNTQoMxi9ZE0JB79vbP2qG7EQNMr34O9SfPYiLYZ84UW5AJP61/3Ib
xDqwYZDxZp6ZOIUhQjkUtaRuepFx3O6PRMOoQZlvHgBakbeyIm0n7NpHR3INOaVl
J6aZ5fQEcyNYep2AoJtYAJcWkqBPJgsMbbqHkYl1Erd1wKSxot6fKbgG/5iwg3eH
gYBYbpDxIy8t2zJeihS1Y39f4KwiE/ZYk41VNKWasZ9LkKbIeA01rZHThGKBukIO
JZYzkvEHgJq0hZ3ngjhkG+xAKgNJ9jbCPZBqWCUQVtyfc+/qgqremRfInbpwl9Nw
XUN+SmldU4Qy0r8Jj1Ly37UU6n2PTbNJKGVpCLZsBxLcZwAvYveWceus3KziY1iJ
0Bu7SGB2Yftq8Bz+RZEdcnmSyiu97eYjRt0osxSLzu7AL+E5A8D0YfY87OonxM6J
WjANdjWGq5pG9Gua2YULiEIceypo1Q2+Iv3iyUSoMxi2xh0QjN6BUckJELeJTn1c
B+kItNY2pQFlBaq3SUEqPuSN0y3J+Ewiqz52/wfm9qfN4JXLJaSB3f5lXrzuV3V3
xS9qEz8eb+xq/izQhE8X5ykUIYx2u23e0htLRIdZjnl9zPyRYTjXKofegp2+r+n6
dC6Xt1TWuHKahQZHOrsRK6YijmyzN5N9lMHYRnYDo2tLWu6pdz4MnMH3vMmbfFy9
Kv0M5p2/d+dF5pwzdOylVfaqZbEq+hlV2vZwC+XeK8E3n62jUOnxXhn1KcAbIOlZ
x65vkbeNpq8x9Vg5HVx7m17A7/vvimEGxFLfgAd4+vESsilzwcYO9tB9K7kAQH54
FQvvnCdtGLGBE0PQF5WP+apGL09hqzZYOfbbQ/zYdDcunH7f9R+WCSBlUcbosVcP
sxO9ZTUSUKOuAJEe9vhrO+wSzbagJyAKrzkPvzOjq6TMF1sruR7tSpbk2UX0DbAm
qqPR5H/Q0V7Kxd651GSatxT/1UaNUFfDxgduC05KubcfGzNY+LcTsg6O1wRSHVL8
LUsyOWMkqlkxCcvx0sXx+EYBZsjsIOWHc446DGJZylp/BCR9/aVpfUDfQY4Ju8l4
k/IhMqwXJEPfFZY/bxL6GVK8fkqb306BGkOrON2fwrAV+ncKtv0Go4hKAVGrV2rZ
3f/C1EmB82yVzxVcqPJR323g+XELtjaWJrEjhBZOzhdrogjMHLjYRmQBR4Dmsym2
/YttP+8QBnu3XpGWzJJwnIVRJrKR1oSuUdYitpkh2Lp610gr5dMKimtom43Of8r/
6mYVMcW7Shon+QxXT6NJ17b2Jlc2n5acZVi7SeoaGclCUgIwMuLfLUc216KwIlpy
qac93yz2w8ZWSjZW9qCxicr1aDkq4xhHrEJvanzXBvGJhr+rYQ6Tb2nh0lPY47/c
Ev+NPTOKbNYEjHa2+v3RPjkdYEZUiFTJSWKca9tU64IqV05s+03PQNob2CaSyqz6
hJDDjANFvgkqidP7maMCN9Z5/NDBAiHBAZu8xNujoRKwY8PUvlLkpcsIW2UtI44P
yschlLcXs5BFH/W5RhSqsvlI/hkfz2psybsdonXaNkcMucluXfHUDFI1Vk6+f4SQ
OVsEfWHEZnrm21df28+34RXcKrsxUYXvulavsYK8iB2CYFEJuHiYSalwkgndQwI9
6QsljtNUmT1pO6C7c/g2H5ZC2S+dn8oSuag3gu8PzQvQtFvzAp7COEoJ3ySKWAyL
vse41DdPR4jphtV8lHWkNswNr3IcJAabU+5XO0AMVE3ONiWGB4NUsOq+XV0ME2W6
KXIkfikC5jINXhWmS6Enuif1H5/bHyyViDP58qFHFAcJ0lfz+JpH1pWrthj/wcOT
V6AcEYrqm/Uf7XPeieWXsuCDQEIvqK2F/Jy8/sRXfLxmqqkXsmqxaiMFl8YQ5FpB
I0Rq0OyVraNPz3UAZlyWknmc5qNBCV79u1kfFAlxdwwkK6NrJKVMdYwETQd6W/wD
ZzAFPMlkPBO2yQUQgXacR4laYX2uN3R9j3VBHxh0fkDngWIHamtKTURfVS8PvzFY
w/L/sNrpCSzp2v/5sqEiuBeThKuesTPDH4Vs1jV5FC1UudHuYXrWln71DvxfIwCA
hBHQ32m33AjVsCKh6ErvLQhZGv3+F4+670zzSMTrlfSpjLR8aNqqKmSXwQAjaJVF
dBzoiEneNmjoKi/XfmT8zbDAIKGDUkyZWIrxTCqr8Zpz0YcSV3ZMqEpL+/q0ahWb
LcFZJ1WXuHv3AG+OjHqDbG53/VuCNhIbYhkNffFZyAszBbnFxYNgeEiNAal49h1L
c7stzlXNIYr8B12ZqJCpVGJRaUwAYWXLxREwhI9pu9pBmJxnJvWKNe+q04MNxLka
fcVpePDKbNcvpSVLnXCqRKDslaKl4/6twPe2Kz0pJOoO3BlQP8fbRETz1OrbBG0q
we3dBeps3zIU8xRKT5tPStYNnRE8SV2KlbzVj0lkliRfPZvntgT+v3I6Ag16Mh7h
HnJckgr6nm0fP7NFkZIh2pVvgwP0/a2mQUmsU44hs66fY12QtbV9fjAIqgE0lIx/
A6anKqMu3bLhrbOZMAVGzylwgmOMomXuiRIAQMP8e93tve2FHT5sfx2VJ+O4JpnS
oNKv/sJPPJkdXn1qpv1AK1+01jO9I4/s5VXLRj8NoIKeeNg5xJfjphqh3NgdMq2u
nGnBFFA61vuPIBOzl33ees2IE4BjLfCtTk7P7gOjwPiM/mNR0+XBLFvoEmrajD3F
0XKEsa6TA7pR15Zvb1gHmBTztbr8Hr8mNu3mo9OcGPzT6Zu2gvKyNlV5wuIVyHol
3ycd9rIZTvCz1rxM6lHC3eS/JEr/iEbnjpZuaun4956gXOISvf575x2gxUDP+6l/
yB5Rrdwe4OZ82EEbIvWgb8kmzWdiGSYAA3hari05yYjfbfUHZtrf+gE+K+k8Lct6
QHVAF+hVq9MmxvsQrv1EvWB72TSIuvoNlpe1IYNFkaBQ6fi8pR/Ylc+jcl3obGJ8
hF8fqSLbvNnl7OrNRqzjoWlscnMMMW9bWwaUVnW9MkEIPgRmwuDMlQ1V2Ovy6L9M
pM1lV6WYWAfr9QO9SxAsyq408eUs2EcrvHEz/VAMIxPo2MTaFFKCkVlyYyKYzRpR
LxYnR4iBaSLExxDgTz+zcwO0R96VjqYOcRFwJFKLW+fb1AcPnH0itH8s0sSKaX0Q
B7BYPJLaQ3iO3SJlHl+dz+CWxpe4YEugNDomLu7F8LOvnf5cRBcOdmEooJB41U/8
DO8Vib22Ve5Vx/Gr/IVIMfXjfG0gQWo9iOU/yzXaJBWH/l5ooMZbo/iaqICTEMDY
+qQSesHXItE9Mqcp85H4wYC4BqotEHrmixd8ca3YgGrM/a3bHwVBJOGwssLCZ7wP
MHdHwW1LRsxlhwn35rRxpjst11QoSvvI7eLzjQhh4so06o7J7wgIQiYAkNXDmREm
TRWAa/LmS2ClXFp2ProW5d3oK+VHiUNH+Ie/4A2FYnHq8cicJwfIN0Gfc0Y75zrv
83EnDQ6OoB8HfOg0Khpq2U1jwrvgNcwsv3DmPZjRv4CgsoP7STHOfxtTurXTffvZ
PyfRaGDO/41ErwYx+/L2mMYOyPz74i8lMt1QC6TsiGaPvazMFCBI0BviS3VPEoEh
JgX1HyhfZ/8zrLcUDzZ1QKbIRY3WVcte1ZJ5c5TBG6wGcu/XjmswGZKj2q8Lyavu
RUOMOOPjDsMNeydT3GCoxNVL4+TVnRjf7kXMw64g5EBPhzQSKEwDqwzI73tnRxD9
FAzla0TvUd/Zs6BsIXUtbeoQQGoYkfpFjP6ZQCmpHFQfZBcwdzJV7R58KzIQaqkL
YgxCM3ZMJiaPPW3e1s5cU/z0lWedB8VLr9TkQPrwW0DinQon0fKTnAeLdnDynGaC
TslhSg8Vk3l8jkr4Sch53B8aLsETUv3Co/Wz1jmRJAcgLDW8UNo2dZImL4qi0C5M
m3dO57sqN546ae8eiOh4W9wLjTRfC3Bn3WVcPB+8w1P8jlmEXArI2UdPZjd8HQ29
e3pl4XEUhZhxGTVxI76YMAqXvG9jfQt2EOcY+B6NR6LdE230O7PXXVZQiRETF5vF
DDT0/njl6FFA+/JMplz6asjURLRIl/93+tVbSWbC06l74ctX4KB8dwfcouhWbk9L
zbsxGY+5O2PXeebyfJTwefcJyDS0P8soOnAz62zOsZi5EGG8K2Fi0MIbJM2eVaHk
vd/C7yECpctS5t6EZLMUdIWmFjfwFSGMrhN0WFR57Q6hG/XphBnrIXD74QZVdehe
fNSUdDbktdL3hHWVv9VuA8CtqlaiQlRFkRf402U1PGvjPXzaWfUI1E38VmyMiDwM
8n1Oj0mdz62wzZkYWRxA7oRwH6EkP3Cl4J2iUf7bqRu/IfsjAtILV6kuZfu0+PPZ
MIOeW+Nokj8l8Ds7cnykntArQtus98JRy+8tmOZtL4NfzurV1v1VggPEPkYZkqU4
qMApWsxIQCP72fOBVn33lzTHsDItUZT7KbJ+f00GZLlFCJV0vH9SUCBlx1xp9Wt3
XoW4NHnbe1syMxf7PrvwD+fUD7A/GS994mDAg4zh85ZYzsX1zczxTkp2RR05dvWz
QbbO8NQTebGI49C9Z9P5hL51w6dp/vEgSxdzvzM9b1NsVAbo6K+E9UnCADVmQHuY
1GJL78PdQU+zX1snul8mEPIBDWoBcsk/5/B4c5kz9ZvbduBjMAfHyehxHbaXkMut
thIONqvFMGREUnlyzs3UofJfTZl13+oyzhJJsmzGyFXw7SNx45RCSwG3MFkiZlOh
oJh/LkTsOFRk4aC2IiWkX1430JjLs48xLkEMrejH/Ee36DIKDO4PoQSMBFLI5BYA
VYkRXOX8sMjTdI5nY4Z0XPJPi/T9a/KNnZ8N0OLh7ztbv7rl4WOZ0N5Er5cAAmTc
0KqiTicCNhtOf1vFUHTIw2r8EObf8nCwL3Kpot73yHLlMvUrTVlG+q2wOPA7YHZu
x8Wtr8vtDWDz5HqN858RsLJ6oZg2Ucy7d26ctK6h/XBMy+epzcmrXXbs7T0GuS9E
Q076Y/57arNj890yM10H2ItZeYa3IczUzEovMAVRNUwZFDrJu0oBR6zkwqulAQPi
10s6vEUuxhgo3lSv5zpbpyqQ4s/MKIoDk90NxdXAmQcerz0m76ZIbYXs39Or6vqT
0QWS0x0uEPTxMh8GnN8QN/dIQQbkoepbqNpft6qCjhBr8D2JsoxImy6FQjIyCzEx
/SdyGoVyeKsgdCiqqUx9SG/MUiJT0BJR0fO4awRmkO6PzunzWk6kkqAgxSKXmSRD
wMTBy+n/X7jJndiQmPq+Ykx/KlrpFE4RyDGcGELGtL6Wbfnisb/e98+uDvYiWXzW
j1YQAwVejmBGHTf/x0HBNs5Rv/xuG+lWZ9ydtFkfqGbRYX00zawQ12u1SXr5Xlfv
nMSnUe7HRDvW9C3HzUq2bUR4VmOMnSjZ99SN7Yl2ssEo4kDp1Bmo/72uOKymFdaP
QUmU5NIgjYLG9sdXsfm8I/kVOIF6Svy/ndyYwax7llV12XIS2wiUg0OMC9cZzkHs
GIeifrdbwHWXZb6BkfBz402l9jc3wEV/K3AMiSb+LnVU/i6+BQd3flJsAdKc9k0G
pan7MqHDcdwJ88ovmc7a65mmKqiJCiSDhwUMQbUrywKuuiiqX4BRQZ94o02BF3x8
JIj020Rpc7XYHNp2vjM1N04cagmkQS7smPks17VWa/tRzai3hsSHNQyRcwx67y8Z
TzZhqYHrAvc2owzgGG3HjlI1O74XRrndFgG8oC9H63l5Jgb4g73yHAdmOP4634to
tKzaZxLReUddMX1AqR4k1r5XyQgvGB+IzPFk7702k0hW2XEbyFYuu8XBmVTrbT77
4Bn9yzlR3CvIAI8CPfawIY0+3xmcAbveL42Ut5+csSfsQ4lXnDOsj+a0LBNre1mZ
sdk11pY5+schje5ZN1u+HBJ2c7+/Vicu18pQPDYmvZcRAmKSu0+dS9YPyLkbU0fd
FDgjEUkbNW19gnxOS3JnrxL2j7ZIuBKc4Lz+aqCIwjCdQBdM/IgrDkmQ23vKi/nF
iBfo85hojKalrWelUw05VI+sAQbzyzA/DCaM2xI2blxMotwL3boPOL/pbefc5jEG
qmhTf1Fiq1QyY8ZzTIrNOe63sApB78oDhThanYUdTYn3uV6LRKH15nTzzDHYVXYA
vbH2LlejgG8+3o7QVzW49pO5e3cIqcGUTrph5eEuACy4LAlEtyH7Dug/5snjEevX
XzdvIFK1eD99X8yXdJSt8YRXu8viZDUZZyZpoud7wv0RF51nabvSQbRcMEep0L76
Nv4lZx+P3hPHzWichE8oQXINAoT69Vm2GbEXaonxo5OTxSA6ZnOv+qAj04FDU8a1
+lEA8+XTBp+WOGYh6q3Pq/sIMc1v47dXsUoPSFhgE+avu+wu3fJhNOudcJoW88Of
OGeOty9yxA43lyDkEQ1xBVz64F8xzRhwFMe+LeEEiCZ/HSyQH1P2CaTWG22ETXRj
5TNjOrYcAkNmDPJ1x3Bcq6IRBuJgM+ibznXgbjnwQFbTIV+RgdVs1zDdKTzVNPzp
X/Yubhozh437kYE4QVW0c8NzddbI75Z/hTwR2/b3DTpOF1581TanZqva2AcDo8Mw
fjsbeY/BWMVUebhGdQNbV7sQhs0X76jutTcFP8BwA1za4fg4MuqVD5vuODusu1Ix
t3t3T0XriT3aep3KyfbmkqFEB0mZttVMeOh1r0LKyId+FHxV24qVyoOA/qBAsC0J
zThQzNjrIkxJxpVtegdaY4lWRHNCs1iAM1gBUFtvJVDkuk81gH31/dkKSrQiRYx/
gYfKbhSHL6RS83J1gdx7nqCu7riRsMUCfeHolNQLiKVujWO9C+I0EhOWfYjlYuBs
dgWNL2j+cnPO1wNXHe1dckA5SdhjkWuAe7A7W4MYERlaGKD4jgluHriHmXrVTHhV
HjBirkiUOItU4vWZbFeeA6lgBLtxDXi2vcGJIV3VouOek6JKtoRbdy9FyqgxqFjD
YL4yHcn2wFNm0ANWj53b6j/k1QJbh8vtby7wJXlFMg4GZ9yRfPjHPUlHrC4/y8Hy
YlcxCo7UvfCQ7vFNl5fSf1FcW7C9w4VLGH53r3987MaISHuwstvr5J47OFu310CR
RjucyfQIIEDmHIAjfSlbKxZxwiPf4gbgZPXtD/kabtlXx1qCU4y5PA4Tjj2F066J
TQe0bCeqMy3fEsgPYtNV9N7BaRtig1cwgauSF8fJn4gIS+vy5L6pBVOimbOFjSfq
OAgxwTHeRLrFJAAgGmbAMOIY2DnY3ysPexoiuxCOBTcJYaPUQdNCadTP+lH8JHm+
SuE4YRQ7pPxcF8B4y5NNPS5baTKP+xm7kLdbR002ey6MTV3W4IhUD+sjqY9SH//N
UwQzASxMHIjdRlTx1Oeu7eUmq81ymY/GNV082xINdov3q4nwoAk+DNw+eL7Stndh
ChXGKSPcH1jZzb1QMYQtK0NpmQoKxTs2L5x96qL+XwdrkcQWF008xa2VE2trQ2ud
ssxAPansGR1c2LHqk3n9wNDmWdRbaE8EVcjnY17w3paoZ8PBNp6mIRexkDxZmahP
oH7Wsycza5sYHZ+gv/PlrjilxiwSES+FeEmdi8CqnsaT3VIqFqWdIlokxUzLnLRk
jAfS8qHEwvKZZJFSZQ7zrPNyhdzGpX8Z9NDLoD+GF9ogCH/a0uljPf2oxTVSJ2oF
easgVCZjq51xLsxfGnAM5TEggjF0R3PhUhlkcKwJfdysM/zfCg6rI94tqTm/dPTe
xDCv+15i0NzO3HvViZKslOB9zN45fNOivuKLERJ/RklsR5NpeT05r5RLCCMDDO+x
eC9Zdmyj3WGQif4qcPiKXBSSZzbrAtEwtr8DKthW7N3DhrJIZ+DRiZeIhm8l2Q5q
1ILFaxC4NQ3lrkg5B6AUTNlQ7mScpcOzLpV64z+h1AVw4+Ov01ldzWWj2I5MJcpB
mKy/TI8rn0OSvwps1zUrsdzd5C65ACIAj2PaQiYacOqKfJ6vYtWm2qufDsN47ycc
JzutmNHiRNthCC6iRRQpmvVP4PEsBdcwg+Nh3dIMia8e3ncDIP8z20uPeQPBFk2+
iOug67B7cxxGrVQXOAKTdRmPYORks32dQojv1P2UlPjKmapnrdEe3u+EH+r2+1tY
7WtISM2RUGu1Cxbuw4VdkebqU/eBqRmYCKEE5r1vkTK90XV7jE7BW0mG38mqGMEf
fdA1u6MFplntbODB0z+bsf5lskhuVTAJ59f1fQH0lstJPUpQrbQDPpFI6UT3kzbJ
mFZdhS8X3dZIf+w4cZqIoewt0XnzMotuzvIwgm2YZXw7m5A4S2mufmi95UlA1y4q
RCoYaqtz2FM+8Uxh+Mjq4sdp5NQJMf7PcC95Toqu/fFhGxmzWp3NITb4zioO3KjY
PeQZD8RzzwNjRAx/bugmmRexgw59rb7kbd0BIaru6ZBgNjrc80lVBmj4CNXCfUfo
b6QY9R/4LvFvdZJrZEZzuSNlN3Awxgnjjor6pdJwC0R8m8fyZenViQxRnIr3Edkw
fDyVXy99WNO9aDNTMs1TAbnrtsNSIAkM0UA+Fd8H3r+GMDeP0yvlQjGdaZXeS//N
/O8yplOMNzbKCrIX77VEAfwsX/ClSIk64UKsVZWdNGO51KQJGH1Q019E813Y5z3R
cpF2XN/LYETFB+Op9oqXkTccRCGNc7qvBncidDvWyMnIA0rgd+QM5UIdtC4MQKVe
7lS+YOnTsxu9bKuQEfCfyEAq4scpX0MBo1SM97wiGa+qACbFe0ss5lAu/AIUh0Si
wKVob2x2YPFMyDFeE3zCUDOEjjHSRszopBTsg+pcWI0rLGV+4rTHb+QPA0DVPUtF
nD7Z1it67zJEV5Bvg7XeeqIJicEgpfmRYWx3+fYnkocdcmyWIlJjRJNSUOiu1zll
K6VltVa4IBbSsCttV8UgIYuOqRoa1cSq/KoHvUWJ/iPW+cfKnkQHGG8oRYgXfCb5
/GE6UqVe1RjrKIAJRAJIPQCnYbXlZyR1X5OhxCiI3LPBttewYWJmmSDey1meQ8Cq
9zpUi9RbCuiFLPtWsS48Fxdpzb2yY0u+PjilepH8qPkPQjh8KK1vpC0K9FBqIlbQ
ZFT/aQzQIm6WXxwpwcpVVMJS9D89xHdGg9gBYAaofaR3qEkMuL6QnYvAOk75ENLd
lsm8NakxsPk9WFat5BC5OjFJG/9czKN0Iuqke+slxLgqj0fexckvczfoB1yXnqtr
DwRcJUNrBI3GX81UYNSB26p893H3UeHtaaARRzp6oLDQPn4R0ePN28guYeVT5A8u
G/I1cg1h9SaUexnS8Q1bAmvq08JpiMb8GvSN0l+VnlOYJ92fSuwxEN2IFY+arImI
mAzb623rzHcgk6FcsgfS+l02DR+vPVoOXXXqHZqgy8ISmR29Mth+aNekAQJgsxp0
4ew3VTvTBxXGyIWBbXEzGrOkPZQEvHFGQCBu9ywl6TICSwpeoHKUQBtMBPRpnU/f
ADNqrO3mPXTDdHKyTXEs1z/g13fEEyc8I+i5AyImlNdRYr+KuVn8Dzrh6uFYpt2d
QzhTHF20/9Rp6E/A2rsbFNTddXpOxk0msH2CWfvf/SvEiu77Npgvf3kskbQ1Hdt5
JsBPRCIC5z6GEcMD7PXrGCYO7ip2GmSd3otNQJvrX0xWTslPj/0UZluZk7TdMrlW
4p5PnuLjNdeKyzahTpPZOQLuDOdVo/wH4axSFg2KDM/dm/V2XEV/q2KgVyeTWRwT
s2Rh5t+vgaJSQp2B5uZL1ktj//Pwz/nx93Sb9MEZiFHh9FQnqWW6pYtnPUVOTVc0
cJxeoVLGpIJpMD/7cecnfWRj4wcZUqQEdx4UAwRt5OdOtppvYK0uy5vOf093Z/dl
mh1E53JXa/IkhB9FFiacYhPYEPFqtM/RdtG3xYcrvgbfZ1rXV5yHI0HbpiCyBY1y
TQ68mGralyU6vtkLyd6pLgIPfqbvElO4cQoCSSjHclEtVp+OrHxYOEEAu9UroLml
Z/uhNkBpEEi3rMXGcvyTrYqy2m8GXqeYn3rbLd4o+bx12NvFJJbKgzaOob7szNvk
NwbWANqUBwxSNM1vzBMEdNb6BmJNV8hGzNE+dN2paCU086u/IEyPt/EDfTn1mlUj
0fNrUqt/twD7sI3/mRWjAu/au6eh+Unv9Z8JiJnstP6SZH7LMAyWNa3J+wl6gnMU
+wCoBlC2sXZ7C98HULFG81nhO90qqH4GLPllMXCP94j8B5Ek0ZFzdXbf3msnqDcy
OEBh+aqrUGt+q+qMlwi8iJxhTA7Mogp82CT3H9KmJM0VzpGGTRx6ubx9Er2bQ20X
A52y/WuIRaZMGFE1EYvN2qoAtsEBcVblj1HjBVCNE/HeoVAr7RW89A5klSqcGZbh
wxFiLZZLzIF8Ode4Xo2nDAJCIeBGMcXzyKqIuaZwOFLirzascS7tm+NwE9i0Q+L8
DffZqBkfFOa61ysynWHUxz3vU4qeehAWHxfHMGcXlmj8zbEw8dkx69h1UeeCH9Hf
zos+uggtZ5aPfsw7GR5P+A3HVL7uqN+sLmotY9fKi3dYyre4ETC/ffsCyqJF7Ise
8XzwCKsV4xkEGU2xmGsRQRTiSIoDhSFVyZCEQ97nx83ovi3eo6Wtkz0/jeLqBj1A
BQoi4OxIkr6OTIfCAMLMumlRPsE9eccddrDTPAF61LoslhXddfbyZvCUvBltTQSx
bwLtrUXKbTEZ+UJ9elZckZFJwHbqS+vjD5e21/XhbBDw+G0Hsn7lTxlml+BQvQ2z
ilXPRQWy+mDJJzh3+8Y/JLjhk2J7FtW+pSmFD8TpbI3xYmd+MuZS3ULu6nz4DP1j
oqwR10jGHC8ijN8QRlJFvyYZGJgP0nOCBAjyZ2vpl+Y2HS9HytJrPELRO06s19G7
tryZ+MymMNlKqPjhqj3YWNRXUPZGBTlNNGlqyVJ/r1hkXOxKM0EmcUjTmmedOYer
OY6ryRgFP0ZIZcJJ6K2goW6oQilAHUBG8S0q4aKzrol3l2LoouQox3JVyVuLEo/s
dLLZUuM34h6E9npC8FRyPZ9IrAY76S1aSW5+SOeKo2VNsWVgaJ8+99kaJLhtGnUZ
tLmTzXh0pEhthV/bcESUE4jvUVJeJ0fSXKkr9+rc6Wb3fHa2eguOSkYDjicpgtEH
rhH/s0bdHiuetewTQDOYWSaut6m12vn4I6Z9BnoJ4/bo8kZK3uPhkOCeDqpaakbI
YOXQqNFOCK46jt2S022glJ0lEbEtS0opGAAmg1Cq4jYzOzzZVkutD0InV18gCUbu
0CUkqKsQb35Hoba7Nn6j9ayqii6To705Ko0JbHY0gtKPkDsAWk4qRuwBbiHYTY9r
tmKA2Mvn5jfKuC5vSUODTmIEv9bM7O7f2lif1uWVSXkGgjiJpwwjB4OXOn0Y46JY
15gvuQ5SnfA/vTdnpNNjDc39rQFgJBgUz6K4/KMt8OXxh6vZBMROVn5OtJ1c4K3l
cQZ3WKePA0TNhLu7WZgIozW4BGLvCpOSPHQcMPrMzJ+GBlz1yOCcovgt/W2VnZWh
cR4mEmR6fcBp6qg3/5a0OzhJgybG4N8L3WPdZAC1WPAbatyqnzux0RFLFfAdmuIf
dKI+HVMZzPvF8WZCvbTouGgmjHNIJR59cIzWCspuzHsvYVtzebhQlw+bNeNz9v5d
O7ew1ZPfaIFu0m6d21EfI3C1Bzy1ik7blqBqhoTXoeaxgN+ZEV8aT9uqXjjzVhmQ
HE/W/zUGLnymSksbjR5vK32VFQjJ/f7vTe6ZBjsXrIBWFVU5JE+K3+QnkZ6RSfTz
YeumFry9k65XgBT5XkUcbw==
`pragma protect end_protected
