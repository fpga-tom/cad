// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
J7ZARniRorkjgyzhSlfproHf0YLttUWWadr0p4weZmqK4P+2RMJmGJlTMLTyQTMp
YEKKLH0h6Cd4TYQ5HuVqGnrVhObYK1ry1HNcEhNJMM8zrKlA1CcYBH7eLiElfN60
DKmw/usbho9HV2Y7OCbs9Ncr6AgKJtOy1H4Fj4zpqro=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6944)
vwWSLZHi256qfOpIN4eM/dAa5x1FkqLteXl1/6QoxCyx8KRMSwaIQTSWNL6xB3IF
bduQllA+ocneJYqTPeWPuZsay6ThKjg0dLBr1Bq0UEbjwxKA5vCr6jvUXd534FC1
b4AiwWyHIb/fRXmYbhztWOJf+97r6tjOD9pXHierJtne6mffXaAUfBzj0uKoXA5o
TzT14KnDt0KX0g5wZsZI/1xi43e48zQq9kkJ46Cctdrsvn7tLsIzIP6eQuk7FVDC
sJ7KCWUwlve6X47JS3Zx+1AnLkEk47gdnl1H/TNh1lLObHeVMw5AwPjcZmMBjJl0
DY15IkalxiWEJXXivs2fd5gHqoXiiG4313lHFfEIOfqHJNGPjPWNNwiagWyq2LKc
J8t4UlWZQilr3OvaXHS3LGVR/tk5VYsL3Etg1mc4z0HTvL6wYPUujK6FcUiuHjcT
fD6VxQYACGZJw8mCdMpKJ7ZlXEDyPBrKsuQojYgO6aXq534eygYxqKT6HGKMuoQ/
oogdlnOy3qw2OzrxXU4/GkYEWkaE7F5xsaXu/bpXZ72zxNEYcgYHWjqM8ZW3gzFE
ez3h0469CmKmq0M+p6zDydnal3tEJJ6MhN5jckybrQlJRJqCBxFfN9tJSj+YpqC8
2YYHOuSmsTrOH4MBpN6ascXDZo0Io+2ZxpaMLBoIk/fXYXfwdPkzzeo0fyxZULBA
QRpIrdOWQOH7THbhgvjG1deno+FfaGcvk7pgD3LCgKHn2oLepDg7VWhaMn6N/Z2p
PHvoxiibCqSBD8/w0+Q2ROixurfP2bTd5kgcS0jIWM8FScDWU20tzXVUnPCCbaxN
9G/RG44HJOtvconjBbneKU5ktOaaLcBH224bp/mdvABwfxxYqmMhjOuxtAkJYy90
1rcUWxW4JLx2Eh1iWhTEtM0Hw0DI7oI6Jilv0/EGd6rAY3gqdLbuineW0l5ntuJI
chj7laDoU8jID0IktzOSY+Gpf59VM+Iq+LJcPQoZjiBmovBp6klYD6G6ZNAXE252
15mvMvW9sYqf1mGCWAczhkOA5tuEF+PtWLTHikHFwpbOIRky0IULvMyVeOaRwBsv
WUMIOrdFYR6B67GENKVQHa/MMuSZwzDe5ShY00vrPc+liZq5vu2OVGmL05gILFX3
u7w5Ksg3cxBdsnrXta83D68ccgn9gRuz9WLWiwrd911b2wpcbFPxtVkeYQHTkPFX
fsMgvXh3RthCsdjRyLXYHaTKdDcf/A8IK/8Y66ByjVD5pOMdxxtFavhIu+sSIqKz
VzKTaKjTZzgajX8GeOEmCpityGEc+51MDHcFfwwxwr4iTDyyvp/FHYsnCy4srZ4T
3MAamrJf498IurGnBaUQ8uksOxQMqVLA0lokY0lg1S38g4F16lVJOjtTpBQUFxfO
t0ZHEXBdM8qTb1xEvVpkTfHHJjRO5/Uo+qsWgmoNBP2foDTa41C5ndJbyTuoybah
dXvojfJAK3mg9WV3JywjaBKT08xuiW25Tpew809YNbeIhYSheWYwxNCVZN8MG3bh
MjAUb1fpVgrPky+vOrfjyuyhAkIgq8m/bvKNx+Ak89AVO5Scw4wQZZer2acYvTJH
DWu08gdDtGqCEc/1ADVxzi0fQW9fjBOk/Sh6NoduCWNG+ouB8UqQqi81xsVeXqw9
Q0C1HUF3JwMfZHLCtcMj4yyPWcv07D01x3VoDCoYCXUyZPZZS3uVih8OzcwTlNkz
h11yhmnX/zjyqmas/U7TMy+wHdxS7/AxP8SQPIR7Z6l8uWifpr16xA7IY1F8w9ij
hvW9yYXIGcvtx8FwzdsABYxcDAji0uZDATgs7kLL9q7Qmg9ZeQ/TlQnEuk9ivI7r
Hz4ZXpSw8nlQ8rH7LZd1pvcH5rAp/4J4GHobjYhWQehBymjjeUhv+gsAHhyZBpUa
dF8oL8gPzzOe3fRRDnPHuj+gagw+1EGSD7JNASLjRmkUprFV3H7m+4L0covE26bT
6oPlxjrnWOV7PGrI6VU6YSPVHCEN4BwRmYs7uT/DNgT28JEgWzY7n4WmLtC9dF5O
SxnijwyJ/R/NJaCYkIOV859CrmSDBOe8BIGxGjKltg/oT6G0Xp9AUzCBWiMwY/Bg
HydhaX7CpmgICuVZ3PirZmblBVqQMmwNe0UkPpYuTQF9ZS0oSfbtgtnpVpgGGcN9
L5ODlRek+Z5wSdgRXGg63kxFRNJ+HhgVlAbB+9o9Jq1n6NAt5QAnaajSiRqvM4Dl
syqcZYF47PibVsMc7ho3oZOD890wNlE24mFL3+ZZXqVZsL6AgfIsjA5A0/c9kITs
LZlqLj3DMRV7Dz3Y7IX2n2fnTS9PiLcOIUL9eWnk/JEHwd25mOxwH0iuVaLn1dkQ
na1lxhV4OuVQWHaZy8N7EFXDopXz5PXVqtjO3ZIARZiCedrvHzCoC6W2pIi+eezY
ZBj4/hL/649epWwbRneUavZh25wF3DjQj2uLgMp7QCj6C1PqVdfu/er+XjJvUbTg
aCb/Lmm0jPzG8f/z8uUMSHi81sywviptMHgfM0T5Z0lF/LYupvflb+fnwYn8IzE1
HiximnxydFUyxPz+b1x59cAKMAhSLkoq1O3RU7mxeUaI7asFBbFlzQgs0lzSkUBs
1cOp5Xllb596ts5KkjhFMCahb+YxnDGdEZluMv3elFQK90Mn4kA7l/t1K5Gdqjbn
YNSBayBRPMavQHX2vJVjChTVitU2+BQGFz8+v6mGjvWe2BUJvt4fXtKnHhGbFk5v
CaQ2QyXwHi/OOwr7U36LBUHgo7wBAwa0dIqiyLiQLFQinv8xtTOMtB39rcPlwD6u
usl7ogM9gNB82NJT79glJ7bCDwlSkDGs/tWbd2cfn08vyIoRtnfxzD6yC/r7ATgT
z0NM1bJUx1ul+D0198JgViOkAAb8b+CTpHhjhla1yUePjVKWYlPCjD4ynbbLwQ3H
9zFc1JvJdb0/KlYgl1pO7PvWcuV8oQYtwCYx/WZm1SuTSVQ12ae7rt3cIuPvbd2D
HsIkEM7sSJKecfne6eVZdyVbugzzWldsfteuZIXXvlunnIpjWvKKzBfBmRrjQVij
qG00zy5I1eA3Eo06+QEFFI342te8cGIY/85BrQ6HNaD2zr4GdO2HWKlARaZEwkho
ZmATWkSHnSJNjkCljfS5hjxOKkxF2c+D1E7Umjo35qoQyQdm7L/KIKaTo6r2bjfd
DFtdb5B/5nros/ognFCORb+mgK0TScJiZXN2Zu0MF7NbcEtK2AgGOssQptg/tnBY
hH2la0rB68rHnA7S6cQGo4E09KqK1dvlaJmrv6W49frW/wVqlvvFU9X6bGQl/vJ2
VCaYHmNu2MumLNYnG1HMuEDNQ22ma6yZXZxq8uD7uCkGH3gbD6dIY6gGxykac3vW
26FJ8t/b17VNcGqTXJjbV4/sqBR2xxtEZCkrHuRnybRqaKM0KCMIVZa4LP6Rjd9h
B6RTbDUijo7Nm1Ydvng41BNRg5DCeid2thH1eZHBC16e3uTGJuXO4S131fnkN/+K
nvMz3DEKeHlsPANCuy7IrPD7cViul1vGexg7sv8ujOBho8GlAcSct2Sdju4t2RzO
GQCsECrWQXFst+oTBMU5CLbkGFdUpLVhcoGqpG3tMu0OHr0dUDBCGxNKg5+fbmLE
g3ZuMaq41fpbg5QkijWbG86vpae4RB1Y+kS3cv/1Q0vJmFUBZXhcFgpt6O+N/rv7
J7U7w7XNTaSAR2KvnhWweVRWkmP5obUVhB57k8j5EqoYZkk76SuxgC/dMizgDnzH
6ri/xzX8A11LbjGM9wXCOXpU6Z0jo/vhp/0ovqF44DCBW731nIgoe/p914t2YNTd
Vx2Jz2jwoPIZnbkGEsMRPXe8WoajMUFiocUgLvaVQ04b1dGiir6S2463NFpxQgnQ
q00sH5DnRdQmA7lGsd/7+bhMiLdOuKGmRhgwZzPC8nzebKYFnKBkqBJcbxM6egnF
VljNlkOtXRZ8/McWrwlW6MlcUgk8dni6UTosBhsdEII1RajM2xI1WHFlnIXLxIdn
F4+BEDp7k3oZcMoFL2IN8sA97AYmCc6gRkhxEeQ4rdmTlPm5QUh/lCq153NrwZV+
4cOOtwEtVA0tR16KXWoy2+kUkCeOL/cVZtTPpjEmxQ0l4yiNNRRHY+0jX7pQ6oiL
dtUdQy7CIJ1E/phAh59Btiq1lDW3VL6CylwRPdTBnL07kmNzrKBoGI02se50qjW9
oo9PFwCkLWKivarbVc5XzxS7kbOcphJkMa5A/3NBH7034NDLrDE8SUFW/KjXh4++
EY2094radJrvJWRWYs+LHMaMamLiT1ZGeMuIPBwDkNCx/ZWgx7ox/ynHdNiibu4c
x8KVUnVcgXW5KX/2XpSwXRDIcghk3f7A1yQnrFLIY67e+5d+4aB/GEX1KRW6M/c4
Ec/y7wPbxXNcVig/ZKArhYXiXAom1QiTkPdg5mfB72AUvQFHq1pmTpOVlMFWSnsy
amDDV+nx7gE8MqwrdcWL98jXiVhgxHjaDjKoDvUq1DEUcnhth92NpX+6dLyLoxZE
J3ldPj6m4K1Uve2WJaTQIcCyXzXp+0W8QjZ1LWsKF2ktJ/O9i5T+RXxfhwmvXFsL
UGu9QERZcjMLrURept3GXdg1L7eK3Aw6GA8vRB8zXHGYU8c3kwYEj1ePD0S1QwI2
bzUm8c9ccUawNQL+W9E19EtFJoE/eXk23yfnSP8oslmaiYA3PYt1z1F3HTMpgmaj
SzU/QPaQl4vwxS8RTCTk/28RU034+NeBP4ZaDo2qd+8mpJCcuweAwsnneEbGfupj
T20aezXfPtUWHHifGr8xLhGvpLXjU6ffpJO8CW+D8PNUYZBoUEjvZxj5rewIdiYu
aEehbkDG6Y0NhR+nf+lZfv3lPwbw19QuiRVS0BTWE1ZnGRUefZlNFD7hS2wH5lLM
KdY2mt/ToZLgVgdTYx8APTszsuSwbXVvrNKxDWBRhdpsEICP5m4miVETVzmoLDf3
pt+JM+V9zxJZC7IZUOGoAiG7ZzL+MvrAgrSBfY4goY+dgBPUtYYHHnAyssDIKB1o
BMJhjthpliI8QRDDgjRiy4u7XecWJ2+pcN5iLsIKjfamC2Rv5wUZV7LTmlXe/J3b
NwJqCpC900OeAdwq3i28xtKQHQsztzmjygSyzqDcto5KBz85Syq70FGSPO5Sj+ce
C/TQcZJf3ir03EuKjs5DVLcTVgs7oNhCOhpr/1OXtK+r3pt5pBoeE8mfS9gASKII
w5rQqON/urTdXLoVypKc1Vhehf04n5cA57UmIuqGtWcwMVUVXETILE0tOLvIvgz3
LAWWwKXVrgdp3D/xYSRXX/1SnI9BdLTZfV3gx26GYsFCl1iuSwG03nTlhZJDyibo
OkuwgHZYPXBknQ6zSqutojld8JE4Q5M6fEMVLlS2wK0FYVwGVK8U91PsKl28B3mw
ffxAYLVULOUBd2pCEjEJzLQUyb4Dp73GR0K/ElYQOJoj52IWp9XfzN/k0tLjqoyA
Cvt8QxlqBIqI4qbJHBs1cVVavAg0hr0cGXMhp5ZMO15pMyTsIMhldVl8YFkRQ21Z
eK17NQdv3XhUbHC+58/z1NDpPh8HKfmSk1X/p7rUmZwwnd5G50n8nsdV9UXrRP65
K+mZv/HZnxfLIT/Es3K7ZOst/qHmLDsAQ8DrvxGrwodEP/hUUUStJwWR/pXhFXmh
3koN7UQDyOgkWR/OStj/xT493TO1WjXCRXLfmEj2KTsYn4pkAVoyqjoppf/zKEs8
STk0Trmrdw2/8BppS6tJTSbu4V0MjuD9v50cwRlkG5/YjCaEj7gE+fIFOko7WaHo
9/9/E0OjkEVGMxa1ESSC8XfRWky/XltvXxB3XMUiyMQOd/usgQ2GR12iQFh9yiQQ
Xk5JacgefjMXu9aNCgNLHfyVOpQseKA4TdYZRHS397DfbBS35734neQuq8CjwVzb
OVko7ohGh/6/jDNUwfou4pjXHHRkZAEcnI33ChEP7lT75aBMvHnurVklWqLNeeGH
aX+MnWKIsD0zIug7+ht27gcC2+3jPx43YEwRqocVLe42gkUVjBX2Sn0O23hlukSW
98201NW22H4zl0LNwBkw7hlYNWKYp2ccRz8p072y6ICZo9GMSk7SDgdIG5ZxqkgA
6veXIlW6fJ/Ttp+X0WGRJOPMHkbcC5JHoaZARs1nlbUSDz4HhkntN3gdDT7NW8b7
RjZu/DjJ61zxxbfcOVVFrXQrItEwy2s+z16Y3Y8c83WKdtCYPTC+xaRhauj+qoBX
L2W4xp7/OIXSDS144y/WdV9msaTe1/iQp526juimsNP3uHN0xv0CIt1qzdXGhv5r
32pKVPtwqnrWg0VkLCCCwQpJgIwoJJXr1zQTbfYUWn4lDhRiGoiWAYWUAT+GUIRi
SwuwZhFFgxu5fblKiaslsMxRQdTEvyKjS9HzFdrd9HEgn9SLK8q5O98+haJHbL/a
ARYUdabczop4w8o5NeCpNuMI8rw+9Ys6H3xApfGEEOX/5VMox9x0P5Q/+/cb/r/L
nFWUM2ub+bYAfwjq8QRbvXEDum5NJ9zWO+zrQVr+r4izBLQW+ejxqLr3lP5Df/15
tmSvu5iEL/gK3lFVibiztAFQ7VmJOeJkfOskPHj8TcGUVEfz/GPz/asIrmycvUtJ
cBtlFApAWthkrVr43g/54uZdDBTr1MZRFQCiCAOVLx7Q5OCx0UdEjLwXvYiG+Ax7
JXdh8A6fd3sipBnwu+SVkDeEuXtsQU+1QcSajBKen8loSlIX2bfLcTrdUC1RBCv+
lkpEV+GRZ1JBq3GVqpE0RYI0rCc2zih/KnKhVAe4bGeXjt0HJcUoa5At9fXjQUZ/
IqQemlLtgFzQd+FMyZdsuC+nGp7avuimTNHZXiZFCHXMAUe+mlaWc35j2HWPDScK
j0k8BceRmH6zSDbGXmBxNmT+ysiI5ypC6i19fw6I1LPlgqTspsL6WB6c18Hc83vE
MudTFzPlgqZMwVPFhDH+eJiPyd1E7B0hbiiG+xxJVRO1R98HcefwcSey9lbkIPzD
HiunEDNOlwFmQpBV0RPjlDWxOpZzz40v3a7/+yu7tNup8iXE/WFBrs1twvM3dA6c
hQMpFhNKNUIMP6Y+fKxzY2aU+KtmABZOLp6I+dCBjOCESeXyOE7GDvqz2dwKfxW0
4ZrTFflgkxMYZDaFWRJMOxfhqQpYMp+Y1lUs/S8KwBGC2QEWxpliJ41QsfBplAia
IzP8t+mYnpvExMD37q3n6O++EbUhHUeqRw//xCrLJhRh7tLq9CmD3zHUeXzrXQ3u
MUeaikr6uqMnDoDSF+ZGDiSxepepfJ90doE/skRl+3xtJir/Hw502oQREq+6OZjB
G8n6cWMqbmZAg/xbaTNk+QU7pnSraC4PvryNoYcW84U0xZd0Cn7SyMMWlKe2S0FE
PLIRTR83SHKh33iufBPD33kxovVa2E+RAXahImv5IecSdwroCZlcZpWlHfQJ3pnH
d5qG2Ee9PpHuYj6L10B2NJZpc4GzfcOTSj5bwogVdd1iis+PY9vbgPI0XnQQi5PG
WJDDYnmAL/mvB/bAmQ6pVkyMOKlACODmRdSgo8yOXK2tTDKXDlwsB9KkOEjSnZRC
X6npbEm39sCu5rh1CezcCm3lFYNHrJjRggYGrkltvkbubJv1TS6vlriHwuclv+nD
L5AHiNvLeItaA1x81sOa5LG2vhdF6NnIh0CJs2EeEkVtTOyhRdAFRS/S9xFta4eS
3hpjoTo/N6xhTJOweh7kFjVHY5xbgq0SOmzUFS3vjXRjqq/hD9cJFri+t27m3sxT
tF4NRnuCK6o1+9PeY59hG15cBUCwYYul3/q+wqlIzN4+HC8/hMSRE9SSGN3eYwSS
rbY6V+9kXSks7S26+FA9G4cnBHFwHtWpTeXJY1JwC5opKXZr7MwaNvoQlA0STewj
5Yz9E316r/uPFjCz1hxZGSCXgTPgbxHUY11s0eHL+vFpXyPnsf0dcc8Hd+rUhj82
s9sT4DyNsOWpbORqarKwQE4idxp0ZGE0tEDlXilrygmuLd1dObDgVRYQ6RfibzU5
rflC/y1U2TNKzcLTZ/W8oklIOT6Oz2SMmXDvvk6CIid1YC9szQSe+9Y+u/3sI779
Mer/CFQcXQ2axIDT1MVXm1TiO/KRyqEATIPOqSZq0739b390YGB09uU7TLuSiIi0
hw8efAN1sgYtZY5XmSZubXTjfAi5T8Z8m1wXJGCKf+u7FcZdd7nTfsTLmGUBWIdD
4iZe09UU29TOH1ZBiegalC+MONqvgkDvkImRuyeBTLeU+G4ZN8E9jsI7gKsGd+bX
kn0WHLJ60UA1tWMqwyxd1XdQXg/lkiWuqm16hZ8PH/b3oBteu4Lg4MXaRz/0uvZG
AmVJpSkUsiRp3dBFbcOzbZimCCaJVpEuL5pOW/oC6uAVwYob+6sYT/RxhjzCNtJs
Lf7TNspnPrzpe+ZiYPvJH22lRIhJdWB7Crf6AEitErnsC08GXQgw/z+72tl/fMT8
j36jkYK5vQRcnIqLTli7OMFohiLQSPAHuMoVMPbTgypHNeuwanmPA8gTroKktq0Q
OPOH21QkroA3YNA97lL+Cb4fWVoxi5xEsZFaDQObdx7PN9HU4Z+K4Hw6fUfbVn3+
LUHOhyaDZc905Rur10yqVWOwWjP4IITsIEpcUtx1IvgnpWFwEORpyy26q7klrStz
Zl2bXfJiulD6dLqaBHlVZUhWBIJSrRLqcb0ddZfMJlg4yhJcUcmXBJOd2I9WurvS
LkUPSUNgpXhE2W8b9zUsAFb4l8gEfmq3e7qjGskhMNL+8mOa8fojxI399DYibCEp
LWnkHla7BGXm8uGZtNYdmTaqzQG4DFgdHWe8jNgcvKRupo7HFitajiPitnDDVM3/
rf1UeMp+3bp+INbt1bJlaRyWj8voj/I0aNIlyi+fRLk8YculXLjb+kDk+UMML5Gq
LvmLf+R6w4EQoegn6YWRO8HoVtzMZzJe6jE2ZX9+8Mc8uiK0dHQYTOJ9eCRnS87w
qyBB4xeT8y6lNuxTGLFujFy/LkqLKSqm3DCeqHL9GG5y16pi31YCNxCgnSjPJybt
FPHnEql3YLW+4FpIsbM8G62DSQvxQ6IH7dgBAnlOiHSeVKV78W1VVNbFgO5sSD0k
c62IkxMjym+I1zT5j76xRH6Kk+q5fGUv3Pdt0UZNko3LpsGYV3AvOvqPDUsz2B2v
nxzyL+2olDJ4B87UJBAsNDWRTgqy7ZQw1Xmsam6KNzg=
`pragma protect end_protected
