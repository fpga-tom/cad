// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:31 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EimhgYIsCGcbBGG3nvjCQRJE0Xu2eKYgrhC8DbzXzc4nLPiQqZnvdZoL9J+gawZC
SMhik1J5/UZVwd1VvA0ldQqk2qTFt9hv+FHNz8Q5L7eSZibHaVEDJWvlIyy8uUEe
HUEycwq52bQX/ffeN9QUTy9GKDprXEznMngFScYC2NE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
IIsIQe20Un8/sbPu2pTmq1Gx4RChnItSjedK5WI3a0q14MYg71Ekp5GPlwOI+L6e
uPYLo+ihQTBn/BWt8rXycjmKrPsNzLouNAF811u9gIZhct1XTCOirK6LTQW28p8T
S4rRBwHqMWCWq9e7WDA4xiIKrsfVeH12/MYuZ6B4K7E09JUMM53H/RxUQKv8ytmn
9Z0mD8SeVtPgRGpdgYLqktOGbkxJD0mFRX+8O8aNDR/P+x6r9u/eF7OVjvCxm/m9
Ubh7t3DgUqd/N2irYXRkCsrtfq4eEsrJQOaIkAvrgboCfYb7tbDUT5H8c7340UzF
fOt1GIQkhNGgmZExCtsDD7YQOjpwBsDcX2JFRpfDcNrVgvTJEpoLbTnDrjKK3VoK
3DRzjXdAU04qRzCt40ny+RVI8tx41GWwEfSJD127ZOLuXIzrHPtEj6xcGJ7Oru7B
8llBAL+sOambIYuk9pkNVflL3/8JvTo50xOmjxLgSNiXQepdMpXAHNHRTPeCO6bO
CYOUPQZvMjiNrZpSLRTZHTK+YyL4IkHy+C20qQKCy0Y0Jh203xCbQEau1VrEWtBZ
JGbmm+WUXOY5XFgBVN/yyRKgr0pNjRXb5BNVsxrlltyPolOT45fCLyMtIVQZXakz
NEQP+rX9Nq2U9V5V2B1uIfdN27K6K/vKveUDvzKo8MGBDzjj1DP37Q+KrTZTYCg0
NxauLThn+LrXuBuLc0DuG4bjgT6jHotVrF6G4YY6rnbQDDWFf9Ip8ZDsfHDuSlOt
BErY9fP2ZSIzb12VQyit9RZFTPhYXKtUjI5G+qCRTbkswr7R0qg8XMaqb4yjJOiE
+xa2trvwlE6guySJFVgELJqQMazlFybdl4vLdMFuwoBlOX16oAndpmB+ludRH5F9
NRyImfJjuRH7qvT8lnRK8sz1ND9hkDhTdBdwjrlKhSLif0WdP2sToks1M3p02nkg
nNlGSyxmGBOLuXiuKtmtiYE4LQNrw0Hozdciw7L06I8UsRuvEgVGAegyXVkN5q4Z
r+cUjKQi6bvzeeLYXHJ3Elm4QnTOI7xbTclfUalNJs1Qluw5HZpIDvZiquaZTZP1
lhMJmBSiBbuEgi7RKgdc+tfF6kLJlu8atvKMhAAQ/dAwPz1CmdKmcaevj/22G2F5
RV/SzAHM+YPFhVH3dvHBVP5NNxoFQMlh36llN8BS2DKdB+DRQVHH8XE6ah3FVKB0
qHERnxMRqeXKb4k9hNFkaY/AMTor+BdjdjzSNw8L+ntkLOD/wBBHfsGbquBYahto
/MNjyXjkRlhpPiKJwabYRfzr6t2nFWNB8Zx7LDshj3Q0krOyF/4B27Dd3Dhph6lT
VHbDgStc3t/dQp0LygTl/1leIK5rrWL7XtXAXJERYyrY2jI/UMjxcTGxdZ3rAp0/
1XjJz94oYTJA3+I5UhWazGHK54fvkYXEe2oJxYDeYr1+/cKEZROzz5l6dMyr4qMi
QjE6NL6XLZld49a6MWkdJfiTXMYd+tVs98W+ZGx+8dZ1Nyd/lX+UGyJrcJZXWR98
Y6n/juHMqJFfFWt+qvjwXCm8SEaZKPAlH2C2fD4u+xSFB1lkRo3XT804AC9fXmwi
y0oelqKDgx7o+P7Ey00i7WAVKgNEaQ6xwTJHccE4wDE7jv7eHpT/JnIWAi7Gg4I7
z8OClOImVUaN9An9g+aI5vYMoZ2BQ08GIdo9GnrXa51pkq65F6mGdcAH0SgtCr0Y
kaMwWoYX0uWluuzs0GRJzeIzVyzWca4Grp4a+lNsMtiy2n/0Xi8Jijk9mgvDDLex
0aFYU1YurmPXkYlkuDkMT+CpKL3c4kbhg4Ra9TlJ2LB7MFSXIo8s3lXgTmb79Lsi
WL/A/CEeon/bcSL4Yxnmpwp/7+VNpRhsY2BBfZiX4DMNAgZxOhqDCeTOzgiztGau
MnG6DV4WdxFS+r71QtfxTjnk2+zP5MP8RiIJuBqHVcbBEUIQV18U2MZc6WoqQ7uM
lG8+LKFOjlxsVJNLSPAgkMxOG53/vi1UHpLvjVxhvtILFcZH2cOfK3Wa7pgKNTDr
Y/1OZZeI0t5JUZvL37sPzqpqcPa5WqilOBbj7YeBvErgmY+hkLaKoZv5/yJYTVeZ
8ml2WiJ8q8ie4XCmljo99ITSe54xfOI4u02OSeEUpVv1hzF1Sc8ej+gCWCCGDlvr
Ej6tfYSQu3CaPXRSEOhyTQQFNIXSlD0P2kSBykHZV9MazXZ/06QYkDW21xM0qp5x
cdd5dgm8CsD4rR13gZCTuaWqeooEgUj/rTAZgGF263bUBbf/8xuIRKROJUIiGO7+
40EF6rGlKRcYZKXdDpIs6iTmPsNlzFlmHSkavMVY6nm22lWP6acbEekd4q0GgSQQ
c6h1+HtHTvX0HCnVDhG7zPzJRqsBVAAP4e229hoZCLr7J4pN8ZZIAhUk2a3pwAi6
7hnJ3t4R3eYSDjbCauis/B1282thdhjdw6ufamTID+CezJVNRqn3BtcO64B56bqk
6HhSlrb62R+VCcvaiygCUvcI+zfQPGnY92IDslckUfwONun2RCzqYhA2NXYcO8aw
VnlAHzF32IA8Guj5bdkapEfHfcAGFDWWan4t1LsGGhKSaeMbru7durNs9TZspKk8
10E3q+XjTiPWdHFk2JNTbyPvRrQPUU7X3jaS7X1bWJeK6V1OZnEapkFZp76DIdK0
LtYGMWXeiP49sFEjA42UPGB/CR83KSv0DDb2xJ/bleb1LqxIZkv8orr4rYvQ3jYz
YuQlQtNKVUIqzsuWnptpRMQjupmAMrjsIrhHnuSzSnt+Cdp5gKUfcr1xm4TEHBlJ
Jw/YIro08vFd/+2ioEUFNv/R71lqGnnhejyJISyibWCTafQzXIuSq+Zd/gYa3+bG
gdX+MfIRD1WmPhnBb2hAa3KnQTIvjVthXlEVBJjl+dTqf6usURzx5StGEJatsKo9
PnFwsiej6XzsXhnv22yGectDkDVOZoIexisjKfRLvTMI7H6kSxAqN6Zupm8EH7YM
Z2Gs4ivBy1UbTisnRlfYTrsFrMF/ROOOzL58FydUIHQgIbF7quD0mj5anuXgTE3P
K+sGjED7+rxl6qfa/Qt9uAvnnNtEB+ClnTK6K1qFFZcS4uUtAdhrauzsDq2wtQri
YNyCqub/AUb0am5kxxCtkPUxlEsLRdcyeegVgGhBi8EUctuMk7Kh5f77WOoxwklF
7TzRIhWujxBMA4tbJBhxoHLxN5IjUBrAhwi1flPN+anJ6HxA30itK3HdCEdm0x5E
0ztyc0vG8teC6PjZw5ZUSRiIbufwBfxC5PBBhqm0L8zVQ9GDHVlzZ3pSXXvETMlz
OFaGsFKj02pEqQVfEj1rGvbNb35MU+ypp92k5PhrZ3B/bHja9qj9BYt4mkRFdiZU
o6RsQ9kzpN3zEVbUNZZGeiSkYIcujl0G57QQRCifgiEw3/pLhXs6kPt2i+IEIr6a
ja7ZI0VCvlHQShDeQppOyE5Uezq3nb69Ww283gK8bYYD7LlP6QqC4xCIILD1AU/9
Zwh5KP7blvQBwtW8Af0GbO79oClF5nzjBEpAHxcRLDJYk4vyOjQN2kaJF4OVzYg9
vWI8T4sOD40yoN1B8z6Eut85/BWDyH9zaowfyi3xY9erc9i/BNdptQlZ59LjZAKF
4eghcGkeYskmJ/PGdmB2ylpsro/QjgqMr7KRJf5/9hNzJGrvRpElJ/XkeiisZwp4
BwxUguA07giQbnMP/F5GmThXPYiAEQCLBxlFysSrHR4TJ+7qTzmOgNJVJ2xoh6Kd
7VGVU5ki9fdrXk0XgYjIk3cxvFF1q9QJZOMRvASoyPq1ygMR4djaOQa4vTgsOYwc
PXYX/kRQziyxAPgzLR4bT/eWMzwV/M7AM2dJFE1MVYaQkI9vNGxxucEoh30Djy7w
26uxWjYe9u6OnOyTjZshY8uBmQJq09v/sWV/2tQ5OQBweJqf2UXX9v868Ae2xqIN
b8QwGwRG2eCPgDUvreUqiRK4xeYO/K3O9TAxCHOuIf+RkIEX/X38544fPtYVOx6c
m5G2Bexqnx27TdlaZnkoRyfBlOm8h2d5bh2/8rzHQTLjhd1jOHsylKelZ8O2qro5
y2K8lHI0Q9XxiMj6/BTrcP/BmFcFDSwEUpD2N06BtNgJ5rKWTk1LxHYVB7wX0OaM
+Ie5sfjv9qYwxmzdf0Ps3k8KVFbBHoavC3GC2S3x/oL0i3h94dozy4qTb6Ca/bYg
XulPCE0FZx75LawjhaDxN7oWOelxzFtbF1cnK3muIF5EnovHYx36L3uxE3afgY+L
shuewjtYOBnJb+lhNI11iu8mizbNw1j2GMk1f/3MnPgxf8HhUEjuDKSZPjWzKMsR
f2eTpVz7iKitPhcYn80ruxPMpAM+y4FJ9RkofCMbGJs+O56/b+A9dNfpdwmMq/cC
LGLuylyx7zo6S/UEku0dvvFiv8H6tABI+Eh3jBg427q9VFt7TY/SpGOK1gROVSh5
Pvbrdd5kSPztTnKHxc+oxGBfk4sN00VlZqJLwxWZX0vWNRlfNMvvvJLdzgY4/ngc
jEbJU0w93dwg0k2KhwM81QrX4qX3c02v+ZFc/htYrNvrQDeGHOlKRv7mxyw66zWU
lNyIgSDGShTsN6NzVI4L9s+1pa8bdVXKdi+D5mLhv7P9PjDykPnfl4Yvt2fDSEi9
GvqDTAvRvErUq887tvTEvcy/Ck+7BPX9YKHR1rrnH1fkodYFLovgkkIVjACLrWI2
179MZ3JsgiSS9vpVvgoh1Y8CH4RmNK6aXsO8wPIjaRGTvviaXTeRKi5iyOxhpSkU
cKDma0reom5ZasYwi/hNcFaE0IR5Dv7TyIbpxm6fpPrTFeH6GRk4PJvMyk/yfYIa
pacUwO0kQ1IA3I7mJM+XkV/mC7DsNPFi01kKoCIgzlt+RfMF85n1GgjsikRBYKtv
aYeYw1OtyzumqOXQ4a2ywg6tRPYv/4UBF/M7R7JYnMPSTDjyWGztYk6IK78nmE7t
LLN02OCBBGV4zCSVdlD//XL1aETGEz3X2TMum2vR1zxzew+Lr7/goW/dB1gdzwkQ
SL/N1lniLgavXpejzPX+IaqfAfzAHck+iGk4KWaLZiT6MBoNSdGUjd8L1ZKD8rq2
cQvtAfEmApwDXNMU7jyFbcSYttcH6iw4iM7jp222isdCMolB/ixSQn7fN4n1XuT9
HkwanYbP4Pji5C2f9ou+ZZWJPNcgGqR2pRSLLco8LDntZIibk9XDaZyejefM2PIA
bLlwvqoYdFyIxqBT7gskYXVch7MBz/eyY3JaPBltIMT1HKXALBBivwd7r/c3fEhg
bhlByp6OmKagJ9iZi4aIV20sFojRonby4UASIphR0IlnkDCtwqQ2kukpkEvPDX6+
7KSgvaN0EHtu4OX64a/mityBrE1mPoBafDMdrxccGAxFlxCPEHBsv+u6o3wQ+euK
jtEUgcPSo/awnWv9h2tMhVyL9s3fz6toxZ1sDZIDSpVJ66LrmuMkwg77N+0fuvOs
F9awKWwlqt+6yFF9p+ecADQE3gXvnAG4ETA4PYKWleqKjTDw2zOPb7pHzMEaeKaF
+NnZgYmUKwYTcyOGcXwjcoGRe0qSs++E1iGizchdzqYcjFVps0V9NW/QM1WdzPnS
itCOecCEfu9DPDl+0Vjo0DKQOHCvP1+ZF8/xxH8AwSBYRQfh1yXXiZ0BgquXMIv1
fF03oCzwxdUMaSu3R1jVZ1TIBtPhAmfQ1ahDszISJ0S5ppT5/n2u/EXcqbZWiteu
OPHs40uOgz1yNuhbdS9zzb6MVI091f0FSiNGyLpcHBsVQbdeT0+f6mnst/ioeAMA
bOpb+LoF6Og/POC6AwRdFjMTHPPZoQ1EC/Oxf4i3ZZki5CRc+AMyundXP8MP7o71
mKDu/4QdWl09Ak1b7y3nDqrGR66EdxlAaFoSXDG66Oxdrvh82zVX/iovvWw35zoU
vXf7Y3MAAiIq8KJegNnQQ+YENXPRy2W9EnxwRZxxO93kk6M5TG8Hd1yqr16/Nebw
faOB094F8MvA0DSFMjYOzaQFYci7MiFAydOUhJCfMSJrA1yc4ybnUC4PAqkBHs3b
eNB+gHXnweMVCENjuuthVIp4pdKLoHI9kNFvpmBA7lu3FcGbn0kFrW1klxKuUlTk
MhBa5+kEpSstHKthDI5bceq5BGod30OwD7yZKOvsLvyIsWim+6YLIcDMzgzvqqAU
hdMsbKvFV4pRIVahpq3hMm6W1zmVavnGlgvfkiBj4BejTHRIYoAo70tWLz8VKMLz
ZT/wmthjH8xJRpIPDMuu6DBpruBQNCslgeXHcVYxHjnBMr/voNzPtRa5Z5lQOFHa
5XLOUmYIv7chmDFPEM7ufH8Jom+2PFYnnkYfxxLibGrmz941q2R8cImwwIojbFPG
/Isd9Sx1L3kmFevKnZWAzURX5XGnQuMcTI5pxSd+iCHA+CPBf6Qo8Wj7fAclJbqk
OybXY3CePEG/oKEaP4ov9DaIVvCwRhVUW8sz5CtAYhANiihR0rqlKfkyqu47hZz3
ibFRKoiB9XWc+RgjXy+zDAVKkXZB7DHj8PC7VSSTURLOr85aBc0ibIvMcnxWhd0w
7vLZhSS4RZDR7A8g4MllQSxDLnpfbERU35MbLGXsckxj9fphE6DLEaa73wBDMGYi
0AdvRnsGu0+ghfgrd6B/tA7r5j4HMxEHvFdawSDQgo3cDbrSH0oNYLuvejg1Rr8I
JhOo/EjFhd/F7h6Qkmu3rzjs4HC2Roo9iOrvJROAZPR8ru3zj7LTubniuwyZhwEU
4zZmcqgCjLcIGENk3yvTY4TORC2YJnovxMzmB1e3pFinSrgZdAkTwQxX1eeBX4Vb
o9tc59dILtL5wm5GUhrNKTW7dW/RUY7P6B7smksdtsPDBMJE/x+NWQwayxg8dOGl
hjE8MHDSzb4EY8tRwlYmSa95rCVueWPS4EnS8pQORxPBjhwfWdELKsCR204Q1hHQ
z/OB5bLLTDWd4b3aytaLgqyNUu0cARD27Uk6GV7q27a+flDMfZBfUgQLWemymInl
RfjvhGOPVdy0ZkpqYmxOZ9YhRNKea3w65tDuoqD7Zx5j4ROcHvIuW6Wa/1aRj5lR
TULEtJCfgvTBC/G11dyYPVkU+sq6HVPuwZf8gKoEFCvz+cL8jQZauUvMGujhkuOS
fs7NbSJYpzIDCaUcbl7h7iMIoah+Ck2lYGH8LI/JU6raZE9O5tEHvmigLmDgA78L
7oK6xsUnSmo2Y7kifJ/Q+I7mSNQwdzQjUWu4OmVTdg0jYKGFIijj/y01VZaSjKjj
SFAOoDi1iAVbQ3o5M2QaH6U3OE/CAsYYCsrGI/Dz/D+bt6XXrqNL2pGlLdj589ww
qfN3qJx7mGSq94yjMIhFTZ8utNhtO2t+9VTw8yBZm1Yaxc5ggEy16cdAjuLVccPA
OLh/VpyP9gYr5CI7AsZwP38JfXGoYFxPkxrQKf7Vw9eOT0kClUoGGGoDbyH46biJ
/2jMiknvJsS+rMXzOJSIntlWg2ZOlvhEoAwASGuAz9IDmkO41GMDYwe+oIa+rxnz
e3rTHQ5L2EvF80GqCObik1RPIa/iJUc1Gb8eVulSh/l+TLZPvzwop6DBYKOdwwqB
7+vmf3E1Md+YssSxuTxN0870RjhLBnDPprjXVumXujsv0fvDcwWAbXcQs0zCUEDj
WnfPMYS/BrP5sg1xYRzY0pahK0tW1UJ+AbXQPiwtLRY=
`pragma protect end_protected
