-- megafunction wizard: %FIR II v15.1%
-- GENERATION: XML
-- channelizer_fir.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity channelizer_fir is
	port (
		clk              : in  std_logic                      := '0';             --                     clk.clk
		reset_n          : in  std_logic                      := '0';             --                     rst.reset_n
		ast_sink_data    : in  std_logic_vector(199 downto 0) := (others => '0'); --   avalon_streaming_sink.data
		ast_sink_valid   : in  std_logic                      := '0';             --                        .valid
		ast_sink_error   : in  std_logic_vector(1 downto 0)   := (others => '0'); --                        .error
		ast_source_data  : out std_logic_vector(25 downto 0);                     -- avalon_streaming_source.data
		ast_source_valid : out std_logic;                                         --                        .valid
		ast_source_error : out std_logic_vector(1 downto 0)                       --                        .error
	);
end entity channelizer_fir;

architecture rtl of channelizer_fir is
	component channelizer_fir_0002 is
		port (
			clk              : in  std_logic                      := 'X';             -- clk
			reset_n          : in  std_logic                      := 'X';             -- reset_n
			ast_sink_data    : in  std_logic_vector(199 downto 0) := (others => 'X'); -- data
			ast_sink_valid   : in  std_logic                      := 'X';             -- valid
			ast_sink_error   : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- error
			ast_source_data  : out std_logic_vector(25 downto 0);                     -- data
			ast_source_valid : out std_logic;                                         -- valid
			ast_source_error : out std_logic_vector(1 downto 0)                       -- error
		);
	end component channelizer_fir_0002;

begin

	channelizer_fir_inst : component channelizer_fir_0002
		port map (
			clk              => clk,              --                     clk.clk
			reset_n          => reset_n,          --                     rst.reset_n
			ast_sink_data    => ast_sink_data,    --   avalon_streaming_sink.data
			ast_sink_valid   => ast_sink_valid,   --                        .valid
			ast_sink_error   => ast_sink_error,   --                        .error
			ast_source_data  => ast_source_data,  -- avalon_streaming_source.data
			ast_source_valid => ast_source_valid, --                        .valid
			ast_source_error => ast_source_error  --                        .error
		);

end architecture rtl; -- of channelizer_fir
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2015 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="15.1" >
-- Retrieval info: 	<generic name="filterType" value="decim" />
-- Retrieval info: 	<generic name="interpFactor" value="1" />
-- Retrieval info: 	<generic name="decimFactor" value="20" />
-- Retrieval info: 	<generic name="symmetryMode" value="nsym" />
-- Retrieval info: 	<generic name="L_bandsFilter" value="1" />
-- Retrieval info: 	<generic name="inputChannelNum" value="1" />
-- Retrieval info: 	<generic name="clockRate" value="125" />
-- Retrieval info: 	<generic name="clockSlack" value="0" />
-- Retrieval info: 	<generic name="inputRate" value="2500" />
-- Retrieval info: 	<generic name="coeffReload" value="false" />
-- Retrieval info: 	<generic name="baseAddress" value="0" />
-- Retrieval info: 	<generic name="readWriteMode" value="read_write" />
-- Retrieval info: 	<generic name="backPressure" value="false" />
-- Retrieval info: 	<generic name="deviceFamily" value="Cyclone V" />
-- Retrieval info: 	<generic name="speedGrade" value="medium" />
-- Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
-- Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
-- Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
-- Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
-- Retrieval info: 	<generic name="reconfigurable" value="false" />
-- Retrieval info: 	<generic name="num_modes" value="2" />
-- Retrieval info: 	<generic name="reconfigurable_list" value="0" />
-- Retrieval info: 	<generic name="MODE_STRING" value="None Set" />
-- Retrieval info: 	<generic name="channelModes" value="0,1,2,3" />
-- Retrieval info: 	<generic name="inputType" value="int" />
-- Retrieval info: 	<generic name="inputBitWidth" value="10" />
-- Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
-- Retrieval info: 	<generic name="coeffSetRealValue" value="7.8731E-4,8.3969E-4,8.9334E-4,9.4822E-4,0.0010043,0.0010616,0.00112,0.0011796,0.0012403,0.0013019,0.0013647,0.0014283,0.0014929,0.0015584,0.0016248,0.0016919,0.0017598,0.0018284,0.0018977,0.0019675,0.0020379,0.0021088,0.0021801,0.0022518,0.0023238,0.0023961,0.0024685,0.0025412,0.0026139,0.0026866,0.0027593,0.0028319,0.0029043,0.0029765,0.0030484,0.0031199,0.003191,0.0032617,0.0033317,0.0034012,0.00347,0.003538,0.0036052,0.0036715,0.003737,0.0038014,0.0038647,0.0039269,0.003988,0.0040478,0.0041063,0.0041635,0.0042192,0.0042735,0.0043263,0.0043774,0.004427,0.0044749,0.0045211,0.0045655,0.0046081,0.0046488,0.0046877,0.0047246,0.0047595,0.0047925,0.0048234,0.0048522,0.0048789,0.0049035,0.0049259,0.0049462,0.0049642,0.0049801,0.0049937,0.005005,0.0050142,0.005021,0.0050255,0.0050278,0.0050278,0.0050255,0.005021,0.0050142,0.005005,0.0049937,0.0049801,0.0049642,0.0049462,0.0049259,0.0049035,0.0048789,0.0048522,0.0048234,0.0047925,0.0047595,0.0047246,0.0046877,0.0046488,0.0046081,0.0045655,0.0045211,0.0044749,0.004427,0.0043774,0.0043263,0.0042735,0.0042192,0.0041635,0.0041063,0.0040478,0.003988,0.0039269,0.0038647,0.0038014,0.003737,0.0036715,0.0036052,0.003538,0.00347,0.0034012,0.0033317,0.0032617,0.003191,0.0031199,0.0030484,0.0029765,0.0029043,0.0028319,0.0027593,0.0026866,0.0026139,0.0025412,0.0024685,0.0023961,0.0023238,0.0022518,0.0021801,0.0021088,0.0020379,0.0019675,0.0018977,0.0018284,0.0017598,0.0016919,0.0016248,0.0015584,0.0014929,0.0014283,0.0013647,0.0013019,0.0012403,0.0011796,0.00112,0.0010616,0.0010043,9.4822E-4,8.9334E-4,8.3969E-4,7.8731E-4" />
-- Retrieval info: 	<generic name="coeffScaling" value="auto" />
-- Retrieval info: 	<generic name="coeffType" value="int" />
-- Retrieval info: 	<generic name="coeffBitWidth" value="8" />
-- Retrieval info: 	<generic name="coeffFracBitWidth" value="0" />
-- Retrieval info: 	<generic name="outType" value="int" />
-- Retrieval info: 	<generic name="outMSBRound" value="trunc" />
-- Retrieval info: 	<generic name="outMsbBitRem" value="0" />
-- Retrieval info: 	<generic name="outLSBRound" value="trunc" />
-- Retrieval info: 	<generic name="outLsbBitRem" value="0" />
-- Retrieval info: 	<generic name="bankCount" value="1" />
-- Retrieval info: 	<generic name="bankDisplay" value="0" />
-- Retrieval info: </instance>
-- IPFS_FILES : NONE
