// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Y6uYK1Mos1rgbtZd5SkJ0mc6Ggoh5Eae5ISN+9YCAFdUtQ5fBPnOb3qazzzOzON2
uQIa6LGZjDwZ8LXNCFQqe7cw/m3YUf/Lz9mONO9yIy/FqYoFaEwqPXPy/Av44Ve4
B+25YqE+OP4lEdT1qOebXEgT+JaaRCHRa+Q/FqFxj/A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19616)
SML3UcbEcfSocQZKpwh6DDNUoQPJAPzGzTkTaspVo8szn/E78a5b4ziQEJkOzDTj
tXzZDz07VfRn/lqDb04WvNakENS7qwb20KuYJJsQ6c4EZsyVQA0rAW52N0eBQNc8
5eQX+u7yPj9cv/3l6IvMGnZm7RHHyZEJi82dMzaFdg6nUtmOapnNP9UW5wG3kfDk
NZbGLre6Zs61In8VsBfnlymKCv7B4WlBGvwl8Dz5MvwcqwZRCnC95uW80zFZwLCk
Ke86amKRd7bVep8JnDuQIVHheVX5X2SDFCixXr58lWgwWS+SETLspEl2qb4mF/Sj
PzwTuqNyPUb8+ApUMCp88CTTh6A0jx9CoWT3QtmLZGlnvhK1AHKGMoCE9W4ovh4j
IFWDoerpDkfRcWgj0xjLG3h52HFk+F8d+IRkNgQi/zTl+tkNsQ/yDTeqCzqeS0HL
himH4duxxBlULGTiJsgss4cJCU57h7aO0YYVglvNRNDVZGOc4imaMlE0+JT2lw7i
DHbgm5WP6FGBagmHxF2+hTTiQj2qlOgFYcVOey5qhfzZCS8Wbj9w+exm72XMe6DJ
MEoAIMwBUNDlP3iyHwV1sw5DwccmYKeKSI2zo8Npyp663jxbwN7MojURQYljHQbj
gEcr9jMebTj73Q305/iP3EU1uUDgwqug8F0dRNk2zqZfAhl2NwW7Qq29dMuTG5sS
3XXyRSj93kDnH6tOxI4l1dzN7nZWTGrJaXAodBZfHS29OQuM5DjIdqES21pay0Ps
qcEUBF1LXDj8kP88jdoy0pc4H1KjIVFGB+iS4Fgt9E7BryouCWrHSZkkqeB6x9GT
go2wPDNlrAksN97zYLSZm/4xSUOxGFxJf6SBdHFn96hSN13/LctDXjzVJf0WB1n7
m14q8BPhc+D1/I8EXctDdRtJ+MjAe8/AdgqMHWp+vTwU59G8boAYqFjmRznPCIGX
OhpmPaeUc29DHZU6RVgMtsE/LvBCPHvCS+wmVUDvinipdY1EruODsom+I+r/EgXP
lycKtwP1IRzFrKY87W/sg+mPomyxpruN8KDY6e+pg1LLGi1BlZgN/h7llIxOv0NS
e7Yq7N7XotSfc/64OFPQHfLgwzWcdSxF9LehIDfsB8PkO+ZbOG/A6udIDC2YUolq
NV3V9jN1636+Y4euvAP/+KSa9zg3q8yKpqlZFBNymzAiMcRGffnb0mj1vLmyJ/Es
rFerzCoG6LuOmH+g7rI7VPgs/DytYt3B3EA04hc5wTbkO8Ua2keUAfCwXZdo66kC
+DENxdgjPcpGALCPXtgtp5ndyVE8VxBAQnaBMcpCUilp5lSEMEozaW5GO+ECgcF4
1HTY3I48uhqNOxHnzSRAVrNNkE/8w/vOm26ztAWxFUNOltQpyATYKKNulb0Z8/y6
jLQy1xNg9e+XZ811eD2ckFJBRx+62cmfj140WRaQBIjBwzcs1WiktVDhEMTMjBGc
HY+nFs1TuOlYfLhbibXPHpn3xOXvA3CQ96wFoE8HUJ9Q1wk2U0n9V5Zgq+Lk7Prt
Jw7AYvsxGafSdfxwMO+l/2nPgJ1spVGun1gRcvEm7Pj0Rzk2HtZhIw7LhdMS6Ndk
naCFGW8Wcus/7MnjLtnvV3gITvOlhYQLXc8BpSSjDngwyMvx8HaVKydQ8CZpYxOy
GO5MN1TJHkGyT89JsW6Lj6Y8wUeDIC0YwHKUo/RjrFm9yMu1oGoIcg4Tz9Wcss8L
Xfr3ZxnSiVarViRxHBVKSv//EYzxE46EKn45xwK7DKn/isFbGF0bUmOiuKi4xVbR
ix36b7extarPxqMYeVFhrzuszYRc0RX7ABD7wLYni6X9gw+INjFFW4kwbGhJPYQX
Egs2d2HclK2P9RaF5LyTQ7oxEZQMSHH18kLNuun1sDgZmF6kPayS22Fe2Us+MwQV
MtY4+zvgjdGWoS90WPXBapTSA0j89gG1D31cEI4Josvpb8+FpL0MrQvpBPYEsFcU
PBJYcEgq6j6qFUH8Fv+sGwA6RDiXuN0cEpevrxR7YwC7UU7QPPnTv0gvFz0CkDuM
pFjVCnrx/Iv9pv3Dk0oMhskNTdTKv6AlnaSZ5zQ5muiBOzY+EhI5g3XWI+b6ZiPG
qMoQsCfVytvoYvYDSKy7Jt+WruSaWUJgD4lCGKmTnYNDfRjP0E6tqn75XFQq/XAu
8ub0n4dp/BdYPTgGvCcndawrHMvmIzGuzb9xyGRILzTPr/T8wjrrN2GtR2gtfNw0
G5INZzEWWwXe5AFRldNXrt4gMMwbLW86rvMqRVf1phU/1W09u3faGCEhmMDsg2rZ
RIiZwd8L9xHupOPEOMTbvlj5LbxfhXxROuFaVyXJOzvJu3DXfk4e+3xlsAdCNf9k
jhg0TY+2mk+7HKMuHVUWMXPRB09JEQ3cN7W+NQzxwK7OSHHZoERJ1MaSLnNc0Voj
a1Zv56dwHW1hC80Qg+JiaQ8nJIpwH5JeSBdjcrWcnaQtbKoA8oMGt0vMptZAWdTF
pw+b6/15UpWpZP8nsQ0iK1hr7Y2crLwLwbwTI+KCRsSPHXaWGIx0on1IsKGn1gZj
4Orlsw57SPDRX1bpxc/63eV/av3tlcm7jB+/p1BWfvy43fqtuiKFsuMNNKGWygyl
l9XzLn6AExRG76qiDALjuF/41Dpp0kIAE+Lmxy25RJ/4gO60sr04xl/idmRvdL5c
fI37TqEFOTBvWeTdiSEt5KPMz29Sr4Tbsu80G3WNS1CIMLpJDvQN/GzCw9OmG/ac
HMMlxdSikJZ5mNuSKCDmINj99j3jYX3jRHpMWaRM3/J1kc16g4erGwZMQ4RMYQ2r
Q0hMPPuSg4S2T4/MPpZ3SLSwBxSczBhiWPuTkMdmqjhvQ3Gn5f/SOzO7D0nBBoc2
AtIeus9Sos5V6Vf6GWdU/lzf/x3hleCKuDwhMd3zSCFHrZYhn8uBk/t1PTMauxQO
3wGTZDpWVtd5IJ1Xt/udRxWzS93/7ktyv3Mgk3oU3rCiZc45hPBuUSGCKjtLEouZ
zTytKEF+4gjx9UkN4Q7YOY+yyEqWTDBGbmAqZASLvwnYCgKq5wDJncMC7hk0Wekc
6v5QLOnN2NFr3nq9cR34k9VG5s6eDa/uN+hgNPorUiGZsEJsZ2lUwZ/Qh0te2gKs
wmbms6RLztYpLlyjrd+fkkXA/rfwBavXwBw5wib5o/ay9Vrtef3ed0kv3yE/cg3U
f3U9ZznV9MbPgqaOYi+1Xxz4+FuR42/otr48Bw0dZ5y1gE64w+jcrJ7BnMzTpj7h
C1XWuQQk+ORBLaOUenis2Bo3CbwuIchMi2v6n+hroXibleeGdNOz6zcFUrhVbZZC
SJrJz4Yh6pynguwOkahysNo+UZY4y7v/PzBE0q+ZXsmtjo5XmZ/eBVPPY/84hbs/
tMJvOFXinBW6i9CeFov7dny+9V/s30v7soAmznik6G9+L9oZs3LJyOhtROtxD0X8
wEL4HnDmxy9rQS367BuM3anWCAck/oZthaeN95T4nxCvBAPMfzDJa+8nq5nOlNx3
cUavJ+m5/IC3xxSFMew/JieEfmRKK8TeOVB1EWb+RO3Thg0l9NamevbsMViz3POh
WkTqAGSx3GO8mXKGFypNz8tqHAA4U6+OHTbtCf8NmZJbj8WYIl8UUu3s4uz5MaqH
XnUeRe/vuf9hXA24YZZCgZljTcOjBKLWKz55G2teV+XZfCEpS1ZFUtFUqTA2wV9K
RvMvLv6LUC72xGC2wtam+mEkfmVCFgU4ZT2L1y3dMBwpW8kDiYY12M85S7Q6KhmU
SANEH1mN09eH1lXjtP2srSYI4zYcPY1SsokGRBPkFGg6KP/bFuRSnfj6/KITxRAr
RgUPorhctR3sjcitcCVzjvW1Nd6iC06SHcmmXt5bPq8gnYEkcROQ8qkeXLpuRERA
tb5Y/l7XMj4bR6Nibbggd4fFwx6sED+hAh2lcwaYrMmo/Y8t3D+ksb9CQsDuaCVj
mpG5wQ4/6AbYbkwFYqn/6BSL/xyxRYw2LZRDLLAtDvC5CvmNwnq2+iBoM/nG/aWG
MmsfIelkyzHIFlErlNWQQQG3B0Nigz8tJQ/kXUNagJpPkZu7OlKT8YKKC0XEce4r
TRnMWTqdVS71RPWG1/+2l7AiAPs7nWcKBQQj/4/2bSchb9syxw2Vcd8o3Br7+Bue
i5S8NW3UPN8GLXw+s3i4vQdw5pWsvvUvwhSXQOx7Xpc6uDhSlNme3V7N4xIUYLpE
gypzSxyhzH0VLyZohp1bud61nBXvbEewMo3dl3w3FjB3Gz0teDY3wzWaGQQvdfPQ
wUkYH/+MgWAzmoxb+d/s88KN1zFfHXcgKj62ESXLoeYqEz3/J7xVDrFVwuj012BR
IHe/9LIZkCzdQfan/yxaqNeuhFTFiliOZ+JhLs3Gi+Nk94y9McYhP5l+Q1W9w0Fg
MsE3OBZ7Ujteuzk79+hhsQOYHvxuKHu9394ORZ4nttwMABdXKVX4dJbobcxglwct
DeZhNcq+WgedQNZWigE8b5n9lhEkBRS+iH5SaRfiEU8p3tJyDojoxIVx2XCZI1B/
Rr/wXvkVp+LcukZu2zX1zRClai89pZCAakiiQyZWQJaG29TL7w1CcdB/WN0aLyny
ujFRQBSxwCPOLZhY+tYrzWvGvjbOsvhsCZZ94oxNXMZ836ZFb9VJvolfN+pzrpVN
GDq85jUe1JWYc4v0H4UHvdh8JJfmuW90U3NEjHM3qZw4ysmkkQU/z8CgZkcBNrVE
CkUr7j4lj2uUc0nG5JQq2YhpbdBH+9o1tzH3J/cW+ed3D1TCy+Fmw+qYazniMY5I
QLTAlLkjpMF4uIsz8+aIeMrDbHNN3Mp7hGa2wJDvAwpW/3g1GRCWBQziIigBuzcE
bI4M6wIxMst4XXn66UG1FfFYVRk8mtNe0JeWlkL0pJmSBvq6vq0kq+Fl98y+7ktM
wvJcn+5pN3T2/DZKYpd13kaeYV0FjaER9vD2mXv6vQLpEAxAi3ys9jggVUT1nnpT
BSpmn5Xa1al5CuZypnt6Bj9zlL4QBMoQPzxQb5CG1TgJiG8IBej5wuXRspU409ma
lP3bDg6XNuG9ll4nJmBVdPvQnhCz0PXrMSgSI3gJw5dgdE9vxLBP+CijVVfJCs9u
mRS6HEL72+V3Wm4YdC7nFlviyCgRftLeeEXMDJjbHyhDfpioKZKPFoo4lKy+RI7K
m+nxXYVll9l07KUGh2W51nzsj7sgoQQlhymk95+XYlz3vwwhaJb26Y2CMTmB/5Ne
lzi5Zi1Ay3kSln/yukNlDLDatfUeq38shk4zFOojzjGctEygAyjFiFPcJrQoQCYw
zVFwbIjSceJAsCTy+4plty4Y27nztDXYaKXLiHbLCf5T99vdueHskNHfEOmMJifV
dr2WeLmB0sBvi+N9Cd53fYrSg1MhD7vwAzRcRBJAwsig1miifACWIKMFmiKoMXVB
5XYUprX//HSqUtZtgnGfp40rSzaBUq3M9xmizPy3I0vfZ+tqj2+/IDHumyw1iuvW
AQIhb4EY9Bo4472igYWeFPMnVHqqgSZDnQeBT2yOrBZB8qJz9qKwWU+XFldrvUGR
vuwyt3BSv6H4qJltCR5hb5oCkugdfpS0su7szGulFXeWCgATkKnLcieIZHizhGkl
DLXHPePfYvNf95hx8WHoP/I1vKkfS3yUb2I/7k/LGFcabpRzRCejvDa039Y48T7i
EsD2NjJPTkOQXS3Tf45JPTaW3p5ILwa1VoPabhWh2tMg2FCYEVN6/igbyq2F00T9
Vd8Ewoj0uN9V6q1a8CaT6kQnQNksdsgoqoWCiptdnP9t22cyGxfnM8Qe3A/ZeTib
8BAssHgRS7233nt4SyhJ8eLyArjO+5mPIBPg1oWrGX6/1VuYzRSsduZ3OSfgZOiB
U0pA7FBv/wCK+iceq3FX0myMdnPPhQVWMfS3bDUsEdWo6qnV3ZngJgDpM5Adj4Rn
xhZeTwIfkkUp5JsMWj1ojtFGV3TVBsf6ID42bhS+LAV8oOj1H4WczNUs6/2FTwob
pXftM45lSeO28pB/rzxqqeINkV1ahtSHasEymMYoYY/cmZk3kWSZsa6kwG2u0vVu
buEcoQMgW0GEbW+QZBzKZ0nY/YRYM8UKAHRBuP5W+KY1JDYL4OBYGUVhyg0rLLUB
IvpSx0ODSkxzCpWhbf1cARE8s2CBzBw7pt0NxODK/nKrgL3aJN0Y4X3Wc3rrqhaa
E9RO9JCwQ9V+L3qy3ulTlT2ZY286emgEWE43f97h7sJ4HqXYs4Fd34tToCIraWC6
CKhzPvsnD0m57NodXW5W8/zz8vynZbYy8EP450aAaxX9M/BytTd8LSE6kx1qzQa5
kLzaZQPxBnXuI53ANht+67XxS27BFUcPgsp5T+9uzFw/tMu58UzYLP4v8d4qRxsV
wYxg26afi/mP8TQf7hkswqY4QuhrnK+3i8dnkmJDihpbfYZz/VVxtPKKD8AAjDuG
7E8PMfv9uwPWBD60xx9ApNjy1VSU4H62TzR270n70xUA2bfh2lRaCnXJYBWM/EG6
df7u/Pf6oUxjAv0YM0Ns8ULKuxUE341/uXzBcdCu05Yff5KI2J+4Lop3YI0cq9Gt
Mbw49eK/cw8ruuPRUe2Ds/pYQzhJ0621V1NLP+OfLBbtGCZlECHPOQhz+5ihLyPq
8vFxBIICwoseA4YsofMcUFd4c+sr15q6v60qDLA7XRYBa5ywmxBsdEhjYcNiXmYx
GN0ADZ34mM2GhTIF+knKEVQO7CK2TDlWP7t8gRkyo8Q4AImxsGuI67SwxRCo4Yqg
PGuay6yOLq/Jr5BQElixaGCs7YT8Tdc+YLlfDIWVtqER0shBY2UZzGH6xXpMMXIw
jcjyQzpEetsBTs1+nWVEyRyEEDKV3l0Rwbc0RyUqJEKejRJXvn3azq3nIEKyyrkQ
Bku2oxLhI4KBebqDgK1fy8+iAvV0zejzzKZYTZvi8OrJ3npD1y2bTbIhfAERA01P
uES4dpm9NnMVZ7btClkh8Xu5hB26OmUdt5L+k5i1Kj1oaMYnF4mdivs5wySV81H6
0uhJy6TiIsZtXnrRISOcaqYnjGJHPIFxBoObiqehm4nWFQqK+JVZYQFIfKge/3FQ
ZRLeod2ovh46dyXwx2Yc2gXjccQjBIomyFAxpke376tX4BX74kxK1L8t2v9BHObD
0sakcRx1L23xNSsK29xeFNAM55qkNPN6uur9WgoCFvO6B3GU88L7pQssQZKgXYlX
Pn8f6thDTpr8vD5VH7utQRRc+r59Zrm1Pcc72Tx8HDZtscbWK1tAcZKGsDAPMRs3
8QSHj7yQJSOJCBgvc7at551y9oujyHmz0UzleXFineEYtewAZa3HaeUAzGS8fcEH
W/MTH4aIcPJ7de6V68rQdduWOgewWDifqSo2i4VSGrB7yohAGB3jX5ZZ7o+XlbAi
K/WsWsBOseidM39v/QGk1gb0RcdZfn4krw7wlkhyBGALidzhmiKXhBUKaJIyqY4v
mYWfVC7pH10O8xK/y7GhQFa/R/HLny+cs0scQdCzruP1QJD1CMq57D3Q8hvHCfJi
33mSaWSKy6nWacTmjL6kdJc50iXo/yJIhSvIcU0IUF2jST8ZEiFL8baz9Cp4uT8a
rqSn9bPrPa2tqVvMo/7xyzMs3M0TUhZUDYB0FrJC55VfTANc3qxe9CBBGdowEyAN
h/aUQhZY7j2AmbhPnnJWL5TVABDtsPTVXt7oAEvzbZkzhrF7A9QlfDpW9itxfb/Q
wlCJ9Lk+nQUGkuPdyZbBx+ByHsAwgIqD+Jm0Zq6xGZdWYMZNlnEFvomnX6Tc8b3e
racpggmo2J0iAdqZ+52ojeUDYYm87UJ9lmC3umJ6jyZ7BC33xgrWyFHB6KwMggqs
f6SfIjOdFWpQlCoygnAL3E2swVgS0zmCQa2HvIxlE+uZjq+0qEAcsL4UoIuueHWX
uYZCE/zSLn0yhIJVJfmUZzL1BZJ5C7DAX6qo5/i3j7pRXabK6/tvPPqtOyUr7iJy
ArjQyz37wxnc/RzVB5nWbu8R80av2RLZ8BfAByPhVmLiMe3LO8cSoZfJw6vb6z4g
SwbYtVyneR90eXFcshTs2+gXroUn2bcEQYQeXfLZRf848KBh6aT9MDy9SEu24UZk
Q58uXhSoMQujA6GGPqvJN7wzvEgz0lxJFQuLUZaVB5NE7mIdse0VyhPt1l8ngv5k
ZvZEnRrZNqUI4/z4LsHNRgL7pO+gel64KOFNwtgWDoE0laCJ7RwH2JnCfv7V7bnl
bON6hrj1ncDfB9Nbyl6Q4zcDkLo7ZL6w5asKqoui6oW+/aEFKpIokwgjA3kdoFpz
7gDL2DbyUVT1PCogV4jwH4GoEAbWacPQ13KeX9aBzaihncwuH1IatSk3Z8fRMXTX
EISCvv6Mthgvp9bxtv3GH4fQdBldcj4WNQWMak3RvI5vTigU5VPEiBwU9Zoe7o4S
msgtdnld4VgaIj/sEefJWtR2iLwWj43LTeTMRpLR0yb25+7He3fmaGVeAM/D+pK6
+zgVL+K/wQT0rsi8MJc+a6ukX/jkwAk9vVwEosMpeM/um3Mska8OafObpJr1d2AX
jFcwsjJFHOse2l+ZuBXnnLXMJW1y+sPb3MkacAvN0PIu2Oht4XzsbX9iuHwqa9Om
mfGt+QzOSGw8NwPyR6ba+T4FzcIVCXO4jmE0OsXfHApulgtjnbMAjw1cq2PNBHUo
l/mtcIZ226Z5Bk+Y1e+05qbGDhheMa7nWgneNYJvhaxStO9w34c73gYRf1pDWPj3
/v5rxoFY4yEn0NH4FYPJVHJOR0UF9yXzpE4Hb6HRZR3bA23y74NfMkYnU+9HC+G7
TH//QlJb6E1/JoSUkHmPipkc1rGH2MKhautU6z7NvPKG09Bukp140Q8FTTqZTelh
50eSK3U+G55hGiXDtzdW6did4m/TFfneo746Xt2VyXhhfxytQXeCnNq/d1IWxBCW
PCSFgPOOukNaaGeEqb90OaUeixN1Fdv32xSHZ+03AkBMiT7A7RI1kM4RlzwBpxw+
JR2/UEkIY+5DuIOiDg2KhYJps/7IjItvKMfQPrcXNhMdWObV1ORxZ2lRMfRVmZaY
Cxbcs13KRBonM1gIdqu8VNz3cYPGqjnASMVUYDQEZxdA+pQYN8zx7NmSdYXY5ATz
uT9HUvyKRWKgaIomfyTVEgZ2YABBvhMeHGCues2aHDMS7NWdZb1i3+cXuEwrLR53
LPPIeTmSHxvN+FiiDDfFj8u/6TU5qu+MRdxZklWF7xbAK/5ddPmwEOIQ9JZ+fnlu
CR+8AaRZLJNsWXpjIZhc80+EzHuhYoa+8K1KRzRgAUjTKqaDrSrWpohSEYo51h/m
ydSVNC0axjfFr0orlNkqDkVBY9ftknREhNL2SyN0G7ThzDNyf/Fr8M4yMpmAo2WM
fhJv3CcBc14YgNk7htDhUBgjO8iBTSJkkd/7bwLbM50dafIMZDeZL3v0itBihZBd
jSaczGvCUpgCiR1qgWmykVAV64SsjvUcRhvy1hW+BFBFdgIbi/rE2PJAx8G5DDok
FbANQlXZF9Evi4D8Mt5muMzpSs+nUpDtbiYJ2sWRjj7Vx0OxQgI9I/G1s54kuKqo
1EPVK1Zl7FLWfHSZBob4/Zgbs82HvCWs3JXW2CiCbyLsieiP/QgvXG+h1YgrOegm
zTp4Q9E/F5BSZeD2w2o6zNoy+PD2BjgWFZ77fywuqS4w9AVLcIme3YSdOwCHqiTr
Ne7UBENjIf0SFj13Bzol9tHm3XOQ4RjF5d/9txMSpmAA+HqJ5ItMbruilWcLGGhs
ZWRMoDS0vB32aEiuhoUQKpdACwC7+ouHzbkmLGJsLJ/1INI72dHSesy6Xx5M7L5l
R3iSRodFfN5svYEWEyguB8cKyWpvyQBpIS9S+rIX5VdHe6CC7gIfJDjHfK7JGjxa
tsGpToh/IlaEt9tmlyFYg80Y0G5DS1KiC3DMyJbKKGKg8V/ORgccSv7tEHRyq4pj
exKtZRe7scuC9ehfYvhtnyZZu4zzGtr54TMHb8xBTQWy4RGVzBHHK2GuYbznaohq
zr9+o/4Jyfzfd4X7mIHuhYtofHB8+EtYIIzctYm1e2EJGYMUKJhW93d89HGLDTLy
Ci+phEoURNP/MP9yaCBy6xuOiORshuSa+JCGZ1YgcjxqtBNm54rDJTnDqud78ivc
03pEFatxENEfVAaR5yOQZH8YDePq8b0b0Aw1U1A4bXSnymroo59n4yZ5mJwRLu4A
88jZc0xWv3owEdbizxtw2WfFiu3XYO/YE7/3JGdGJkyJ96uHu4QlXEeYCaSeQZDl
pLytb+q3XHsZt6mJEpd+vMgAeb7zSNNIAYo4NuTj4J/Y7y8k2N4IsJj4bFHhX89o
7VmUzUpRR7/Sar8ukIIGfQGc0CzmtxIQI22/qHR6/bBP7uagENk8QeiHvUWNEoMb
s4DZDlbHSPFNWgXz5h3L4IDokOQBKnW4Ndd4OdlcT2TMZ9Z3Gd7Am2K14Cmxlnpv
iRF2KaONV0jDh6090R4jqoF1w/OWzm66j4DzhE3DbIujKKs7Uvw+mg/b2aClpP1z
FKhYFrcNvkZfSip0s9B1UZ/Pn+oEO5AJi4mApYg/sTerg/KADXP/7j3ZCy8wJB3U
YcfjJgi5RWERLHDUbdJYVMEi9XuoAOvlCov/dGB4jTltPIXe/dvsw2HEgT5OAqsE
ZR8WqkCGR51MrjsiZB5ePPRkxgJZENmnq4T5//vkprXQZuYF80iSge7qmSmSn1qN
eUNfxy7XtdBWf4Rm/qwq5B0DdTT1tXvitAj6N8CKaZd1bGrE0vMOWI0pLrQJ5xLy
Li3Wjy9Xm6uWX3EH1Wrue+I+m7Vha3KrPSZwcQCMsDb6YBBi7EQpPMWdSKu58+Tb
e39vG/lTKDujZUdtNP7O0oAeWHcerrVPhZUy0rJo4zJ5ZhuEKLddMDbkDpofbbCL
NuWfC7UBH6+scV1B6eA5EFv/fEUgJksdFDh+X81zCOOCENwgn6h9JMc1DC3o2w8w
XjQxMsDPgDawFjRb9zwmzasKZGLrWwDMJBLZL5d0QLtsco+KRn1U0flnDTFCYRWg
E1yDdxFEeXilxVfOGwKcsSUAyXiZ9ax9s1atw5vY1P2pXhTZVn6Vc3FEp1/sQkal
IquVXECzFDuJX+QD7U8P2Q79HWC1VVNILhtOBjv+VqwvjY9Pmawx2Y44qb+Yg88f
S49RSNMlKivEw89QE/72gzeuBtXBlQNRQNIsd1TFz7jsqOONbtQbLA6yKRzMHGkA
PY7h9h9Ajtq3fsck3ZwkDyagSN1al/N/oj/kS8vfNFb3K08NdEHI+nT2zcQbsPeN
P73gt8Jp2Ue3ie6qZmFzEQaYiLoBpu4yBzWusEIo6SBpSDq5o7y7T6FG9mkF61Px
/cd45kbMS920Q+GsyesZJN68yN9Q7XHUru5pBBY+Tn2Y7k2BMm3FM0q4faArT2g1
iGn4wYeXfx3kOKD7sm5s9vblBtrTtCP59LYhpRCkb2i0DPoOf9rktV+FaYtN/lyi
n2nQ4s6x1/DNkw43ZE+DuANlllL3w+7lZTTWcAoH82lCIM1Z+4eIEXXnKgiSXcQ1
V/O+L5n7Zs5SvWmjAS0eAY+XcsSbEORoxeXdPFVKttqp/nsNR7v9yDaDb1MhvRBM
cZOcDxmdpHvRuteCKSc7nYUBIAl7WgSu5nDeP0NRE5S31hD72WADBVsf2ne/fTCV
IepnB0+E+ZP93qs30+Cs2Nv7naHB41yeVufZQlAb+kFcUhNFGsghSM83CO97kTBK
0m7TT0+1qa9Ql86Fp2/FlygDnADKrFN6peWIJzyPqfta9EWNFB8aubhI71IH6O1q
wqclNr5HnmBgGCMbCK1mQjtU6rGy37+k/bGvQOfmbyStC59lpkca7cbnAR4HSFBI
4JATHVbDAoAi5I0wOpqmXJOMzVTU7OQzlhgLyeKINa0nht+0+ZDpWUFhpPAtK5bk
4TxFIxZwTCKBmNOdWvY7MvkfvW6+UPdOaTntoLbZP/iBhFmp0t1FFNQrBGF7XsHc
i8HzwoFNaBrWNzBgzGWuFsYlqHWYk7ov/Iy7SJL6QDjClBtj8QpLIClSo/3YGTjB
mMtpmhfCg8fnawr1HCzgIQ6515UESYEYKwPutBvEVLGWEThFU8PTsRLUbqolbNOl
AqyXRm3dhEwa4aLpySIsGgrribhM5U53HFfgKX6ktTJxZ3hoVLDTNujv0JTc4djb
b0qBroYi+ipvi06qj6COXWO07RVtOgCbd2uJni7AEUZPDLrYIROYYUQrvkFT4+CY
Lk16AMKJFZBRAb4BiMVqMPdM+ow8e+h2z8O9kOPEy+ck1+B7Dg4CoBNdPF98WZvA
lP0y8jEyxWlnwdbct109Sw5PFsPQVZeWqY7vr8/ukQ+cXuVE72IXkQZKLYKs6Hnj
1zRYzUHhVEGp71ZP4d5LSGgypHtZMaOdy64y1qmf3czoidaBU0tLLMcN1KRaKbwk
ZeXlS1pu7x/ctdVZ50Pb41RpYTKx753VINxm061xd/y4VNCyjMBkWwhj85dT/+Ad
K1AZHWbj+N0H5ILryRx2c56JNlMJY7z4+BEqf+VuSGGK213gNekqLhtz683EW5Ll
IgO4Qk5hZW8Y6KT12rkA49YfjKCSLjVjlT17NJu1ssKkltoZwaT4ZQWOdqJ2iRD6
rt9pnNHvqdNss1pX4UXMY56ht1ioRTds80eVPoeWhkDsS1FNt3P5II88tV5Iwbog
kf9G+eOLfEuW3ZHmpwNvHEYB2W/JtJ3THfb6pa27baHqTDCj3WEm0NXxzDvHN8w2
GKccSzyl2seq3WvwKwQD2mFBMQZQPmd5uoortzcBxtdHhDcAC//ozrUZd/5dOox3
xHF67sfrI1wN0SdX4O/HReNT/xqGXkdT7TRUFFM+Tnq/wdfWRklLgDCfiIB5JPd5
ajT7GEyRQRKdF7zgMvBAMrc4XMHMsL4AuOL6TQ06xGV98lAB95yaakLWyykgltBw
0ROpCjfXKlaxWujIxuNAu/++rxOPVJ4f+MtkosF7qGwXdlKyZlN9YhPKB/GJtpTj
ETmb0LYWeUqpZZDkR3ODQ4R0PeR/J5WaVLrrLzmfPysS7GSKrjFuSxrN90/Dp3Nf
J5n5Q5mMCFAgCuib9NYPU7nnXVEwtXrcTpFLSxxXPdMVspYTLrvFEuAirAlrmFhd
Wo0D6lRpjiR2ErPLeo0c5tyo7SEjRSH+FkQVh3V6dkoxnmHKLzeYZ6F/fXthK+Bp
8lp46prIbKNwZE2dbQDemSQhp/0M2qgWP9S8CsEaVA8C1yO53ArfeHtx4OEUhimI
GYhlVNHC0hiteJQlSrc2C7SO+SO2XOd7ia7l6lwZOi8rQTDXpGAkCxBHSih7Y2bX
d101v5MMGNzL6Arad8+ruKAghvHSrr8G5xHk1D8qF/t5GVJVL+LCUJ6JT7gEwxnB
phTPWv0R509Wf/8U5InJwSDPFLbLAqKNEcN9/MWwYG2yALtndkV4DDsL5rbV0u7j
CnDAfUHEwYdahPwnJ5orRCmjgOKLqcMiEP9CeBQEX148R+mFF/uxD7kKjc9dIDW2
jquE7LwQt0OkHgNqhc8Wr2y+DKeP1FYNI7Pqre8R0AM2lR3T8n1ub4voyfkHN36o
qHVb3byYASp2H5khcxLRvtxLcAXzcMg90kBYvOH1E9qtg2AEQXPvUdAKTiL9Uzgu
qklcrcZfofXLr1dSRz5SfAkdNIa61XIBihURqsi+IZgGVjcDhV2PWHJ6G/QdJ6G2
g7KrPzcphzL1k3Ez7x17BTqdiygypDFkoM17HoeyE59cCvv8Pq5nxCyCSsJu7B20
/hE81utS8eAsGqnA90poxwQNxuCX7JYsDupPaNhi6JiKAFyZEMXJum08T/zvuKSX
xPYHOekxrsZ4Yb5QuGTgBzEuZIxLW/z1+YJd0sZajRIyzinC48ZNL7IOX87/J86v
F/LihInph3UfK41NExHtXoWnD69jbfYSewVHabQi/eYUq3iQot46I5f12ruqQg5P
DExvPug3zo+jBeVAtCOs4NGTxZz1o9Slox+/HH66ilfHCDSS1hGKVf/6huwYHtSU
VGEnElfXPvS8xKZfQmoYsdwJFzb8gRv86QmYvsAMX7bdc2dSmoQoZ4ZkI4LuBRbh
mwlRUjzvmhd7uJA7IghwwIhc3BkmZeKm/RnpFeVQIHXOi13UjP/WEr5ZWyHCRU38
5bsx5VMDp76Mf7ljpcJLz1+hN+ebVcBe32l46DCJ7T0zaR7AVbtbjFxfcO1PWkyW
fzXjg2VZCOdinWLTk8AuwfnckVgyZdmO3IzZe28lfASM9x8ENmoF69btwn9HmWN2
JW/9iSE8Q11VStHhg4hIAekzkUZ37RVzKazvJPZXlI/8JhAn3A6q24v5n2V62+Sr
T7WtyZeulnd9aalZ2w9sw4ubhKJeFcQ/07TaZwycXE+I8zo5kDfbEkznwK0wTY2C
VhfG4kg9w1RFTWcce5rJBZ0mdoQklxWwepeWT5HqoJ/goT9eFD2TT6yD7mUh5qO/
NC5SdUoThOhIYQRONiZmxYEe3AVHweUFx3mETPGmCub6Cja6RqvbnZHnVF4ueGU0
jYY3z79YRO2ZiSOC0OaCo76BmSY0bvGeHORoUhjmz5jHf2WpGZOw+bqaXduPn4ug
ydNNHLz1kF+1FuQclxB/hv4FH0A1oKR2Bjr7Jf9SJ7h1FdOQYnezrZzb8nGU/wSx
1ercRaacKuy5L+U/kg+mRfnjkS6VfJVAVymhQOEuLldbX09K5G2R2t4gQBsUcAMk
UkgkC5QVF+ggm9GB6FJzbVOmNy6YBcGn5FG95HNIDPz4hLITuQ3mAmq2H4OAOtFl
oplyt5yZurhcIl2mluVYMqTkTnRx93mJZtn+Q7Df3sNL3GpB4Q4km7lD6eyaAgMF
9HNeZgOeIJJ5IaD2RNz4L1lS6VzA1raiCRtYmEJ0ApXoze2lglqhDiuz4+VVq1r/
TEJKYHvzhi14bXAOV/RmRlJ9vhnub0hzEzLIKdM5Dga34+feFg5QFcVRtN4vhb9T
NuK3tOgMRFhHFhlUf/wnGiW/1AJyQ/SgvfWLDo/n5fo8HVrWmVqTztfQaYe5D7KH
VJgW3hPw/axzcC7dZ+Sey2e2c/zs/2cqpMLEdnYDHjjGdfRb6tUWOcyQk8CA+RkU
9A+/DmPhyYpBtx5mNZm1C5fZ6jGYko5cy2GXNX5zGugw+rVA3hcro4rq/zpuM0x+
URILyGNtjM8Xug5fjGeXRihUYLS2u7+imUSu1vReInxl4J3Rqs/WmW+sXww/aLfc
eC0IerDDFI3X+6dGds9IfDp7lpKSUQ7YOL9rex7iGg3ourf5TkGI4IR3RYTzfeEd
kniAFdULQacAAMYBJ8SgDQIgkTPzs3PzzxFYEWQizzwZMGrOHaMAfcMu96L5Ytau
IlYLm0J5SNR0yYQWSznysyByGN6ccqkiZFb+GfuchN2l2tdia8rl3MIGXzTOQOuM
+WJ5PJDMhpJ11ryW6ZEIakrQZl3smHn6FHSHd1l35dnwFIXjid9D0iY1HCJJnppm
oYdfXuL+/95xdGwApuCG2N9QTWfXUHkoOKDhNoF2EeTqm86oweb9pxEzwczdxTtG
dFL8Go8vqBBpOYd76yV5GeS5vs8S34ALY/eI/gVaZR9nbwQoJ+YlNRnNTH3UspdK
iPNDzMb+pyH2KDnpB0HmelwYOkxdl4aZX3zLDnsIkoWE5CCliAEQQlI0Fap3188P
A6CFv+2+3pP/fgN35/cyhOjV4FO7NUO2G59QUdyDctEfwQ3ixngbHNeZCefjNQ4s
qhzME+CFFnLdh6vYlrD2mf/mwrf5ZP50KP8XuVOjChUcRutMZKA6FVyqITsr2pWY
hkPrH14UPjsOYYcQVXzg5R0+LNw+LgzogiYs4Ed2adW1r28dX5l7SltBHnJB8nK7
OjvNZ/VOih5A+EFJDir+FHN7hUJWW6+JCoPRgFrhIscuUrQOuyR8K2XyF/EHrlAI
b70yw4J6jXTBTYjTH6BKQpr4j2u6cHpSPTTkhvb3PuLjyqU188Oif4fn/4aco4Zh
oDvH935cFXRCGlk8wT7nuD1InHTrtLfLdSSTfplLcX5G7LedDCR0NgUCWvYzXOaG
cDFjsUKFaV+8XS5Mk+HMypTiOTK9FAKgI/ukhXskp08joToY1qDr3AeUCFahltsT
rJ3IIku5I0bQeAxfQqHXE0PpuU/76AdsVdu8oUhTk0vFv9l2UL+jECHs7+Fu7WCy
WVmV34Fji2fIKrt0qtTU5bQ3p2/8kOuGRHhrs64VQNDPFJX18INb9kqceW7nLKwr
lAcA1Pmbv6oGBPfv5sI1F+8AUFO6hTRqdTIq93KqHPEE9d4IWaEg1qDH7F6e/1rQ
hIQia41g5f60Kq5yZb7quwNFEdFlY6NdnhCOUBw77p5Z9ZliEg9uXU5okvTm7IaY
+JksIy7y3VtKr1watLoGZ/AxF7nssRrNz/D5bpc+Rz5eYYG1+XsHPoqRMp0sT3Xc
QkrttzkUDW53yDpHAWVkZ4sS5KvzTrR8UUZqbttpjoulGKBv02cLBdZWCCDQtiyN
FccJ3u8+iw4OJjk/RMXi94fPzrhqm0ILWV023tTnQiTUOmdiLNimH4J8WsD0oCOf
oClJX3LvuEV3GWGtg/VOilMwM821PzqPMG6WM6c2bUBe80ZdjbZilMj15mQ8mRX6
Xe3VIsg3k0IRjuZyI96YUeAK9DbcK/fgg628TyAFiq/2dREPMvOXzv/dofc+LEB2
KBNQbaKhQns0/QkPY/PiPJGZ3ZSRi13vQW6XcFtjF/S9TlYWyYetbPR0Z3g9SzLu
Mbql18XB/GWF3bhjL6x5q5ydpR5jxlmu0Fg+PJMxnVzfIHoHiV3frPH+uC+bV1c+
dozdiR+xBTwNEI0zcKYNFi3YFikC7HBxjJK/VivrfSSK5BUh+rrxD8N+ovKqf0Mz
U3myNJ6V7eUmNKA3WSQDB6zCjrckEYy7r8IkD0W6njgaKI+K49YNISOQHmi0o4SD
hd4i0eBSzHDzPF/L7G+Wn0gzdOyoYMWYcodIimsWDigsXptc0S0e6qogeUAIbCIn
JHT4svz9nQ6F8qhFRxs+3Dv1vk9fvCAPhP6qdZCVkxRQ/buh8/ovddtPaCPvOTHL
WllSexUdQ43HssnQCjh5crCmYSvkhX9LKsSLYfE2MQKuaMkEffcwH3c/k64SXctj
f61M1zal1G8wT4VM7Hy/L8VFLVC0KU4fB5/HyYQ4CxHYqXrHpCGS2B9uW8wJkDDU
zq0vOG4HPmgaLCV0kFkpFt6PQHPx4jbDhNhTMx3Wxy/nRL2xfnR8r2YwnoT8QThj
XhD8P2HHXnvNsdnDLdBd+o5wcxtS/HzbaenhPq0JugbfDiecI9g/KSuqyDGL2l7H
ksLoOvDFH0mELH3jO3RpMw9MEeiQ2KYA4El70CubDu2WFdKVp6iraANoTUwUrrWC
leKiYNQCC8C8H9+zrdtz608x0VMeQUmuDKnOCwwh3dBLh//XdE4S49W5vXWOcAfY
yFU5QdGpK/B0xXEFHaq9a2Rh8vcFQRMcVmI02pV523wPlF/ef2ossSd2pBVYVwGT
LJk5EvaoL9IKMTb9IYesgdUnv99RLGH2et2J9C6SOz/hgdkBZzFkSSanCY2lbJJQ
b4o5Am0v7a5i6aeOX3sYkw+YkAv3m3EvkxgmEI5YKpYy4wJ3JexB2TGj85JMTQCp
xv2iFX+NwX7TAd1UOssgWWgVxkxc9rvqsopkUMLZ5bY9diGatZG/4M2dJ68YRP0J
qdEh3/iCQcaZGTW0LwD4HGq7IMWz0c7hA7Exy/25oROiYO6fYvwvkt5KAMdbMil/
+Mz5zFB3rB86ct4lCDA7V/TSzv4V87auFpikco34yayKUGVYIkGE3mC/5SjgD0G3
s0qYj33G5HB+/eDXl3NJnvSsn8EIsAZsFYedqOM2nN+PyOX3gpJW8oTDpu7Bi12e
PJy5T38GXksCu1eOQT5q2C1gm2PYH6LDkgROeIe0hyYmlEMCaKGftRZVcRp40HFh
UaoaSIWHWnqdpL5xA7wZfqWO6HsITEYuuVwuapXqOHCXV2YqJx7jjnLChLoUaDtr
/kMWpXFtjC2hkJagErp7WtbEDGr0iGxtAgBbeCLDIEwnkZ1bG0XAQHPlT8BOEYzx
FkEklE5QAn2tjOpmeT9VIyfvepnir25f3uDx+FiG7VC+qX8ZwUNTEtUTATO9loQZ
knG7aimOE4pn+br8H6Ff5g0v56dTHm2nnkp2aXhyC2GHN+PbrI4PadjkDO6nL7EP
t9tjMBhcfP9mZJLBoOoyUh/5hD1Ozlv1KZ/EPy121rkSMx1NxbHjDDR/oOdjytQY
GqioQFOwkLLk5bXcvFk/uJb0O7eDNPzuwOYaWj28MgLcuNZ+zPjqhpmLc1k+kBUD
hfOj3XcQjLEx52jyd5MBi+tKtGg8Sp+JzWDybRfF7IIWTwJ0cXXStC/SZhvG+kDx
gSUjPnp0UWZNYc99nKJSrX6wpa2y0G3um+I33hbzmMlJerqaAlHO7FClziA0Cjkl
jz4LTHil7VvjZc7wDDDxXeiNF/ruv3qmCHcxGwgWf2WJn8FhS2UyDQvv3Z0b0BSe
TdtRGb804vqcRHPptjph3jGUDz1usecc+Tj3D8xP1zSmH13FeOhsFLcfKx+Nj1T9
TevMMxWHAtKQtLTFE9vn6ei9OXQexIJBDpfwvl2JNKiKP0XPXCIvNXS3q3RnSBXM
qE1YbsaULcGgwger85RJfRvOgCw4Av0HbjhIFyxZUZiIozK6RMIZCuKBjDoo6+Xv
BFa6TkDrIocytU4J2MxkRIChheCe7aJuZB2Se+8IiNtfMMOFoEhBTmEONpJjNzQd
qLOZyF3M8oe+CIwzvl/6qz3JeeNx6M+8KKIlZUqtLqhTEZJe/5kTcICBMyWRP0av
2dZFAFOl9zpUR0OtR78h3DCjLT+srLFoKoWpPIinCuWtNkZX+5rqsGwN6NLpW/il
TVkHdt0hPFUQGQ8Y+f0XjgDzQE3ou9Fljprc0+TsWADA/jd1aq2W+AB8qRl4mtPJ
+l+Ylg/KsiadUg/RyxQ2YqONrrLsJjZaXEl3soZyAgdVsjzdC8DRltppf6tIX6F0
oAd94p5KGBAa/1ubUE6FYOk4CERHxS97jsRLE9N7WPKtaK3KuwRdlWatno2ir+FG
7vq/fuZIw1uE0npTPVVj5/emUfXVJKPN5n/RjFn4yoLGNK4jMtXSwqercAHZS9CS
EmLGXxJQWVjez0B1867GGDepwx0ygA279IyP2lq/sfiZuBFJKOh1l8mSBarsQ15L
nxOVEk9zFOWwsKu45tearA4A4Yyj6RRJEVphNzTQLCutB2V6R/8dh62v7l+/xQWw
LxmlCmBBwkFmR/jCzuBze/gpYC58hElMdbtO43//lwq3qcUXoVAeppepLPjxwqXN
EdlWkYFZgS5iWcvXba9Q3+SRNhJv33jPT5U6vUJoqWzzQfDKxn0hGvx9/B5zUA+3
GmbF3jPyQe8F0PmsELkyG85pBNjUBN+dVxtwYe0l3xPoco4yl5D8xznYztjioEhl
fTi9u9i3hfmiCuz6/ZtatU6CHcppV3Jjgl5KOXpV/LgebF0UNE022B4149eN8FqF
ORPcASCuXtYdT9l5hTMRC/07EpNqYP9LhJ3fv/C/Kpp/vNAqCZURzyq8pySAeYyl
fPseOjQ2c4uhMlE1nXaWenTEDfCi11lEXtv8R53HnV9VEjQaLz4fvIiG+Az+5YXx
AOipp0VYdpQjnIJKDfRTrRGvkasuq8hcs1x70f810md/4cK9q0uY0H8pxRivlVZI
2tQTsKcNDAiANeVGOaQfzAQ6Ueyi7pM+s2P/YH/5MaooSKZTDEcrqSA8TCBGNZu2
IJpmbwuZK/PWDJv319ts08E6YeuI93+z0u5qaVNL8xPm4V5uM9FZPGSiVTo7muEP
+wEp9illdYOwGTyoCy6dibXbUnBEUDZBb1yj/TB+KKedgQYokynceictm/hk+KMv
S7b7LVtn6hMJLjPgkPBQ9U3L0uqJrz+Uz6VyIh9yKqv/hKLLCpT/PSrvknE56snp
eLaoa5MfL9+2+3f8gtTfNnIiiP9q/gXuiM0P2q7y81kew0f4EoZZtOOM5HXppZH6
7lFrIC17BfFU4NXs6hVLCh1o9uDPKFwOUorf2MxK9F3jXxFiDkyqrD0U9w0gGB6K
tnhFasNfQ6j1RD0s8Il4Si1FwCCp/3aQW0fm/5NAw8e0DaZisALYzg4qMUUnuuPU
EMtPhidniY4SrxFnnDfFUVM0tWY6GEma+ZArWhVmqylUWqxmBD8C/2OaEvrhD0df
T8XeUt0Z16JZ3cr7YZzkGclf1gfTNkZchWp7UCUF+aToL+d0gOUZVSBAYFjSHZMA
U9/ZnjdIhnuYnw3dNlCjq22UFYFmHJ5rR5kWk2tj1I5sbnV/eK1/Jx4E8H2SQQuX
ZZFjN7v/1BQOij3PopeKXt6FQSDLCrdDp9HpCucw+DFb+z5eClnruUqVfhQXSAJE
66g8+yAG4L7jfhKO5509Bb26LDgAaWvwWniDkclTBbdbLiDGlI14BJ8CUAks8J3B
yfEtorWOuvm4Wf5+bNdzJ4dpKnEnyYCHhdT7PbZH4u6nJfdF5pcy1s/c9RhYYFhP
PpJ8oS1/rp4j/wI/ZI3dWHOypzwIt518KogfDJJr8uAoNZpDcAYfIHvCWZy9Amxp
L5Zrnia3ZepWqkH/Hv49Zknw5l1TUqWi/Im0FC10j7zV5pU5xbM2m87cUGUC9AyU
6oK37HHeEKM6kfFxSfl7myCXOht2QlfiO3xoYsDlGJkQshbpYd4/qv/iNeAuNuKt
xsXBGtQ0y+WWN48mKDlULHWIn5d03GbaLBgRa58kU4DJ2puwLv4kYnkEfbqXc5iY
gJit2z3Fj5tTHG2hIRk/aeuQn5kLM5lbnafILehpFqDDeKOtUUm+Ex/xWO2PW9bx
qITx4tIhWCGb713/TKorPd7fJ59/30hWVPsvTOMjbwFrS6Tf+zCnBbpMy7NCrxMK
GoVY1F1mWVcuCBQgqpiUpct6xKeQCTPN1HgSSqB2nvu56NkfrpOxbF4a2+qTMsaN
XjPq+gDg38Pg+IwAjb8klWfuZmVSOfLcnFA94QjXGxikbIKjWglF27B1PySTLm7B
DlWRhfS/GVYYRBm1Lg41YTiyswgaFIFMds0bjBcySeHVUIVLAm/N/InO5qrXAruA
HpJjpsHQE9twUI9jmd4LDRzwIcfTxxlUULQ/pY9N3/zKcVu2PLQZ60JghGV+Ydl0
/JKUylM/qdLXUXJAsaHCxN2v1kRvyg5V/ecw348UzKFfq9zvQLgekRQjW+095TNp
My2knzSc2Pw1moPINfy1sjmt8bDqejqP+pRnQE1AT27gWlOYN+XeVRq6/IXPxMKv
woBNtT+a8B53Dh75MV+IGKRyYqRwpatmBNyQFdTbryRrZP49U+9FTXzo4fqUqV8c
aO8ayL050QvqbR9xy/Tdsui0d3ZsEcZRPLkLNruZ/dMQWa56RbF05wmINvzSUImg
215V/vre8R8YY7nmBz0YUIJXoxD+XokY+/774gSny/2C7ONUjdjegnFihqeXHjkP
w9eBn3RI0bu3BT2uLTKN0b/Rx7Qvq4QpHhJ8iBLph1vJlB8bTKZYyvviF4nh9XL0
3z7UDQMKt+B3WJqRxc06sW7Ai2tI37PNmjn3DSvtsQSKnsCVN8ENInDPV60Zk2rH
gyIIHxaSGqwtoZpnB463nE6wZFo/pW864Bzi6mTMGdM191uv9oW1vIxjJVJujbQX
dIEltRQf/TqWCVgbh/cRoKPyVi0MH+Yr8TfZySfVrLT2GAnGJc/vGbk+kyDejtmj
twSZEWS/Hsmm3LaNfC8YAdWPs73tAHZgtxl4Bg5Wp3Yp+wP6NmbHR2dlmliy1Ikc
ToxVssfDf5LcZ6lRSJQaWTDKBfeQe4m3kPxjfjVfghw7GQo04gFxOgRBP+omtUIc
mcDCKGKu+2W7pTSFNBaPVdG4+RPWcpX/x1tuElMTGmelVbgpI1YTW+2tBdvYj4G7
GdQEuwfG5oEfvCH3JtiomB0nxTvWfof8z5rhBsGNIjyuwOZ9Siq46m8cUTW58u2t
V8hFn2wVNjF7p/HfqtiafEnfu0X9i7dAh4yRI+qw9iFcKk4EVk556xZ0fOAexEC5
s61DMJQg15mRJgQv5Jjje28QYpfACuqusbQ6DzpIqM2M4FR13rlkpsu3ZZsMSmwA
T52fSDI8q+P1FAUzXf7SQzFNo66c2eTTphAIyTDonfbEo3PN28yVwbJ95/F9xQ5r
xLXRTfhWbdia27KKPxTShy072nXK9deIxp+ybjUEZjKqRi3A1c0zAvEmymgsqnLM
t/iM6LtOieJUw5B1iumjzh0n6/XBuzF7fjgmg4qMsFqHSk6lZouLcVw0S6GE0lWi
/6M35ajYJaTITvh8i+3cE7MGjIcXfSjJ7qyWayKQeDVB2oqqOzEqZTXSSI9W5qrh
g9Ll1RykAHa+ajWypnzvDwAEphrUO0ZsGAQcFb8fJU9L0Y4ZVtdC+s8ju7IS+551
zSpXPkMSOVUedjoUBY5ckXFToqyIuf9wCrsVFWw3eyPwZHT9qe3PeGRBgw+Z2ORs
8pZ1EUUSLzQrc54jwtESSxlyiJgYq6fgUuozgETWFNnbeD4C3KIOXjzXUez8c2wj
IYTNU60mT+8VeCGnCeol0mXuB8j4A43C600MZYos14Tsa5rSoJSWglSflSVyph/4
DAdkBY2ao31Ol4E2lv2bWSTPoattOsbjfcj1GPdINyebC31Ak8LPLB2n7/NFPOtI
L2Qc13P6ISQwBRkMHHlM3Xhtym4ywQJFyQVBuXC3DyIEKJg9bgYRBWK2GMWQB/uA
4gWu/YOUu1Rrk4uR8C/WWgIq3Nb4CqVKKz5nCFto3tUfHfCsGVKmtjn886Kf4r9l
W07w7a9Ekh05qPOa+tUuGVQ8CAgZIisOukqGogDolwhKigH8cs2Ur4L29xOWTixJ
uhSxjcRt6jiDaf1eM4zFG9lnwZEF27cywh9dPFwdiq6yB1E1oECq3Sycqtrn5gw8
UdaIx9/9LNYkbSvVxGLCPIsuMZg/dBx358ReHCEJbhLYsmwPlLzvwx9MCy9jwL64
MxRrELXp+/PyaPa3NCKlkcff4e6W29N8ULBCnvdS8ahpaXxvU3585wyZRNOH4xNQ
G70GKHQ7w1le6ORmHYOfHA5YPbrDmXupwmmxXtTYPBefDBqBVIURedHEMIE28ePV
xJDJYrX+Jq1Xp9iKGk9PJ/gGxUC6DTQgQ1JXVuGynjvSD/9DjKm7XPHlYrr9Bdqu
8KaOwCxxFUWniWYHK4fYEIN9DhFWWyRHHXAmcmNh4lg9kN47hIZmx80O5gWFsLJr
7Fmy6jI9HVxwL+bkeS4u8t1wxDlQQ/HUAEJPP0frpALZUTQ4AQXK0TMwwVbGjSdC
cL3cUcY93ZahoZTVKt/snI2qscApt0hlIbd48F9htEHeAzUUd/CLr2a7QvUZbUTE
R6domq8l2qFzysj+opcuEU75OGw/3l+MLSd9we30Z78AWRdZYgEgq15kvPpR/zDu
nBU3Nx9z/DImk4qrv0g4DGwQxYfqDoZcshl5T/XexqwJQjiuYspNn/VPyLbXsVZQ
BXWSIYlcmKml+QU6wShaKWAHq9Q44fiqQTXixLSxcRjfW+XB08xiM9xsU7Keo+Ns
nVG4N16gOa73/yXw0BbbvJtPOoaemF60D4Qx4/d9fE6GMtBTELup87RJ+9iZDk//
ed/9AImlrYnc13/QBe4Hk81RV8sa6S6ePXGZeRxcH9VE9bfsB1TeT7wa3ehX9K+d
oRoC3vR2lif92tu7sIR+s/bS7kefwcJU7E6wANFohqWx3d5BnO/AMBiyp5MKl7XM
hX0+0+wps42r+e6dpiJSy8/mq82dKVUuLRagCxz62WBJnIL/BUoh1YlcDAtsiImC
vlUkPIt3dFvqPdm7dgYq6pllvGaKAz+nFEQ22arAqQ4BYPsylFLP+EFhT3FK6hUD
9QY/KF5qf92eOSgWzMlEBiC8okg/PvLLGoFL4B50e3CE3hGTJYQF71YsgfbRG/95
3dx9RIiJv2bcL77EBD0e569oF5YfqsNDDYubTEZFpNtAIRoY8hC8tQvuJUQJrppt
9SuXcXVHZrCe9RTW8LMWxrwLBOpRF7dsDP0z44iJ4uZWkF1qIBOHqYN2OnVzy3nO
7SUSdr48UlJPcwEHxyHwrrzjuoRlVT89mqSPjr6XmGjxrECljOY/aRUOaBhGvhaK
xj6RbS+P8Cmr2XwDIk3/55UsCHJADztQbPEyiaqYsDZFpFEl67Qy0xQV8T8KvnIW
mm/0XuUvnrnEI3PKiNFFXDsKNT5pnJ8OZJmmt/Pr8soX6qQGjVAmEpNTtoij4cqu
Xetu8Y6s3Wd9Z3cxx8bo4cgV5FDZsiv26Ab8fa4GWwxlZEGc9UGvHIga7nQVGyRj
z3McmN4hc6lACBjugM5+YhT9n/4Eowg4InRr+D6xlUrUsSMo+gwhSvijCSuIq+tH
L26fxB8srBN2FNd8E+gEdJXMw+x6l0bMd0e/hPylxa4xtuRJzeyKUdLBDyGTv6iT
oKqx8gOOqCr4ul8Xj8jSiJMh42J6/myWucTCDbg0tXjWM6aXHF+mqssSxjDqhyOo
gltFfpRONXxvQXC2FfYCufGqlBlalMVCejHa+QSWbNldM3RzQI+DDxVIOTmCdhjl
V0XKeKEalJPkux2tjtnvKhxkL1y8ORp5xUYgqmvtzXs68E7DQtRYxMqquIt78d8z
79xgs4J8bSxdPDtq8el+BmKbQ2pjRt/m6c3WrVbdNf3MUWrcNnW2Dys5NLY3e5kQ
jWlA4lBRscoqyfMJW/yDqvFdPVBxr+BBsR3d3RG7GCJSTlBj5C0Ms1D7QC9wyfaO
eiBOdOT8X7PPxc8XxPkc92c8ns2qlh8gvSmaEs01nU4s+U4rnqXhLSOVo68Vltdg
3QAxTJj/PMlEygxBhm9Mdm69FRGvSNs7J2x/L+veqZmHMCDeVn3wffhisoowYfvb
64qaC+tZCcvEPToJ83SC6fhlzJHB0E9dFlr/N4Qwl6oQMURxz1EXoXmBWlEk+Qxf
AvxV8kLzPFXpEsynab1Xb8mSgzcPjiQKAJKugkZhmCC1+Wjh+6EfMIMUGSn3OnGj
cJP687f6XXtJvaysnxTt6VztBC1sbdmiORG4UZq7CmpX2AjN2sDMUdhoxJROPJ+M
zwZRdhkolzPTQ4FUDbY08ZTWpvkNjUxd1rlYZGjHYAvMm3Wqsma1rki0rQNUwcDV
EA3KvHf8hy3R0VovB4OxR2XV+9l1fghKv1sZrr7TJuXjpjDt4yRl2rfBzWIrZPwg
T6UhhtdmhRdGjYSuHcp/keGUHJxTcQSQzEucQSyLjTxqM+/QpYcPLkn3iADvK8Py
5nr5vpWHR8HeExJnzO83viOmET3zJKc7OCR+9/5MDv0/FcKmzSPbjXRDHX4nd7I8
CpBLXYzsPacrW8FsbIDkhR4Kf3dvSo3N3kdBNGzMaAkoBQJNsK/mBN+Df/f4LG+d
qjJDaNpxKcJ/9Onp2kJC8zOow014X7Gz7H7tuorbb/Ieh4ejcUU82/JeXoT0uEaW
DFaqIyKDt1B3y4+lTdd3lPpNRx//FdvwTrPoDinIC1PGydQIZEYE5mNKPdgLXVrt
/Sf1lGLWq7QoS/Zb4spg8/e1WpqUTiwDc3uHQYdvXsLo8Jwb14rJ9cxLYol4MPnE
IaSli5oa4JO2WIcElfOItmwh6kmoBOXxEcLF9OoANOeSYBpxv0EiuiQwoM5bXsS5
TB6HHGebU83Hcy8EiBmknchUyCLut+cT7Y/B5muUxl8A7MojagA/K3eP71ajyD4I
cb+O3SRblywVD4Nm3Qkn7+NSJYEKPAg8sUg/bONletnWNpzQqlIuRI29Dt3lnCWc
2Q0F1TUPqgWHUItTw5KfPluihqsJ//PTMfSy7GMETA+odU7g0T30SfPbP0EjpOgs
7P5CpigkOwLQjDCXa4sPte9K7EdG3H09M7uiwDO5TSHLDHbnkYe+EyzPIusTTYBR
AxODWtyhbfVmyxZByMwN9yffN5GAspoPR9WPIWgGM6Y=
`pragma protect end_protected
