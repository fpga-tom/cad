// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:29 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gApFVRQzu9cCO67Qe9NMHJxySrg1Rq4aqXaQyrvFKYPTWw9zULNEe4dvQ2rLlMUe
2WY0n48HzOtg7gPDvIEYe5AS84Z9gKsF5EGgE6LGcbYTaoCc++MOKfk1tRe+SwEU
iN1SgHY7OcY+ecLWuUXB6GbE17aqFlqB4R7IHCbtST0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9184)
S3NSdx7YFNNwnNigS3ror6amiUMfbxWdf2nMZthtk7G9jTlS+Ifum3suxxLlnzZV
7+w6svHgbxD4Rw2kTzv2UnlcTN3SIPyCYDDmGKlsRfwvKUKHZFOBNY+oYkDR4cm0
wH/KI7mO/gJeUXK4p3y5kuOakXC7rS9VRrKEegEXdbW83mIgayR+eVHX9zoIdCVj
4x8BdRMTng7pGkTbo7WGN1D8ct1vmX73KwOuRG8YzpbSUzuBa+Zh9Yl4ci/u8w0U
SmU2kgXzSQhJD5SERmctBamDo1JhVgmWNap5HCUGWPyvM5R3L5f+h1UHiAaZ+TYZ
an6flooQvPFtpR5ulnsMi/S0nQR5KR8ys7vnb0aAOkOfQDMP9SwI32tC2FDmWkVl
+W72zhLVSwB4SUKfGnzDIGSVfj3FI1ia1f5H7rwJiBEIa/lnq5cKs1ann+N2cxwv
MUguFCtvINorBiPhymbIAgJNGAB5WhCqHdZ3a05v1vqdOyMMyjsBSbohv36vXiKV
E8mI+349JgiZxbZ8+L89D5IOiEGAF1CdHFjsQNAcHtX4NBJvgAqTL8esnEFKLC6B
N61F7n7Uw1dYkCIgAkhFYhst/0Q0lkhgoNekDePMwq62myzSdqCVwpTbyfeSbH7F
rbvCRHG+edhqmwsPHmD7BCXkFUFNAkM9IP8sBu4rYGJNLeKlUkCXFJV48AcnAH/2
326f9HibBMPrIPjHN7SYbMDVs172wbK73tHQRPbkJulC6TeXtbUtLiva8rrwj4VG
ujMPRfssvYdFh3HhcOqWoyoHjGj3eVDi10ln64UsltLC3wEsj9hkOm6DCJ6+516l
P1/rLjphaT4MZ3HLcVRfOkMNSjhWP2aDF06gPeSHM9de4RYCfFltyR2RD4RhToUQ
F4qtRlmq8mTeQifa4xOUqPJIwLlCzyXulK7NO0R1r8pOatJ0n3VavDmjZNyNZsnB
FcbTi+jYKKEmuBqD8IX+jhcq61BDkOx2vEO2sz0KVp91hhTSmsgUki/gGZic7vAR
FHj5j+3AU7KvIclbKImkiCzhNM9onLoRQRZeMhcZErB8LbCruRDwP2mRui+jk6TK
wklGLVfFbDmZi7fnaqSiuEI5F3yxsqaur7MYZk632QZvP9HI5ku1cbsjF2jf5Bsi
G/eHwlzaQa1ZsK5jKT9i08cIjwIe4h9tcm4juEgyMKYMX6OJG2CYTnRoTTLNepT8
hbAlPXnm//lNdvctARDsqQ9sfXA4UPzwFTr5gd3mGKT2CeYjPqG99ehelCF5ujA+
RBLDB/2al0V5GyqUtfQGqB+QBndhVS+5tcRwjU2BkoOeYV5RLu/knXnx3imbdGSJ
M7UV2QTXTsP7gHTE7/Ngx2HxxDdvkW8hRUeUIrs2ss8GB58XxIUYiY/62xHsLhBm
0DUh53n0D3LmZ9cDU8iOu4sFCEPZwdd3+PIU000nUYoSUl7i5fQiWfHwfjEO6wcT
HK75hLqoODK/zbSV4V7yNE554z+Sto8xn94DtLln7Krh2KGTX2QQdwAaq0nNMmcM
pMWdBNlaraJ0D4+KHnOMdyCROl7qu8dcuCRa6Zg+HjivWydU4gPBkpVmXheTqqv5
S8bAyfmyOZ32a2T/7Vy+iOmzaSBa0PNUUUPIx8nz4BOmprlnVxz0zhlVaOWzdvhP
ouG8bebPp5vQp4qvwlilAHYIFeWmLOKaVpkQvBK+x9/kdOOP0wPTzWrq/fOtj9xT
cxuupdWYtGz9dj7rB07JlZlKyl0lPKhfVG9YcjlSfvwzwbQ2h4bAJ0jVEw4CS7If
YgqQsftlJeKFrdUT18B+o+N15Rt7Bgn56OU2Xyt4HK65N5wZ52y83AFQbqmxHd/1
hD1ZPClnFBiRZME7u6NOmPTYPKPe+jOULBKtdMPvMAhuDZneSdmL4XxbnjENIOB5
cZYzGuqdPh5fhBK2b07bieEk2NRJ2ol2xOpVa0hAK/9U/UGGrFWK8yAm2nWvVfRr
OnFu2BVMgDogXbxB6Eche5sb9r3IWi7n46zsktx6IehqXzZP3inAUWmvt2YAdejI
Oh3brFg0QBypE+Vo0Qucjml1hKz7BnDnfTb/6rCW804srXH5ysiqzt8ZIRho2dj3
puXdav7m4jUIYP48sfAyHUxLAyLhT0gHJgKbOVm1ZyNlJypNb9rnhfT7WD6kykF2
FcZigNjwJD4XP+T2u1Btp0UO7qVMS4z6eHKmVNIvXABD2G+ezLMpaLwBjTRWCIOR
7ab5LzVVLtgCnhpoGJO/2mIkRbItmSuD9kmR72j7mdbHGc+PnTFYJVA9d2kDkRif
5LS04G+KJBpD5VHjYsbFv0xHkt9ka2qngXtYzk1QOQ1EPQyonUaS9h9kTwXwWeqM
XghvqQTAmkK0bY/JCk0hGjKstQKACpfRMML6XdSbKqQ6LjDQC6EtcEf1icQt1T3X
OzcovMXlwYe9ftxry5uwgfaciC0mYIjkcrSthHMS4A5ZTVqa2i2KkPH/WDZwUqax
O686mTMTtNJAqiNsPBgxzUxdBeuagtJqf5xT3zjhYTt5urHAtkNmz5HezKjb6piM
08b18Rk1L8+xTZ8J+N8LixVUKHvRVbq0f1SpTAEN3CULP7wBZZC2mdI12AJU1cL9
z+aotYuQjCkXegjLwnTYbh/7AHboAFkJot/jOFVYse0UBpReg6BReUFrvwSoObq0
3sdFpCuQl6nleLLfDhOj2QgPJKS0fIi150qG6TIKj5LsN2dsZDUlZQNZl2f30Ay8
l93TBqdVcK0KQObwApPgIKCoCrViBkFQ7YpfN2o4EZE+yWlWbP2h1pk8hxwNOk2P
rIP4yCcf5m4I9sU6WaxO1MYuIUSDSMj+Gdhb+3z/HNHkAV1+1ip1ZXgMmk1XhQeh
/2aOgoxmZ9Num2OMk2efpqLPWN+xuhNk3B7Jn4tZcXPucWE8rMwJRU2M45JWKY2O
3TzF5WE4IE/YntD4jhNttAqCSfzD0DnB0V9/KUJttbufELv2dDrK4PApy99Q8nNm
1qSPRDwNZCPzdVbkgnLMcQA1EkjsZUYnepD1dnI25aisPYH8LpXvB2ZI75noHfXR
1aTWFlMG+aKnPoIQBPQo0XTR2/m9P0oxHjp4EY/eAO69Dh4mnb2Z6qFZMivXzsXk
ITXbgD3RTuPTntPIGfl0gNHvpLZ3/r73wWZQE12QQxsnUtjgWw1oDyTSAXmD/PQY
OlwoaaUVk6Q53Zz1HJx3n9w4cXl5WOW7P85hHIpXAsw/2wCf+rKXDBYcS4tdkygY
GY3ci6aWU09yYaJiBBn544q4C/mLTnsBHFZYlOcy7BviNxK8fRGf1alXPn2SFHr9
2gUupVKs9GERcac7e/NbBRZaosnFcmgg6dilMoTOG1yxiCJBobukhJg7xFhWN6rQ
j5JlX6vDEm0EcvzuQAzTZV6Fh3WR2ZNH3D/bnXxiM1sFV+RV7OIWbgttPnDeoc4+
4Ha0Uwibm4F8kHTSO5DhrJpUtw7btZPco8Xr0vW+HoUbrsUlRQULiMZfrTWwL+VG
vDHDDTdYD8pm5V1acwFaOAJBBFf8qqeSTXBblxnzQSCSZssMieOprBjYtTx5GGvZ
zw6HRY2xd1vQY+BAxBnqId/361MJPr+ZgP3MuB7/ta8YJO8zeqs83nbdwXM7GDPW
HdcB0AAcdEesOF7ueu2mYD3fUVK43Nft7dgjAAPac4AZ6D0EaqDyPD3B4v5fiBD6
n4WfVGTIgMCJW3H8M3/ozKX9/+G2BiG6ZD2b4cS4F3rmbcZzdM5X/S4ZWU4L/B/p
X8+WUnPyqBLAEWhBROfMo/Kq3LRqxH8FK7qA9jtirTxY9Ec3M9DGhI9MzTpfRLq3
4tt3Ot5I2A5y7RVVzyYsSWHG4rpO0UwRPmMzcvkZplXrQpnD79Jr6AAG1vXat8rU
eH9Xgd6gBQeVy5ths5GfZOEULDOHmgwwSOkBiEMeGniPih+zHJ5DLru8gRV+6642
ii/Se1Q3Zueon/VEOkR6g1jZ8cAJ9yB/PhJN5fbMrkU6VybB+A8wQlMGDFvCwucN
7JTtlnM1f82pcIez9X34z+3ENPa6eWQr1NtsgKs+JUbl8m9GBiKrPuDW3cWQiZ4x
tUZrtiFbcsPh5NSDtupgkhqmXsJqVxKCjpAcy0wDl4ka6QUAkugcQmsCWYc+n9Um
XW4NSiudoRIKopvE2A5Sd30azGGhK6TgMBi9OPUWWMPi5P7+ha8re4BprxSNJyj4
HJ/eWExHXczJeQ2AXeocPfa7BqLnsQrH+4djHzfdDp2+h5P1qZPx6m2EuKPb8ieH
J4BTxl7kLQRowwjCwvW03rPq8sdtC4Rpg3U4empDyPpNAR6ddilsueqlrv2tqJfS
36lbXHmny1SIgvSjKD890+JbX2K12uU4Tmz/NyGd23DfqcUmznWPx+3HS0OVBZPU
avOuSYmLaMErXvmiYBDZrmYzjv57EzGImibOvSSVoClJ9pg2Vg6EdbchenT5OkKO
0Sid0oQGPgvrkguUvw/3in9HbSUrvmNOJB+Rwh8NpidzS9+1h/rhPio1YC4eXQ13
v5rNqY5mx77VxTuXoqZMDOiHz/Wgltgg48bJPkttEA+MzffRc0xg5we2yYM4mdSC
e64nf9k+fwVEfbI7y51waktI4KIMYZMg4bn6udTGq4DF8tcasGouAuCJKxHvkiPA
B+5RHq84nz/MQK7JamiLzU9EHJEXgkphnBj9otNy5QFflqYXSqs/ZTgaJiFBqvI8
XCOkTbnF4/7fsPjzxJYishPJ0IWFFeixYrqEmyXEvMOl3pPF3p+Vr8AGdzi8exJG
d2QyGcNFygXEla+VLgCaDhNhosVELEr+k41OoYXI/N2kh1H4C1p7s/qHXvZsYduD
WDXt+cHpp5frarxXDtVdNMAQK6f6z87cEfNlYJLAJgvEyXfRE7UCYQh4Pa+9Vmyu
deoueottkkh6BCFiHMh/Tsr6ZcF/NWl4PROX05nqN39QbnJVct3J2CQ0qX0HAFnP
2whMwtJTDBjuH1h661o6ORqGlZxnlwlBBwVyHCh6CHgeseHJk23TOVtqAfMipbcc
vuqDqehoDd+Aij/KwkxZrQGWl6J38LpkXq6Mg5Vg7RMxqA+u/BPaSsyOu+VB4k7M
Bg7pSCGXqpIF5OPmgLVGsi29e8H//S81SPyau0kkAI1TzyQjy2IohsR2c3pPi6dT
kxjC/7bVIh9haEn02DE91HD/r4kXdezq5GGnDxTMb7TkTeBg1VKR5lWn/0U+1GP/
s5zszAGLhulF3v9ygdAhjlpeNKt8pgRxfPbJHJgnczCw7pLZP8XKRtVVLS+nPexN
bZMkQBVoKmYlu/v3y+sPCIzeQOqn0kNuX0DXSDaHFtuii0j6F3s4Rqd3WlOL2+hn
yeGvOCsJJVeaJwVufODYlN0W70oXtXgawKpfkrABtDzc7soU5SzLyhX6q04tFUbg
EdJ96TH2r+/UdxluIb8BHIGHgPnPe6+HVf4qKYBS0Ucg2SC4dnywtrytaBoV2NVo
s0ohyWQwciQyUtF2TgEWO1ZDziTWmihLbDi6DkNTH49ykL1tFVzQ3UDfulv+tz+/
KZMwpQAV+9XqMy5Qaq92+6BKXRAWo+OzCtfncBy8mFxPIualNSKBeNp8qHz2KCmW
STJ69F1Nspdl/uxK699gAiMl6nvYRSgpBaYta0fRp87tP7GNDpImvAAq8/BMNAB4
QQmdfYUOdAPINNJh1xi5pRcUxT9Ac71Dhp7/HYIE9DADC61hPqqi1Nh0f0pT1BBq
DyrNfa31AWCVp6+jlfg6EP1AiKrn6eCL6+LaX0Tvb+UmRu4fN83IfHUBcAEpBQxE
D3EJQ4Kr0ZETYF0tUxttGS8cbqNYTwQjGAYAWLjT4RNjbGMbcMBLbAxJ0fnxw2wO
aSWVEgv72d3GhGU0V+5mdNjXwVMh1hzOmFBwipq+smu2T7k4LBchAzsS63VOOOve
OUEe19y58bOcMr1/1EJ4HXJSjBJm1y97VfthLxYvzB5QUhsPYeOO+lcM00gpdp4X
ucLyF3J/xlezlBmiKgKNtE/LbAeUDC2KXSN/V4y421jebQgGzyeZOV3AYV2ty7o1
wIr6gJoMOZ23Vdoaejvbu0IpWF11IUKEPQPLWp9ZxVr/6QxJIcn0teQ2JNco6e3y
PsNGcjcc70NcgtE6kfUPtEELJrf1dMvQtE+2VA5GoNBwXUeiyWM1EwG47rIRHibb
XctQSvoTdMzjywVZo3ZUJkq8zivhYrGK/0zrznHjs46P5S3wDTt1RglO6+GGUzGn
dNslzdph9Fw1EwnIJ4iHKYjecOswQEtoV3TxcPW9d+7wdcrqtRl3vqwzIsEQjq6g
sW0uHpmwaoxwwzm8L7M+hL0zQ245SJ+tHhLpR5xqRM+PGDrG42CP/X7i5v1S0UhF
VPIkVCpRWEe8Z42CFDy9CkUzqIHJclofy2lXxFzJMXEiU4FyzbPvjsiofyK9SSmh
t2sDn/ffyqWTWrmiiY30Jd7NBlb0QAlYUpS3CbO2IJmfnEteR2GgWDV9edSy/aF5
EpK0ISBEdn8EVGGPt0PQE9Qb1FMr6XJiFGPGA/7tfdqySyoJ2R0Z35FdXGGxq4Eq
cZcjamK3enVjt1Uc8aMTSLeyYW18B5LGZRh+jc/+ubP4291EMQYidDm7hlcpmV40
InLhIjD/w5ESm+dL00lRXncAUfpqucYU5WdTIc5IHLgrJdRjl83utGijKgyEqfkl
AxlfdtTvmIxFLAVgHTKphXLh7Ai83A/zAkyJes95aMo1GfC6/dRA9s57+8xAhi10
tKpGtfP3sNd1QhTQ05UF0H4gkScFreC91OxrzZnEQYJ3n2b0LxpmAtH3Uv4rHRPq
JqrW0YRbryzRWn0rL3QT4CS7sBOlKDg2xCoaS7znrSfKh4SK7RQ3631epHCUoSDB
bgenzhoDxFE2EazwdLprPsdTY4ANPTp9q/Hnegj4npYOE7OBEoJkYWha+9R2KzY3
nVhYu6zgovow5DPLbO915RwVrAa26B/04xgssYeROIDWyWVaq/vYW1kaV4kA9qb3
sxMOcq4OqgD1irCpEJBi6U7WbM8NLBN9zbAK1+aB6AmKSpSv6Ou7kHQ0OVxBMPeL
bCpyJv44xsBDUcX9WJmI2J1hAcEbXh+L92omL1jwH7cfbxMcw5UA6pUF064A9/xu
HtljMOH7WNe8FGQoJUdW/O3hUPWi2DEY6+e2Ns+5TebHc/QPtwGzIj03CkuO+08W
vOmxlN9No4i9W8p6Kfrnky0KdPzHnvu5QtfOTgcu6UDH99Nq5tfdm+gK+tyJLcTt
RhHs3ZH5JP+GPZ8h3n9CcQ1EhtKQ2qjpiKUsKKf9pXpwn/dBkQSq4l0r0vVYfpJG
GFxqEtMnubCksnuHsSw4tUb8UpWGDYYnhvHBflcisb1PZiR3Pw2aHBDDvo12siZW
34QaeGGwlhmNRZF3VfHVj2pkkfIG2rwVvMklLXkYv1RY+MLWBXLdAnOrXFQrw87Y
tXoQDnCdaUNjxOdbLICqv5hiwhZc9GOvHiiHeTY/CAa+tll2f5FGlLpipshee3N6
Awr01Br7SE/ckabJZAtQ7fg8Dev7EKbTbYDfSsrBs+0zPjYn76n+Pk2tk76qIJIA
mDO32qpTKsdpHmOJXJoUo4rzxQTcuyVK2ErNABXdQfEU5myQBpM/8sBiEo2Ps+zS
70f/wn6A21b5lnO3XK+BK5hC7NxvuAdAOASU4o/9yYBwsO8tqHdYZnnu073tgHV1
LU4CwK6exjOctt1v1qWhAuBg+JMn2dvFxUYiqzVrvcDKnakIkghOWE61IVR8REpj
8NbvoChqBbRoOxEyCcmOZI9wlP53kqp5LJmvN995MiaMYwWia/nHjZRi6vHI8g44
N2BXYBb2dMKsYZbvSBU3zS4AfhBk1NniVlM39XK+swYBPQwdWeIfev5lU38nkJYd
czKJm848oCUd66yRpeowAHttGWTHI8n9k8PWzwpoMbQp/+akli7Ag0easxrJDWC1
r++IOpC+Ej3bdtKcinOMx/k224z12GXtMN7Adec8NOMOZc7blqjw0msVOW5OatmZ
MAo6VKZpd87r2RJ6hQSGXMe43c0NGY/ERgSOvKibY/dD0dh98ROeQV/Vt/S8YegJ
heTNjTvZCe5Nd3XZdnXH28KdKajw54ib45JMt2TCt1PxpoLolfGnl0IhqdpROmfi
v0d7phH11qljceyMgjhG+4qaOCZAIgdCgAVhEkAZ0E3ero0SLHD9KdgjrxORG/7B
MBpFYZjC3hvCe0P8D+oRiBN7hbJe+fi633LP8vUMT+GwMz+wxky/ogpDsi3gGWRT
mwg/o6J2t5M1gMcKH3wlsmwbq9iICedSGgLAIKg+47VpCPD+kVlLRZsFzEXrMDDG
fcirZIGrwf6UpvWKrX3j31U1aIAkOsAYPy07xlH2YuycbkMXgsjQYlrMGArHTzEY
Ab6MvO3T8agZgniBiLExqQnWMPiyvkjtpzopyLAM1xEQvQ70CqJ4ZDLTyJ5Z/ozN
+EmHv+58fmtUEX45RSUs4XoNGxw8hIxVkI494oQYcs0wC2fzSCRVbSy0o7AvqrDh
2c+0Z+xOMuWDLqk5wu5ey+bpgY9JGhH2ruOfwIqtQsseUzXEvMaMMcuyJ05NdzG9
LUCfd4vV5QzxghcQWblDBYZJ+zPQYdfpr6+PpJTtoC6y1ReexIKhxTbn3J9fJuCg
l+8RVv5f3PlMr0d7PyTNeHkWQzoka4IV4bQgRgg1AjxCfTPqHWKQn4+JfkUUTlP8
dq4HxL2X9h22Dew1Ly7gi0pI7dWrjwchDMMn74UOJivqj0+t7yKthCvlkc86pc4E
TROFVshit7gzRpgBRBSlKesO9YqnBZmIJXS7pHibHpaXzWO2Q53m6UWl4JUi6Ken
fejw9MgkAGdeUA8MhMBYNpLqYnakLXvsL2jW+3/wMS2+ffehe7SyLL3djtO2g0aV
CmELpC6PnfDYdnt+GC/dolxwlEBf1lclH8/tgpynO4bTVQzLUWSktdnHUqx5igwy
wwLEN5yQ2tzFQJlSpenTmfF1wwx3HWOvIHpgKIIs+ffmVM3uhbTHXe7J+WRM/nUA
Q58lGNHFbuDTknwm5XyTboyMuMuK+DG1BlgofOX2fgtNjxErnT2O6CVeWX77SoJ4
bOxQddE9+Esg8aHovEK/Xlwhf1DFY15MF045KkZ9rfpCFJEn9JmPpXv0nATF9y/K
H5qLkabJ5vz/lZIcz8k+tIGNCioN88p6YQHVaFrywL2RSxZafpWNj4JVkzZg0De+
vBmnu7lVzTpR8tCqGL91ME+/R+P+Ac6/J2qgOp195FxR0A3iY7R5e2fZX2pti0YZ
q4abJiXMIE99W9anij2QAG2jZPb4Rt2B/L8MDfU+EzblhOvRO8RKue5unKNO3ORM
djtNeMmRF2pwfu68rUQh5t1P7TlmJmbmtDimEpl4qRS8YHNGGom68CLJsB8lSj9t
f48DQwthNLckEPa5Xu3FyG++1cVtSET2sIIF+e7RU0DVEfjm6yyO+xn/RoWfS9A5
+hArHPuJLjkD5iF0+WibIF+V43upicygWAR/lTn5423JDkh2SDL+QSa8GReDcA0b
mVqVS2fnjpLky3HeAF49rDuiVXvkvFkYGcQl2/FbosrBTFvaa/XsZPZWqIrbDMTd
frjKaD14OR+YRXHtYfNG50HNEfdi7eHfL/tC2AmAcsI8W5tYRmbwIXM/2WFqaKRi
7cLt3rnBmK+TgVjxcxr5TwQllj8zbMIvm5CmSM9c6QlYcDwLKTiCkBuJS/JYFAGK
JvqSH4lN/khn6RbIVovpB55lajDzUsYVB0q92Jq9GEFq79NPFerEAHK1Uo+smNa9
vmKl8XB51TK5FNW2oe2xz0ppCcNrjqLAoOyHbNuYywHvvNx2ue7esT+49G7i9cuJ
Xe6gW7STag1PXdyvSCS70H94CBmmMkcGdgppb80DlynEm8a0OKekpUruDF5en1wi
jgFEXli+7LcCQf9Ry7KLs05yWAgN/8+JEv0gmo6keyaAazwvMKP+xpBIGe0tDMB5
w7//KfeZ2NMdLHz3+x2IHbDknJ/XaYgxQC/A6Qt0VpVON6RHjEEWbrcolR0hKeoG
XKiXM+eJZa8Jn4USRCHb66X21qmm9BXNLxZL1r6jj6sCUL77iEA/jY1BLbd0nlZG
Qa0OSFmuleCaNeRaZ0/Ku3hxRlp15TGDzT9xkRyOTXGYKFEGSJf+NrNP1jAwpRQM
YqnUgVtKkaAFJ58d7H33YIAqRCWGbXsQcP/jt87i9cmRn64ZwgiOF1y5ph9FoIKQ
xTCj0oSwvpuXI086e1Jg0BN7RS5HXcjKW1DBvQYdVy8f53x+Wn6Id4bxNgFt+UaU
AiikI6NCD2TiHFmxy4rIIldX8sOxtXkKs8+KT2WpO87Hee4Hmf7wb1sGJpTsquay
w0P1QEWoZEe3u8UO5HNfx1A8HaYIjS/n09mx6GUwAKnibCIb+wTvlIVWAJcZW+ly
TZZ1taEMqf8D129EqNJnGdOnvlBjl/MHje8niNTkPVjd71K9rHW+hehcgAsX+PC6
BOOsh33oOnQ6ddaJiTrShocDGktMBW7eFucgpvj0H4Zls4jomr/9UTgYhbwF9sYO
9kcusQ/nJpn2CTdE4iZcO32ymlASNim29pZeORqsd5S1/AxlFxIXbsopCYP5iUHl
f/iISJCJltJd/z/6ZAdbjk++o6dULwU0BeMb59+q1GC+kKiQDnUKdD0IVhItGBvi
AX9Wgymji0L4HnyLPNh3Myhb2L8YovKH2JHAXHL0wdN15nmaLoyZzRnf8iwdfoSN
xQx8RNBYBSNfLKO0DP0vLl63ZntNBkrO7usmTw44WpcMNFOfxOPh9jEAeWTSsNUS
+xKK9kNuEgVgo9mq5HBkcvzz77w65Y+/l04B9HG1MK17D2/0GZ4fHjXVnLPdVZqu
imCT/OSUXyn7Ri/8Y+dNUpHPNVGjhJlKwXG9yUVbh2PndP4Vq2ktzEjvHCbRx/nX
X2sPPJEcNm8sQeI5osiul4XkKxf31oEF8KZB+L5iUe8rASE+Xw5y2i3kMFGvriWo
ZARVm/qjNT+yeGTsK2LZp7CASFzMprLd53Ke6qQO5n7rigfgjg1bgQDaUMULIdOM
BMTD/2HFJIi2sOElSi2b9R495dCdO6n2TejZ+9cx+lHOtYn1VJ+Qf+wX7MJDV3Ag
49fkoVNK7KsgKAgQo2OgLkU0SwkDWjVnj8v3yZIVFuVqVFx3aQ7DP+YxF5B9jCP2
YYCz6EofqZYP5170xRN//L9s1RNCvYSvkrbuX/dRLcUlZ0wHChgUmfkkIvYOM3ju
v9Yx2YfRxYKXt+gRiruDLbyXc1HhfjR1VWh/5nuwWpdij20WpMoRrv5lJLj1G7eG
nN9JpFMgPrxRDmqqY49EBnrT0uJnYHQz8/j80x9GaUJ5FopU3yvcnuk50IV4Bp+l
o3XtdM4EqSAtLdKxdEEVnpU61Oy7OSMhXoyZYOL9ZXhi6nBmmysugtfKqtdqHqtI
x1NFjT0rhUUsP25zdlEPwre38vCqFQg3Qe/AKMBhOw6YVWFz2CW34qPwA3QjSnFb
2LgXxKdCRt1MVJQR0F0ydcyBHIFXvMix7xS06I+5VIlOQp/FlLegcX3ZP/WnRgG2
x1V8k7qX71Pnu6iEeq5WXIU/KWalvZrlYyNJLtyrhvzMona2jBtJqOfG+vpaBt7O
RyNRYQlgyinqSXj7siRDhOCF9RU4f35FnXtE43cNcWXwSenwIdbHleeq6NLqi6VO
S9vZ3ahbAddc9fdMv9st9vMEzHiYYCvE8NjHmTlmz+9yEBJWBoq1fgp6ee1kJ+Rg
L9AWwjcXT9hwvRRY0V/O4ZNL3IO3Pa04QJS5kZNjQc9yBbJe7V5cSAluU4KktC0b
jI0jSiUR1BlovfzF03wG08HWtRQVxdCH4OXxmK0WtqmS33ZdUzCfInsioV0L9Z+Y
41tZ8ggsp0pLsffslZVdmqh1SOOu7dRnl0AeM3mrWXU/5TaAfHKi1pdaGaLoMmvC
qzvvQyEGsPrqsxKhZm1EXqDfUmFvflOPPv/1/LQBAe3/OvJgGZ3SJORTKzxPapdo
3blYK9jUp1ANUJPZAQVlbUgO9I7IXgTOjQv+5mSDvPZrlFHyqAz+TocGYMAGSOKZ
Oli9TAJUFR8EPG+MLA1y6ZAsrusIjK43jDUHjmg+np5ZCY3enuUBe3yKUgOZbu/d
cDMI/xf7R0py2E+gOBvYzw==
`pragma protect end_protected
