// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oTCzQ11jofjTC2DyTmcVic0mW1Mlfddmio8PNFTcal2w7Yk92zpQmjVZHtmeKLro
YwmUKbwJj/DB37TP/H3EQNe9zIEj0HUWuhh1D9zDdF6x/ACY99p0UnCXZFUkZYdb
u2LR7NzDnFP2afxO1lMzQJrsE5g8R+Xb4N01xiWICSo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11392)
lD/izibBXMh8DdSrmM0fXXbPjncw3CuOiesnq9LXXq9JnlYoT/GOIELQG7ap4GXS
I3HQb7230OEblk9Zyp68BCaYfuQ8gHZhQw90JQcm/rN7bj1PNx11xD0MI/90OgOK
qNo9F2Ns7JMD8EA6I9lC1ycy/xKTZjS8tFj/nG/1W61W5jEEHnX/lDK3fg99bQ0z
SVnJOnSWI4b0mqVsgtwZi0VRa1onTAg+veAgKKb4TM9sJ0FsfhXqGy8FROU7EHjD
k08enPO1pkwLYBH2qWl1JAOykFsqWO7dQtRE+g7YTfi6wN0zW97NzjG2K5ND/LVN
JAwLmTdkA9AulzBepgAOdW28bosAYruTEEcpaCUBD8HwP+pa4bRTGbvji7C/ARsX
Efglx4RStpkE9Uce8giSPJ6gpxnjMWUucJFkShyKOpRdS7XhXgpJmH5hs6NG1Toz
tJ0G6DO34TT7u4CgjkCmwupTo+stMX+eu6EEzbrqflUUXYYIdKHfPhG0JjFZQw/P
OtQ9ydm6pP42CAT2lknOvfDncTlfROH15gOwWxWYRGkXjYOg/4smTFofE8Op7aQe
tF1WbTiiG9zVCiL7qUi4h0rNvJi4ukW6ZqQJUZk+4AedTkMstTvHKaQ2j4h43WFC
Y8l80bCjSCA2tB098RfJGojP0R1oCQ7PK/EaBMblSHcQrdszixLLkOgsZEe3jzEf
pbPfjcOPyuSYf4taRfnBkitZOCmCsLo0ZG7DvuGgTUbomKQ70gpJXmtU/cPDe9VE
+QXEEF3SsISB14Dj5NvrUWIy59BgzIuuIdJCi/zuLSdq/p12QUUPxI5FFRy/ABi6
WM7JcoWKB7YccLGgIdqFeARmfIXk5qs5pKGf0yBWJa/GhO6XLKFYooJalgrYt/oo
8xG4cn71oVavw9pnd2ZvqJjdyQkQZcgia8xBrLD4gJVRMZG3uHR+v1wzTeH1DvEk
1HbCKm1SQ3c61o6MtIMRQeowsymtX1hLaESBUJxIyWh+KbaWtsWorAZMA2+ur49Z
fG5jJRt3zfA7T1BPzfG0/VCV7MYJpE/yZfLGZHoUggC8c3Iw1Hp+4jQDf0dZScyQ
is1/1ns/4HNSE9QMFGTahPjEcQb/cVzagTU6dMYtXw7DQtPa0n7Bxlk+dtzsYYQc
F5VaDz7QaKQqwxFhCugdfIUJhdMegd3MZg4k5dKIaHs0iHo2cT+tL5mkC1MJqIxC
dnwYD5hUu8qL20hro4HRkZxGus93Kuw2HSjcKKAdkeQpA4FsrymAs4JuPpOARwgp
DvlTTltb6Gtybcv7wwsN2nRw0or3iygv8FJY1ymrkXl2uZoCcUosu7iZKDssHcl7
mQpfLX8jfX0tWPAC5MFv6PwgNGAnkkjE37pvAc7OyQBcYpYYOUpcBTZZENMD64fZ
p4URFsfORSUDLr4mjYdOIh77LHO1YnFwiDleoT33F/a2qUWeHGdXUxN5PfX/Gqyf
9h4/4h+qxwNmaanWGoIFLXAZQuzJ0x2ZmZQ4Zw1CT7KA16mJsFrJLJrOGnN05O7V
r31ojIsPPqH330X5KNE/Q6w7h80g+vJtSQ/1EwWzOm7cP8Ydq9SMQVaN9X/nMkpp
dFZl3zqKYu11qjIzGh9JFkL1bVMPkh93eYClo3vIkNyKcwNV+4dAad28P1tOf+T5
BBSYLsDcIiDXxTtdO0WWdyHoou03a4OTVFxrt0NoWHwwMrHXhOD4JkgIWdHws+wz
pUWymlsrABYHc7goImZfaV4Kl2PP1bG1Bskvj88WgeZ3u1mZEF1Cab8OAD2l1qzT
3zZFNwhnpJcLYtP97EpTQolgy+Jl8u11JXeL7nk2WPCbgraCCbKWZar7Hc4Ut4ho
52IyTwRhy0oEV5AhtMWLBYAksY6tdWC1HVrJwuTkJc6uFHcVBj7sO5ub8C3EXcy3
pte6qy7tleKf9tG0Wo/Dlbnd7FB8baAHo35Fx1QBAC8TA0wqnzo+0mCCt6zS3IMC
VVBGlP3eRf3YFfVcNqmv13dQ/qFoWKsbWOhEKHPhjkAhkTM0DIzEfMAD0dqgAFbq
ssciprIB5vSLBOpUM2+ogH4zu58wPA/GPo19o+5pwt1Pdp7ZFzpFU15UdBSKqxy+
CoYmOwLDiEtz3xW6BQvWHLG1YM2u/TIl3/h77i/QW+zdS4nSex1Pz3klvPZI4HDJ
cB6fOp1GgKI2jISkja71M0AGHqrOHqiU0PQIa5V1l7S7murmscf1ln6SyzLWQ2nE
QzYZQBJ4edz9kkgVBJObVAKOkYCJyLAnl+4NX8WircfhiQZlj6ytqL5BRcIIbCTG
oQoJb5D6T/ZsoSLXWw8Bvn7gla8MIAyrzhBvW7t3Vaf/MHH5lTPAKmdt+pais81/
B7++KUWDhKllTMNSM7xlHewsPodHj6b9f5cy0HvDrfJTMk96fWqp37NMrCCyTfT8
Wt0AMC5UbiL61QUoc9idQ7g46V9K1fFHmUQyygDPMkdiv9A7ifVWyAnZbJ+MYSxS
1J59GFJbzEXdfxRh4DsviBUUH+LILhYD7zTbHVDeiFKXLAoJQBJNRSCE3YrLcctA
jUcMpmutZ0wH5F907aqnOT+q6QXVbvGGL6+FGmqOip06Op3IRILhaLVfIIHIiJ+g
WNlO3WxmPmx8WRxB3uHWSDerHw2IEnMqK2/Pc9v1fJL/glO6Y5miGkkF/BJU9H1F
sxNY/TWLaWzdOOf0cs9fsTzJZCUcRyp5ugwq6SDG6GEmz1ZkIDCrfahxGlaTpY+O
31vLt4t6WsCF+y+tYNNOU7Gjq3hFtV3SPUWMlduKZQoL3tpVSnFBtNjPbNZnnSYj
m7iMY59SXCCQbzb8vWp1n+hxOLwX1y8KoccZdg6ioqOgl3fZZ2kBVMUB1pCOKHgZ
6Z15mQdyCwePmB9y7qN3bePjmgsgk2PuLXsrIjKpfq1SpCbq90VO2R4640/RtLyO
DD2h3VCVi/OC+pCLoGEJaDVSEiuccC7uDcJKT+Awpz80Ghl0CP9MgdVVltA7LJqi
+O3TEtGJB0wnPTkdutVv2MJJk7Vcntm/fSCnnx/XICy//4zR3LVrB0+AnwWdXdBR
BbMYpwJoC9+MFCvNM77YAXXLCLFIytBiUyOmSZXw84g3VVcNm6aalkbQfh3zNgK1
f4eCPbNnTsqfLumCcJQZdiD+R2oqiUOLwPyjjGldUQmSbAwIAWQdfJDSyDwUpRRw
QiHtNgyPksamzLEG1eUxIFof37dGwvMkpT7AbrpWU46ji6nxnhdhWwrrMozk/Ibr
4nB4nAo6glQds0HFX+Yvalu8tmgl6eIeUJI/oyYujSzywRguTL2UqHpBexpdNFPE
VHSulDEcPsToDzRflcVjFMjs+qdESXT9Lw/Xyn/TUdtvtSI1LcNdcPT5RHf47tzD
71ca/72X9rj4Bext4YF/oNE/7jdqj3ushlD4sm7tgTXF6XQJRAgoOrha4HICQdk3
tbctzxcCgBz5GpEDtWUAUTpkm68eZgYugUxmlOZ9U78achixDWky3ndyGPqmbE7T
Q30BqVEacN3wVAxwG3/HCI7l2msu2yPwOatQZxhAJCfn/Lueuc1QD0igpejSP3US
vBsnkcOfhCfTCcT9uVzMmO2Hj6wTRcSwZQ4C1Yy2BvTBfQaYj8pLu75GQz1L14gY
LVX99RwQgJOmgrpxmLa0EomcVeF3m4m0gjKdvy0rYrZcIDOOpjfyYhOBrHBWulTu
6P/917ikUunzAzHdR4H70JkMvntNI+zULcY+7rtySTuLbALsTvpSMUIxcNlZBdzN
qHr8EO1q1AfBqGef7YGj4LnrhVFeUPRqQYHxmKaJkiVq1oMxWx1Q0NeZLnztRiey
pNwbMQy1wAUXNdmoAELbPIw6pTJOE4QKjJDcdukRpgTfzvNn4DBToFCtKjONikh1
W6aZiwJqyJInLEJfSz5xgzvCo6m6oBzwfdl4gDyu/XJUck85Dw+yErKnhQKVNTiP
3nilcou7H7w7f88UzWllsjEZYQMfennc3UdWVFHOsFgDmLvXtyX0durN7ja6Qq2o
CZDQ+4v8vIRQ09ujQNQaeWARyC9XpJpnEO9NOrvud8acko35CAH+fo8HIFN97zPd
qNc2KdaebQzq4lSSUIfMsgrT6UUzTBdRh03eoq6GsNw+JxAcp1B7+wHrZ7nJR1jE
rdyqzav79HpOvWN8sauLwz1RbFpFxmk7sUpeUA6K+ojZRGCmKhxNKmFbBUMYwNyV
9qREmdTnY7UUim75b/xU9BiMFRJMTBtUfCMJ0ngUh11CDxQlfr77kkf4jaeVw5Lg
JNuxnfiVu+Y2nv1ouBafQaZ9/Ykl0Zyi4V8v6W1/C41AAJfgJvhOYcgPeSTKMavc
Bq29YutcynmJe80W2mNfidW5+L4yHKOPnbn52eqa4FMAubkSXYbep+9eUnVjVHZP
lfb8CZ1kNHmPLsoT9tF4OtHg3oVQPwHPZcNNBwhiOSUvd1U7zGKFk9uVzjGBjWXX
gPFx7pguhHpp4HY2rkKLYZhD2phPBVhtRc8g8VzxfKkkB8mgxvE+l6R5iw5ntsDj
xWdWJYnyVgc9RCk05DJviQhfWXY56hiemJBrUzsm++6bT0UxrvBO0e59ppjeSBZf
gr1FGLEgSC8KvR5PB18ETBCPSM8n0+c6pb4pS1LL4vLM5EUa856FbhSlr4fPCaGj
nVDWQgd+AHUd+HrU6CbVaq62LDLyR0TDLTzjlV0eL4S/p+lf9rTZ1fjkkITZlZKu
DY4Wo5UHxEe+c426mZnKM8p1jbvi9m70g1MHHHTVQeVJ4ckuo8W57qT6oJaOIybL
HP/zod6R50nWkwGjo1v+s2PT1bNnl8dmQoVzufjhdWZeRZTjVK4Y7rfBOzKz09oo
KksO8RL5qtiYGT4AvJFXH4GTJ5S4YgfxuPrfB5ZqaHyWiOr7Bjf9nZhnGxhrz4qM
5+co/WpSRI8jrGRNEujUCFg+DmqSn4KLjWUEGIr0iHYlHFvEa6KJ2QBDktnw3rNw
GovpoE0zcVt/igdKXf7d4/vh8MdSneWQN2FDlpXTP3im1pllMgnDyv//zf7F7/+m
AOX2eozWyijrMG5bEjuW8zB+Nmt65sBXl3GVFZZ+yWEbx1wIXTDU9wu+baT84ZGy
06csR+QCJ5fuDgV6D2mevF21QagYNM+ExuYm5fdcTwvDYQwDHlxm/Ag3zIM+Z+kr
R4uWPMsNGc82nbdiWRaog13NRR87Tf+vrdmM6yIyAVXtpIS4hLbb5uJHoc5Zkt7b
wFahfQS3LNBD3vmcFHRCeYe3ZFGTnoCHNSMStRIDkwJCWxyoZNwOGkKd52Szmgg1
AWexXvRL43q3pD1MLs16ooIWo4+wJVQcFIL/elb1CJqhfq88B07yjdntGWi5Qjwq
DfEKOwQEXqt/FnRG9UPdHSPSwQhzsSvkniqikk361d2cQogSh1MxnfSwZSM7YDI/
If4SFAGJBh3BNUGEFQx4yuhaiuMYvIDZHUP3dMyqlEY9QbkD//VvfYKOYjM62cxk
ngjQdS8SWG3r1XACp2Ib3yt3YuMyECrSI+hTpUl57Y3hua0LV6Zth7ov2deHuFH3
8NaCXWKt7l+3oyWOpn5+74zaRsnhLOUTGSiy6eYAlnKZr6fI0ccnaZUIbAuJCPYZ
21h2dS5kP3QjRyy9J1+CyFcjJdWbEifUSg5fH3cppqbbh708hegXANoIOUTiHzue
uFCxRxKrBiruNEi/nwtNqMeXMrLSxLCqWNwShJx2RafDdrbGA6cOGfMXOfBNm5Mp
mntqqKfDbC6BwAuc4aQQOO2XAOZJTZiukUddjWsEZLqEEEpcZFNWMDItOIYhsRjP
mNUnZjva+hjRd8sdd2Z2DaU0jeewsXBi0jiaATJfUJOt31tXqJISgcxScmwRSUbL
5ClbbZZcs5liNwIjJif84MDMiKxYqWNgo90ngRWK0RZhGz+AK/vsFuHjbbyuwYUL
6q9CHtkuhr7oZZcHzC5np98uve5NHX2ErTFCGKVn0WfNdmqvZ4Llzsjva2kwIVa9
Gp+FXS0EuI44u2bsutem9ZmbsfyooD1ZNcj9WgcINt6YlrPK2ZVXtRTLUXkJAfku
l+9Y8OQ9s1pm5tVKz6S+E1pCaC6ud48XbHTr4epV8yK/tSsmtH0YrpDHBfdgS/4J
spusHhp+DPAYFcoD4vsVD8wq/iXHq8vVbw3+tKGmYo02m+kzzUGrnlE5kPku0y72
tzBxvT+/QqFisvG+7AlL/bh6pWlC3m28Qch/YjZXyMl2hqmsXol2WrYc/PuKJLqs
3BXHLBH4F6t+haXR2572Tveh2Z/Yhh38pvKlg12FCD7GpjtoEMDqdhv2YW/7ZqKY
gIlb9tw+/hZzY6FLCIhAI+bHqTg5OxRpivdm/Vz0gMWHRlC0Bw05gUsgwp6IoJPD
1Dx69pR4ESiM1X1s76DImf7zmu2OMiR1R72VaC9Pip3HycNgLPH0dQMRtbdy45gL
dFd2jfun2rHbc1aS5tdRYF+dl8qr44K+lIx+6oWwtvCPUCwEjJRHtpRffP52JluH
6lcIk5+QnxQiySqCp3HHvcFuBZUbb4aKS9w7M2bIyvqqFaVuG8bXUS+law9zRWV6
th6gRDh/iCRDKqshTTQxCP+Wp97FtQdQnDaAJDJC2eoyWyLj8Lh4lUIpBZD5eEIK
Oi9jgAm7ZOwbEE5kFrxqoyLb5w0eFH6g7DunjIgDjHErWWhMQrzeg9QO5MALXZS+
RfFieJdL1d6pNzcomNIffxha6f89zUsKnFrrPeYrOF0pCVCH7qRX/mh4NN1mlWSO
SuonuenBfM5k35Giw5L9eEwakhIUJWuNYcxVruPgqeXDffhf6OZywUtwMUHebBvy
6T89RQMpYmCdvRDt4tqHzTKWuZ1P1qkm3PbSx6+ELlQT9x7g9IAwdfU/FRfJQr3N
332P+Q9n06zAPRVEW86vSS0f/DjUwfuDiHLyFnM7DdInX/wbDk8vj668QSTXXMmn
8F7Ik44+ZEoigq7GWvGq3Hx5zCMfERsDmi685nztF2VLwg4OcpDmy8+TXCBsEGoh
hlln9Hqfk6xY3Aq1UwXBpSQrGyyNGPVftTpfa+54+6bK7Nz0lbxfetqppbDiaxem
oysHWoIfr8a4USOmNLC34ym/O80gV6Z1r5DF2PASelEozIgFbV32pHX+3c4Yl4t5
+58+U8SugOF4bAxjpaohnebCxJjTzHID5l/VsQwpC22uNe1Nk07Ajco8bd6ff9rf
oQeSOwb9m4KdtD2FLSQMSQOLVN7qKk9iBgVE7LSjwkA0plqXDc869jQHBGrSxKCh
1IVQ5kStfkzINXc6v0EnYUReieprM9hfGU3s4/Q8EbpG49aFZ0b2ATT75B2liM+j
ekf/AcA/59gzua2cuT8aiuebLQUJsGQw8dhmMmJSOJ6hgKt9APKXgEWGiLG7wwr9
Zz+eNHDmn65qh1BBPr8y2phoMBnI1+/YyMQk9iM/H3iTLux65uvfI0xR75B7va9n
QeuAs1eFC42ScQpuqzSVuirKMAFW784N1hHAcMhrPQWGlFtDlolKM72VlnCvjnAD
mXYVMqMk+f7JiZUZ+KYOtjbfwzjck5pt5QuLdlJcWOcjs4Ba+tYZo5dBJ5bt9AB3
R42yYlFfM/wjKitGUm0/bA/6YiZ0liCa8dv4+wdxDATx1oLYCocWGGH8Yi5J3hxk
kVU5i1kKFskOuQ9ZiXwl41EgEc/cWRBmNLC/DNP+P3zUYPqZn/GNdyuA6tuv5NWq
HHu9DRdRoI42wyzcW6xultcQcFuOT+eoH5DH8RTgEtDqLAbBNYPee/usAtDc7k7n
0kpGTLrOTG7jlcX5GrExxyV7iNKRW0l2q5deMQ1yIIgZZCMPFf94/yOhq5rzhEaV
UCMdJ+vL1WwNCvEwrVCcieuKbVaei43E8arCzTNV/SXBfM32j/7Lr4qNkLA+F9Py
GM2YS/rSZnqrz/prtWnNvbfKtn+JhHJbaxzdWMNf4xdW7sSvw+EEndFzLJSaz4Ib
u3gZNkW64GYh24WaE+7B8x8/q1+eb2mq4qsUj47tjSiGRc9/l+/RFfaaoIYvYsJj
KYdJAyRzFUF3ULGkrIMYISwGaP9Jcf25saYX7XKbVJXGmfh6pb3d8D7lYX6z1M8r
SfgsTo/bpDLiIR+z+4Ge9E6Gq4JefbBuEBj0YDVhXGFvBk0RUEf3PQ4lhf6We2Am
lBs/gE3Eh7xqu2QHyYDRx1Gbun4tI4llR00+K8l/cIJHMxgal9xQtmEDya31TohE
j0d7hCYkMcr3I/h+ibcToZGuQ0J6LjZ9ldx7HSFPhETs6kgmN/7+t16reUmaYjHs
3NKsObMI05OlXiLyCQWlsTENym+UV3vEvn154q/s2lASkmTq0WpgkvFy04RJvTKq
rxwGcREQhvHfRAe/uVS3mkTQhIkdXZoAqi0KKy5wd1N79PzDjeBewycthrWA0k1a
sLwaDBTEtZtU7pTGEknOnmQOLEGBQjCOC9kbaJ3SpYrWaS8I/yef0Mn44nlrLANP
hdzC6NR9CDLHYXft1743t0qLGqF+Dgy46EjLzPv/jfIRPh7180fUoT1c68cuNImE
KE6XWsPGJ+GvgFyPPHGgplMV8ZDom2OsSgVdXrVdwo1XLGw+lqS/1V7b8cG+g3g5
TdY3UtueBGQfVhuW/dV99gYq8np7/LMu9ZGw5xEUhVTzDq9M8pQUFLduiRH3L7Qz
aF5KhA4S+OazekB+OPGIPYXln61/Tiwa2/DBWA4DOA7zMg1N6UWKussoP4RTIe4V
honwTiAZkdjAesYowAE6552M6YIgyy0tNZTOrZL/PbPtjDAmUCoJ/LBK9uuHPpEn
GhIlzPgc6W2axzsMojKJCdEkmg13gpxqkbOSOF/CWPRu70ZEuJe1CQoNr5bmNbCr
deMSzLrbLGV4mARFHn1gK9780lP0zaIXEGJfyPXkEg+m1HhWQDuMbkpjgoP8rDaJ
fYXSv+gqQ4A7WRKtgKLN4AVXLziRvJcxJ0iO1gIl+oKpRrKWWUwn3uyQsbP5rZs3
8WQIV0fISgWsgQbkSoblnQED8qiye4TO3plmySKAvQWTzc4Ey21hg4zjnVBTaX4W
20CkaYLVRBQ44oAS6r/D3xU/T92XSG5OfwNPuDoE3bWjz7BkmwdbNKDS3JDFO2If
j/4dky+dmQhro08WaEKFDV08nBcMtZqhMV0c6+GM+znjMtRJ0ZIkQU/ygnCfRLlp
C+w5TKRhO54mZcAxR3MjdGSBcmrtj2cO2CBN8/pjGwbyw81mae6pB+2O8eTtDZrD
SQPXd8fbqxWgkBnaR8tTw8ZH1wTFv2Nz5eVhjFZGufzNGFatDdxcqVsrCdoT5PKZ
1QxgWhhL6KIvAIZGNuQvvOI6hQCzZWc0zBAdQWN65IFKRH+M8qCgRKyKoDBh1ADh
BHRZKu33AJIGxgPPEhnq+vv9pihefSCumfp5wP82g5FGhXAqBa3q6wfE5UgIYOB4
z3X5ywUirh1HnRB+6qJwHJDj7Hk/nU+TdQviUoG6fEePyBGrtn2z2OUSJvdIgton
uVuLRs40wiqguNadr99c1/XFODRk1zs5CHMiNqo5In1foiA2Ffl04woQ4+tz0nkR
angLNPEBcRnS9n/yj+wCNEs3FQWf8DY7PWlfPuBqsIfRWARMXZN8RCl6OzamBb5z
eRrNiVtVoIuHtHhHxnGbtd3Q5kLmtO0sOURKy4lZ3V3WJ2XXikfw2qbwryzUl9nX
f9ASyxGydiQKZT9LtMKV5poeooeBT05gs8R8+/FRhEuzgFdHnWdMLIkReJu1q/81
y8OTERRk8yH2t9+EYVYLEZZSNcCWs+qkmmu3OocjuAGtjI2TQwQgoJEaHBaS0SG9
zQ6j94mpXdmGK5lhBaI47+ddoatNt8rh57suFfCo+BFfLr0VMUIdy0n97+7cHucX
Q39Kn3gUeXOFFAwsnknGTCJCIewfjkD9IS9LpRc2h2UBv25YBGQs9dsubUy3HG93
G3DNbSOYfWRidDrlw8lGAkXaBCagxkKzzN1eSQnbspjdUcTsOPjagzJxSEDTPnuv
meA71TQDps+Y+vxG7bBV6ot/5P4wAECE5B8m9VURrxBxaSxx9kXx7zpoLDfbLgxz
GOltqkA0x0u/F/pTcD8EHyaon1aUWnbUM/epr2urN6yxYyko0H1JbEqaLN3i7uo7
vUlwGv6/qISHleuJy5SKcpvvsoXbhEbImB9fsRHT/ilPSNbQYPXFmhA6NaiTv6uU
HM4fppkIGRu5+i7Pvlkp6TageYNhA5VtS391YlsZnYDFxzroHEiPp4ZFTGftOH0P
c/bSHZHgVb1+rUHnGmIcuzd7ImCIuABosEUCDl923WoXZcNUSBZnRMNKUhf3UH5V
q8E5pFZg+THoJrepbLIyP1DYQOz8XUvWwBh1893Fb10Tr7igv25XBq1VtscGPaBF
mps91TrYhO52g4YuP7ZmlPPXX9VrIIbzlEXWKSURTvH1AuC3LrVw7EcdkZdO3hfn
K9ZBdZdSKRj1ZpnKJksYGRSMXNuVMOu2L2GW8EAEtWIer7TeGgLXGzVXG5S6G5BO
EE+y8SbkFCMRT0md2s56w/T19szPwM3DIPtGeZvR3Q9HAsbBSOF7nJISm1lcOPQx
mtGBpIs0yvHd9yhErdMUZd3RuZOy5JtuYyxLWDDUkqUg0lydIGFfD+KqRXJYzXOm
XC1ww6jwbPslpnCmEKpJQYsIMmS4vWegUsMdsz37QzZ+Bs6oEQ3da6WXoCE8+e8/
fZ8EzxIrHz1u4x3uUcvv1iN7Iv6eTG5OT8u3ihvojF28+c3IFENtJmRNfnlUDgl4
e96/0518nDXIIf8po97ZQWheyPrDB4Ya4cLsnLUWSP0JoRS9aZNsMO9MiJg+a+yU
RrtCB0Hyme2g5rK8YRS1ANxijeHTqExeAB/EDDd1MQjXiFwynxoSQdvJPtOXReuk
k66aUGR5ujv4kUzhoTygVWohZkL5tWst0ifkPscniEcIpxAf97ZGHDdM3xfqyWXE
p1ExB4ugOQmjhJON0btmVyh+G1X8p9g8smUHBpd/q2xQm2VOtQbmqaNorv8IU523
rSrbwvDsNeBEH7UzyGTsbzzpcw42JNMrPhrUN59hlqAehb6rP0TFuVS0QO+aPM24
tZpuJbThWrdxt6N3SL8QacO6JLczPeFKhKb6hQLVdlo2yrPpdnh1NEVhohdJfBc8
Ocy0aAkPuwL9AuOPpuJaylMoXHyLFrzcFfTWMAYgqSPciA7jyh+Caz98nGi6CXst
w6L+987080jeHOxk9Gg0hI/EOpq3ephoVkZuq2jgNbvwcVfDYCn0RK1S+i0JIDD5
+d750xYz9hufxdleRfj+VArxq+BpfxB/pGsAClG4GdONEAx0kaXcj+3XCGqOALrY
M982iGIDGgCsoe904E53FlXy3FiHXjiRUw3LPYEl8FKUR1xOJVF3BxHeHZCvgx5k
88oTIXcD9/aWvHnjzJ30r2k0Qs3jW27axBL2viFQG28+dDnGXKQBrRByrLiZHmB1
8izat0ZFc+nxfW5uRPix4KhQiC+Z9t8T/WvhK2t610166LsWpO3Nn2McqqI9HdZu
ue6ysUReuuLcknP+yogucw+NKE7B3+d8e2AbB8j6nqq+Mhgq6qMnDZpmI7EF6af4
rVpRVaeILJzCXSpTy7upWuXZ+Zr7MQJ1bwAI+laRC8r7ZcLdia2NOFbpEtRL9J45
A8rquRy/1X7UaDT4srKvWHcEiQUbKEsBajDd51z4QzS0C3/5vaM2vRGLVfR/lJ8x
eVL2X+5+Yfkl0x6TqpvxiIsSC+lLlJEwsA+H6q4Ji5dQnTozXcrtrRYgovthkjo1
dlZXVn17xGO+4kaEwdoAShbb2BfAVM0WGWS1dtwH9UF7qX1ogV38KmOOyQU2zi3n
ANwcR41De1qpNr7oVE+95cfwnRGDSXeWLCueDB7jOTsnqwUyGX9jsSFKjNo50gjX
n+9p/IlNT4sxbbwGjSykhp35j24G+IzSG8SlAlpyO/S7JGH/pvQcS05jf7u/MGhG
bcoxBG/4ugA3vs2REbwilvk7V3pQfkHGjaBcbA33xN3RR5uECyq/vXzzM9bd45hr
yibIoh5JUXNd5B60DOgl9oRG7vntJ6NqJw4MekHASmFt5hUob1F1AsPc3HNfWTJL
RgwQWt5VKmU5tcQVGJqJzXU9+eJrPCIHQTzQgUmmv0O6bNfRxSbl15mgDf6sAYYB
2ex/6sUh350EqZ2m+Ye4F2yDPEfkwxUW6WDGFuBX1vsi1na4pyhRnJfmuNBe/sK3
atw0xGS8AYhrRyPAWrbbeN7cfz6+Ay3WX7qxSjITLFPjmFwL7lNE9Sp0fI0AtdtX
6ZZEdBxrBqCkcmziEfJMYhQiC4yqveG2M7Al96VCb1VmeFpnRtT7eCabCURXZhv6
R78G4em2u9geSoGmce8pzS6RbKa2EiSmVp+KTssdGxlCa1tkK8H7zpCitrUikCSB
Y1ALvYBzPsVuAXBPeYFkaCloaaHN86R/ixqJnsQF9e37ZbCGLEKI0XLOBXJyFr75
mUjOM4ixgIfukyQHpV7uzcFu6i1plxrGr9hckdkxfoD2j6fU14iWz6IXK1s44oYQ
sPhL/foEC0j7TUv0fs0xqid5kwjmzJqnzcaBHHS9/FF7Be6kw5Pcp8jERJ3XlCJk
+qeGNmOynisZwOL4Lw6lSuYVqU0VXdPjYTQCpGsq42SAsPjgW5AmshwMAc2Vst2z
3DOvzYSB5p+pfTXC3ypYUMfdkBd4g6NZQNnoGVR2GDUEgfsqSYHZjKHMkfjo2+Jy
jf/Yrxif+dNBVZ1reADbCTD3jScK5dKQw29R88XwNNyCYlTfenXiA1/NC+xQ+DqL
XqhxkZ6D619MFYxF6MTyPm0e1iw7UrIy9gfVUziZnYpvCpfyU8Vnqfkh+f/iKU+e
cSy4iSPFmM29Ic5Wx+b9iVX8So8mNQmqUGfbclLm8cU4UrgJPpIp6+gb6NXHhrrD
q8Te96pi0N+hlNzl2P701kdmOQE+L64OD3RojIVL0Fm8q6fp8Rcpob2bl1mox5vG
WdgFZxDQ6ZeJPL3uNT80Cf8bYw0elZ2qw+wmuHZBxAYzBYYrIGPdlNuStpFM6GxY
cKCU8ayK0FjltQlCtos4mWmlEn2pGjvU2lV5MhlWOnj65uVNvQhX0RmV7CnMnuA4
ZyoRKZHnbtnfp6jjywhQZPWozItSqYU80MRwj9r/RdFs3tOTqlmw4wb51c4oJmyR
O3yg7CIpzy3BGAMJgx4BBn136HzMzAVfKLOJNZkXq6CDwPVXKUXr6zWqUPA2NF5v
ppW1blDroWY7iF2xym1LpCU+ltP8lwge7bDTtrlQheZJqEQhjnMHNdqMEoT26Pl5
cn91+ID/oDDZHuN2d+lgDa1uIIv8wL8WGXaznRi8quu0rJaa0Ywm70UBC5Nnfyvt
l8BT1njRLfKpUT2fDMYm1heXpAdSHSdFnd4uk2zin+0TSb1y+JAeaPI+GumdiPPs
uPZ6Uex32ZALgojQiTcvIdpq+sVHeBwdTZfhVi/DrCWvH0Anz2ossanBKP2ZVeJi
qNOgzq/11VYzcLE2W8UbKOAL8i7yhQXWlfia2/nyiDHFhKTIxIwAUoj1zahCPZpL
skIY+mnHdAHCWUGYyPnqkteLeW/erDH7M96qpUVLq+DBaXatc2npr8xFk5GAXWxO
TYh+GV/iwAGUYc9qxAFdo6GoUq+zdt1BqrnBJbdwK/zYGPJ0C3LrQwdNz7bwZaKm
L9J53gzO3s539FxadZFKeoPRBoYYN6Ciz4NUB+xaiIGwML6rz48iK509nyOW56en
iPq0LmWxq+dTYh/nsn2OjThJ9myln+trE/z9fzXm9xYAfSTA0+HtF/CnxIyf9mwc
Z8tGZn/SYJZkq5R5UhAxFD12zyDv3zz4QL25qKtiqRwTEiqvhDRgtNPK7eX7gdME
O2aZF0jlVxrauZBaNVw540DHF3iISuBh9T2J6GbVpk8pgl8/d8PurnvaBg4vQWRA
AZ3tVtDPtbP0qcxb4wdq1sYM7fbhn0KoHm0UV9q7g6tmwU5bCa3yDVd9SGAQAA4n
NjvLt9uQLGvgxV7XTTQ/aJ+DM2mjmqM4QX+PIQailLtYYrPxdnbNEaJ/9AFIzCbE
uTWBfjjdH5ac1t1dgeygbKzcL9zk9MwOlLgO10prlY3+wB6pABidJpm0/k1Z95jw
19qqAAda3olsZARdIRMnwawbfh+/zDeijT6yDtUi49nH0I0rHFvvGLLFQsD2gE76
E9UX0XH1KYYjlxrrF9KM/N/m82HO51KNW1cOD1Zy7FAedY83XMKY6sR19yZjoJq9
0kr7NehOaZ8xBqc/t6sbwA/n9RTmMbPQg9g0axTFStfeoAkl9rxOQ+hCygT2IJ4Y
7S2upSY+xA0eYPtf7IXBSK+6WaxEXxlc0Ozkvm/pvDWRwn6APJ2qYwnf76PTtF3r
7hnjVhMdEDa5EINu1odVgvg//2CrfhiccJXDWykcjEDtMNwcDE7kPiyPhTInWUaT
ArabjzV2AvOQ9bFuLdfHLYVmGWTrXr7Tox2jOd6I65ZEEvxYKEdvGJx/vz1lW3qc
UPogtH0n3FvwDPpz5Qqd3uAgusgfNpbN+apUAfyn+mr0ptvifCWxxid+4jO+M4Bc
cq87y46LPl5RHmsOE+DnH3s/BM2CzrXF7px9DSiQJBvdBC9D8392rqlbpo2JTe8V
zfnm0v2mt9+wYJq0YmdV0O2imYobwupfg/qTFIXS5FL23E7pp+L21aKSzQeceo5b
HYqPntzDyNnuMRjb7b+RHQ+CUT/eLkfRjYxikU3TXZidFahtv54tqh5qH1Ey17s0
ZaYPSTZcmGpJPxWz70XmlaMcnQYKnHxqf5ubvN0nfnpzXi0co7oKUTqfoSvanSDD
zTLxXt/ZFXUxZq+31M58pIdrtgL74EXCc62pg5r0JQsabCEMw6pj7pavATkUTFIA
fdki2Ush8FKsOqKneTG680hZi2HUnDJ/QArkXx1o0mfmHxumzedWBrB5oJ4MkNfL
gWPlUuQ0vYvbWB9PA2+H09ICyLkODRp5Yedjl9YTJOB3SLbUKGyDX0V+LflFrVVA
z1kyivbKfl3Vm4xB1+lGO4kFHzH9QYxQ3l5z7nkJ+P7ZW1oKsqbMB3rY3OwKr84z
SG5zl1cli/2qk9FO/cpagw==
`pragma protect end_protected
