// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
efGPHowwSYWNGWfOJ79SpmMteyAGziWU3g6HFZ6gJeoBr0APWrqUfIGRVy+LZI5B
UDwKeNle1ngjxM1V21Io2wl57OY6U9ZeW1nTfAw1Eo1R7jDVdgagDOYAVkGRhV2a
/+IABAkEPaSKjvyFh85V3CnRpPNWsdb/uD+0KnzN588=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15888)
BL3M8nIjLWPldHXAZtDYu2PLEFHrYHPXLoYKBTldBm+yMYvtV9hCH2IBObVSJvVz
9A59llSJpH8lA7IUjtJBC4wMGNZzxoZo5EEX6NUktDronJhQV+NxOB1s6CNtfr2i
uBixScqKcxHkMARUd/QwFolZQ4nI6m0RXmzbiMw814YIQqcqHJavf0EhRS3q7NJ3
8py1ZPoaHj9TJjbfYvTm898tw8HVaqB4wGkI/BZQhaaSPB0sFaMMm5Kb6brysEhW
1p4Ix3yZjnFqxVHo7tVa/XVqEGnAlBIjiExMkcHi9v/TW4P1+iAOiQujZaVKUfV1
dIvDFGr1wzXTMwC1dW7VuKfcBb6NJoRBAT2/pGcZmt/QGNBBpZ9SP58vY6o0dETD
Nw6nhTYpAE6ZnQctWmLE5CPigziAgB6yBpNaVvXCTgGH5kwmmFCFIiAXR+C9Jucj
B3XN5W+9zKHX/9txnNlXLtjgoqx3ht/XvkzRAaFMpW+LFKLpWQp7xv9Qwa0Wl3q1
H8hgRaRyLugu/YWP4+fQtaNJGxVm+ZMXicCIyOWqxdQ9ecYLiJ/CoSynlWG2GhIu
UBMls84wDvwrSdtnOo/hwp6xcDYucjOBJZwfOduTTyvMUwJOEC+ZNQgj2YWMudm3
MuKnpT2ddqe1ilbWc8/+Vl+xbFXfYWlwKXIOLK+RPipyfO6hJ9KYet+jRedT3Kcx
50pXfjG47oLCdCDHOTVNiWItN7V5IzSYNPw0/gwNtXxzxlXBJzb+MZJWX7ipVw9L
JyULQ2oXOwsu4QcVz/1L4JwEH5ObTIxUGEa5ESSi0MOmq9yeJRo5zJkhtEKrX79J
mm9JJ+bMcuFU64QunhKSKxTJ7KkrVWKY0Y178GdQN4/w7k1STnKGCFwHluSjt+CE
LbVUig7tXv+lt3G+pIvf+7eSZxsqXO8pWXnEPNQBoJG2gZxgIr7ko4s9NsoEe19A
zRa2GLcK0tro5KRimb/Cct0vaSaL7+w9Ofv/E9EctqHA3dXvDn3e+koGuiwBwOUG
GhT8gEe1epgbApUtlqtP2NraVmtutOxDVOqJTan4razJLTtzBuysD+QthqXBcb8g
wJsuh3oJ2xgu1LtJaRvQgftIFbt/+0XzXOiAQoL+XYgE/BP1OIqQv1qB2JWufOG0
rOhJkZptXBbU9mQPSsf6e402KYif+1aK1Gb9ezUaiLlBJHIFvHxUa1xPqIfNb5UF
vkhH/+r+w3nZOMvBi1z9HCyVnntGvU39UeyYuBIHI9Te9oHsZ6PaNX2Qnto19488
1wNm9Hooe0NHH5m1YufbRouPjqI4jvcYGe3B8OKVAsnKu+KtXMCD0YAZDWS4RFRZ
E3BBrV0DUDVGDHeBHLjwc/vVH70CERSUm/ew50FFclmRDE5a+bsUQDqnW72lstkX
McH9BnlUBzR+56YSK9XYlNhK/5DcPFO5HjpZxc4iUVFmRPCTjkjfgr3GO0RasS80
kqiSl6FDbzxSbmWfOrQpLDLvVNSTShZ7c2HLA+7hboNVFXYoYFfIthc6/1Ptt1ae
VreIfHp2cxjf/7RHFgHmDGpg0elsABJ+gdHtzbmwxtwg6gzedwDJ+Zah7Bhtryl7
Ml8Mk7D82wP34Qeee3e/bbGJo1GOuRihutro+hg3LgT8wVKqsq96VqW+pynXmGDI
ErAw+wM1J7Q90IlNkZ48hrj6E+I94fxYp9nx+eQ7qa7PDQpTu8IuufR1KXwFt1Ua
a5UuQ8sSsvdAQ0oHpZt0KYjRS3UtdMBE7+kp49fvNTv0FZbkcLuEvS+AlRYiS9nx
zpRAhKA2dfTMFHIy9BT6yLB69gC7q7jGeszg1WbjpBzc0q9t15GnharSPAU7QkFK
qiYm+WyLHaO/VnIZXnQA9jkclMAhqopUb8l/ALiBAD/mSsY8kG/DN5lkBtEoLvBs
KgfpOiqfCB7nRwDCxVL5lFTGqM1Bsop8GSq431TwD+mO+SHSbbU1g4jEmEEhNwVt
O5CavC/s3oNi6UcWl+MN8Sqh+EK0laq/zdq3R6vutkdTdi7roAXU81TQhxeL0rdz
JvUtY91tujKoOSfPHRCjOO1O/rS39uFDnOfEcN/20xonZVmBTRBjVI3h/DQIWXGs
0YZs6e1HfUfuVNos5oknTWLMfv1U0+PnRsQKelaEs/pAaqLdu2EvrS9NcT2RKC8O
w2D8cYtOih3DM26mEH2WygPaakiWydpRlLKmdl2MXiZmRx+gF5Wo/QIQYJOCTRlK
itsXuSXKJYK8FAM+xLl+neI05IbFY+Tu5v1bE3GZwF6fWPhbleSui24EaMiQc/H/
YkJdwXXDktiaITuddUcIkskwMxKhZ+SqJFs/WjwcTLvfEj3nGhBYCNZZuHNxidEz
SZUNp/YWRdj/OSLU5FkGQzkVxICRAXLl1+mJ/5y6PJzuC/HXNOpO43IGy7V/2DKZ
mf0q8kTDpPut3H9FrZ0gIUNWOo0qmBPeG5g9HdtkoUWXqT8GljMJozMDOKRAsFDj
QfQ7xwlUT/KG43KgVKruYV42/2F3BQdyG6KKCEUgWhAte/HMidkl7qABkiavUNey
Uy2WCz5jBAf4a8TtRPgZWOXMKbrmtYFB3AlLojYRNQ/ORht39Z0uYemdhnygdkhE
8V5PzakG4hF3N9MDsFYFv6rZwcx5CeID3MTo0bwU4oPYF2/fuZ4zx+qkQw7sUppX
69J43fDiBPdqHQqvtIqcscbiO/5UU7VaEWb8UFpHVDN5ZGzT5VbskQtp4PNsExL7
fpyQseq9A54HABqGyDQb/+CjbX2b7hfjCWBN6cPU2JErAA72eGCKr/aTgTrutjYe
edSQVuRu2wrZesh0GqcdM06s3ZULn8f/QH+sjum+JLKyv66In8KSpc3+vpGWflYe
U+iF7p3JjIFaTYEqgog8pqdxRmP1Eav1t1itXxjhnHXcATTBJ4KQMetmf+T4AGe4
skRAPulRLPO3bEE06/pVy2RauiSAWcYmrWGQ0osP+YnQrcWnip2v4yw189QMSzkb
zhhyaODc+7X7/kD/bKPvcpebPQxfGDFykVVPKfYVe2qZ6IyVYyDS66LW7iSYY+NL
UBR1WT1VsnXbGs5OOzZ3f7f6kkxU7N6cZhij1+slrCuKvWHBP/uRaDzoF0yaTg30
GwegpGYwRdlkRXR/1BgzLhkoV/Ld1nuWouz937RIrLpa5yfPbVa47C/8gf7F2h6J
KyjnYxw7WXHVXW5aNnpV4Rb6UAKk0ppp7FNyB+ZEUacEuiJQqH0hRzQWgZWiNC9e
aY1iGhz0OrmnMdp/N2gqfHrzNrFW5N9WCeIzYa78tylO914snJeadFiuVZpeZQ5T
8dNEEIuHea2EAmuaStFtPEJiS/QiMBxDKenoDjlcpU5ftUpwygGNqFeBAu+qFUY5
n25D51He2yiKWJP2SUVAngq//k91V8XiGD0+H5DSjr6gllLnNuq6AX3uLM6c1gB2
lzClgSHAJCjd4QKMgGvCPwQaB+TolJeJirCdi5t02T1fY8djm/ZXKg3a+UO5Eqiu
I8eh/MTdgJQIo8SKSwYQBInMdrQgTYW8AkuJrESgqnUJ2jZURUFgIsBLaw4RuCBM
nTxBDY9BCmvlO8qypAK/wTscnvrTSWGlk5IO3jigdOmSw3KEvMuHYONpDoMKda/r
wuoFwmO+1Cnvh5EmacVQ23IKPrEy75/R/6zaFMDzWAkm5X958d7g2bvOTUdNqa/h
DmwigrpTuON3pfjCsq77egfXQ8cMaXJa4ShUzubgPV/qw3vn1RhV67ZsxfRr5g1/
J5UaNjWM+kgU/mr6BWzYgc/D6h9w5CDmYaSV+JAkfjkN1f9afwho7hI3c1Gix6z9
FTdG/wtVgfhm/9eyFIt1iCNeKUFa1zO8wDAnsPgkTL5T3/i0NKN/UB19ggrftgz8
I0vPwxiOSviV23xraNCPeCT29JOXNmemz6xnzY/0JCagPgsI/SW0g9XEXokc+iA9
woicKUMGNgGgINC5D0mZlpN1GQfTv6d5vz1KCQsnkX2b9vo8noJ/oCqfJub3mc8i
7Azy6CxxWoXQbuqQP+ZAWMwqML61Icouvqhi/4py/9W1wtBCZQtgdXF1APM1h7YT
ibgWQdLF3Kr+ELkSx9iqYY9nBkPhXwQCTnm5lm947eYXXRjAf2lA+LvcSxvHp43U
S8DRuQFfUIMaZYnqNRA/h3Z7KSpCh3vzqjkW18bz45cimj0PXykLRlA0Nnc7jvD1
ZUgiAGtuUmxx4N0MEIHzJ6gL6LPRQfz3TizDvdd6RrGLP+iyo9crssIuOzn0+otB
xRoSTa2vhhBSIU8yR0gSXJ4C47Azp529Md3QNDiNUkXWH03oXplkSQeAmhCf3fYX
gsim2TLc4NNnrivNWHWFfivnmYB6VENEHxRma0C4ZtZcfJvV7Adgjpqlobka+LDg
R2crdqoZcMdDqfsntVBT9K1WXqxecn0NRvYEW8TeRSOnZc8PBn552qDVM6E3BwQL
HoAsg90lozN8MmocB+/6IrU11FaR4l4SRDv0b+w0h8ZIBvcCJ3njS7OPbmFhxtba
KPX3SqhQw05SK99Wtqr7QrB163c2mGcQX8CvchhWmAoPT9UKacod/UpzVi6EgpQ6
re5jyN1XoMg8JKC6VCC9YhpFwczv7DBcF0A4Sb8/Oltham9E9Kcv4gk3KGdoo025
wCPnd8J014D36pgZRUmDgmdDlRqpgOn29dc4DDHm4k+JsmE0lCziO2av5U+hPh65
8lSAJaJEC3pzO3ugSU/Lix6V1Po/jn9cAdAb8+/WQwY6ifRzt1wN3KOkkJww0UE4
OhOxvf4CQ6zpPvc9ejaCsM4eNfiJL3rQKK2f1xdb3mYFkLqK27RnYHyNtOJ6GTNT
IshoUN7pXFz2IG8p/mhCJcNAOCeYPfLHtrVccD6o50y1z8RgtAv9DBIsl6u0vYqJ
xjiDZUWGg82tUBCBVvI4VnQnivqAiQg5aB0PD2VN2Gp8Cqtb2R582kiI8R9khur3
vT1s1v5ap+1rdCGRrHHePNV5KVhuxcNQTnBgWmfaKGW9w+Es1PKKDdzQsW9S6b4M
yetAcKI+iQLsoS7UIIZA/o8klFcFZ8gHFUDiETeCuTNotigijwWmD/JdBExAcyjM
tQIYfqrerGqH798gKlQ/iuqmTRhU1Qt9RoaWSR840nVWqYvDGNE4k9dQAK0MDWTR
Ac2ydLKpMr0KT47QrHSbvf6Es/cUBVuZnb7Tm1PWO3qwuPTBYD3ej5uh64ZhgsGB
9XImo2tVlCFGFXJNV/RWj9k9ODWWyPshxGBDmlR4QpNKYm41CJLDXQZuQ4XNGtGc
CHJkcuPsmYeopRbMluFQE+Ld9g3shEzcedGFJ4dEpThxipjm5HNbRi/q6Gw51p5G
zOP7QOklUn+R2T/muErlIbET0jF2HDVHnm9j3TEG3zHsbRhkvSIH2z1ROUX2Cw8q
8eXtLmB6G5d6bA1fMZRfGQOk2SVQIC9tndvakI15VKJYLDSKOJfv+r5h9LyZFzPv
DgyZlWHoDVK8HKJbV00qafz8jQlGAMOuwm4zIqEi3rWYjKI4MDfDKp/Uy1A1bUvW
48o+LzjPsj4KRX2meYKPHpr2E22PrYpqMU7d+cu3eL3TaG1SW+8SH6Ocix+AbKuZ
pW0p4llzfNRl92emv4unkmZZ8fwbX0e0T4I2TDuhyuRhDTVNKQKqAncAREThybi5
aAZGOOUXNbQZVwvCEdM3fjtXUQwFoHKBYZVMnzL6X8ZXyZyWuLRAqQ+QqtF1+cvE
C1L60wtpZDajOtwA/3XDpLkSBdB6rQU79rjx5xnIoPLQABae8TtK8c4SPln80Qqh
4wYZ2qEhf+bVrR6CWDypa1SDlMSMciF52Ifnf+6tuZY/cg3xM0UubBEdCxbAi/gl
AHi/0rUM+FQSRs1JMjh8LhHwY9Yj+QYBVf42CQ3IBB/eOXQ0qWXGaxVnt9/IQ2Nr
nWKf9WVE5WwTT4Bdtg4RdzlpuAhSRmifWWalX+CTtMGVSYJqKhEXWrQr54OxHN3t
MM5FhLE9JP88f+Nds6P6XUgcuPYfgOKAL0g4VPvvwxPDvAqyPJ0ntpJqJYbCvbNh
iTXLAIKaLqp+aKC6kRHHLD9tQ5Tp8cT1JQkSch72IvxVv+PbYCa6HbhISQwGgCd0
9kkte2z6bD2cSZezDdkLc6lVHo8dHUaZ/KRehZmqblRWkisj1e1l3o258FZd2LR4
A/XF9xgJDFnt/sbgoipLTLh9n7j+RW17lR1nVBoop7NVMXJHq3jn789PAfRT0q3N
B9p8XJTT8Ty7rCVHk1B3KYkeVbgb3qTqj2uyZ7iT578NzIq3ELx5wYEhFcdiZNHN
8rPlxcTucPlsHaQ10vhC60zEMWLXYkUxuOj/RZDJxMBLuKyN9lGfhcFOUq1Y4G6z
AWoQHZiSyrO9r1PBRMWAb0N6Otmhb2IMvMNe4alWklw8f/sgwJx+I+hExCzoUPJ3
M9VILX93sFf2kkVqP7T/Moh2CBk9Xn9anKPrZp+ZX/4u2EnhdJKsWmDSu8hxPtRQ
GiIjTpKKy2mVZjoLkXKMyULBJqcVPI/Lg/LBAbGh6HryVc3befO9Ytu8/A/ZjXDX
YJmOqA2qZRME1J1jHIqomXBTF5v63WDTlXYJNNhpz8CWNqaz/tP+PHk0+OdttGGp
IH5Ru+ntr6X6TwHBXPwcy2+mX34sC9lKow+9rWFUXnFELsJIOPKqG0nstZpuvfjO
eUnZBirW5VyVThYcc/9Bggc25BC/i5qHTDifsKcuO9vE6OkX6ZL3lRke+4+Vqz4Y
IoTAqlu/yQGRFuFYHxo7tYhsJfkXmuK14Px8aMqjv0SyA5ya3enuSL4tMWboTJJf
NTP3UY2HUziENJ1CUnwr7Ukqln08NlyW/CwiwmxUtAbCFeuh7KUgWqunfdi3ReBF
5BCg6HEzXNkmT95IAgPMFAWug8zr9LfSZLUTaQi/HrlchFEVmWGU1BpPj93TKnes
15CIUCs7Z5KZZVBb5+Dz8O2WF7QwZkYgTJzFIjr3AjTtZqzrzseWM6+rvOq2jn2t
0MV6pOuVYNJ2w4vdHTCyDe47Q92euqVsESy4JLUg9qydxfeE+ED66e72cYZ5I8gq
WHh8EEfb1Jx6tycnsEkcgbFoKTLc8rH0dV5oV414ZszDQgRwZc0ThKJmjTpATVDz
1I2uThyzV5TaFamzw3ZUwJKXlPY+smQJzHnf52cGoX4P49CId7c+qbnM0ce6zdIX
ElkpzM0T9WFg7xMHpFcciqL/81Pzj1RDuaJI0CQYnV1/k6A0dFSimJ4tDiUdhZgD
oBmJHmcPELxpHz0ClNxcSnIRLOECquyMt299CJJUAUPFSB8v3TJE6TqlZO8KTgt3
D+zfvv4SQ8HKuGOXDYriEZ4Uiu6NJ6ZBQerc+FUK2hTde4ja+gPUq+U+/DLJGY1M
Sta3Z9C5OjTw6KGLnfXafY6Ud/6zt8yuyAkC69ckDxyO9tlyDj2RFNwczaQOiwv7
703Sati0JMfeemDpP34lg/CE/9Zo/bCedmhJ/eiXqKeTQTTE/tBwK3RbOXMLJChf
3Jo8sDIyjeREMQnCsfE+RrIJnknfrWCMJqTFmVCjKyUn61QOvxexBV5h3VqalZpi
M60jALT3VuYOTS6ZXBZzlIrGETJRS0DoEFzqZMUu+y38dGzHEKY55HWbzUfqDMbz
vzqzLwry/NQTITYmUspC9qMuchWrvMwIDcwHB4Z+sd0pQeTiak1v5fxlYQy3Ab3i
ugHLdIQhMhk6E5C9dNdDfLU6hjqDRzP5sX34fOT8Dsi9ZxIitZUL4MqyPzcgUyMv
4j1ABppewM8cHBof9ShBCNQYEBRdcOcGlUxDqKn8LKK3wWmHzB10RDZrfftwFvVx
OAYQpQ0cU/PLesB2faNRk9zrtVQ/0gAw0Q/DRA9K9+xg2npkl5GojCo/Pa9nHtgb
Z5nQkG4zh/xNC+CBUeaA9oWjOe521KsMD7ebQN8Xg8/x+ESHo/rgt+Ju0leNluQQ
hjBw9p66pA0JwRWLeGekeYkjWoF8A8n4ZLjVLshmh+H35s5jVg9/Lj/ZfSfcz18k
VSBqwAypFFV82nvqM5SgV8B55IOCRGYXijQ8bAbK2iKuEY00xOP/Ie98ukqN3cEY
K9LYNOZziLhSX7tOQJCMOGxXMbG0MQiB3vEpp8no0S+fzE792Q56Lsedg2gTWJbW
0VlHOpUSGPtM2MguEIBxYPX04O3dmJOJNatJQbL3Vj/6xstSmoTKD40LHwCpjRKG
7pL6IR7YMROzHqO4vDtfROdh8r1UpqplpdHE6sCgNuh1mudkN5VOndgLrsnlu/IH
pqd3XzSqa/CNLHUwO83Gl7KVaihHSGh/DMmfD/5Yjgoh+Jq5ykN9z+G7IIiw5gt3
jIogEzqhfzJ/ImvVmIiC2a9dV4B9zGvtS4aheGhEKf3d4cRzLfPp+qZHWka4FwMR
QuxGE36oBnPFM/DLLa8+37C4ic9cCD62xSKhNRLEvUuN9mlM6sxZLYgVq90f/mFy
fMO0NoBBv41lFNzV7AjmPm0tVPDhOkI+HmrhynhZ/BSbem2RnA2eq/AYB9jz+PkU
IUSf9GhikUZABMK7KnGItr6npaQJyKrodgVq55S3Ct0Ar1fDdJ2KsBxBDwZNdeKT
NRQoijJbsqNXw4hNaA53CO2gG69MkRlZGMiygM18DsTfEouaGuwdfP9+ugqmtFCq
wPhG0plg6aQUQtTyZBr1zeDnfd8dyo8g3nvrrI5AVephLpWLAnz72Sxfj8PGomrQ
VPscYTKTevxxzgrloCtTpdDtvUE85Z0XJWv8kakf7rvFirbKXOXY4bHkaXrXh5U9
FGiRTCTBYWVMFnWCegt0+sCA6zRXenMI6g0UTZTTVaUjIiU909+foxgowZcQB1lg
EXyWJ75pukFdRtki7QsN54IX4IbVz1xcqFb/VrxBjzxoLyI6ReKdvr0TfOJAHvjd
IZwUOKe+debbQnDEKFTgYcZUqYaDfJm7yusUUifmZb9G6uRQiqZ95gLDK0RSO344
DajtfhIGJa0I7j9uWk1jSB3oawuHype+TQH9ThXfi77gKf6t22EPC531kZFGWCGN
hhmZLfOa+jQGG/s/tj5mlK780xLfrTHfBTA/eo94W4Q2Jl53zw34A6KrGI/vwDoJ
i95Q5y5C6H51mhGnLDJgBtlRNZ8pITIQx6ca6oKn8jNsOfic8T2DfdxOs6ymiGoW
J/A9hQdHsUmT1kHk9SaKNEizpCH0NjTvMIsIQK1d4D1xblygZmqs8sesEiEquyep
TWGnmjm1WbJuVKF3ExNuWW4qDPBHqVLfMIUbvryme1ihPP/UcjuYjUC8djzTWTDC
Bh4aCp4jCCa9M9Shvl//Qs+h/Nv956M4y2IWL0YRQF6KSIhchmqhEAzGQR+fvaSH
JCJX2SjkWmNE8YzARUbZGSTbAMOVBGxnRaPzFo6CA3NAZKpzL66/SI1GrRcRYhSC
TieBoVN6poPWTrHy9Pcs6P4oHR9awKaWHXbml6CQxTzONsW8Yhx8RyFewYvq15cf
Wos6FJEwR+N09ZLfNWnzCodWFRwK90ATlhY5T7sgkYnvYAdC3qxgLkpmB+m3c5BI
oRY7wY8RG+abx2ySL2lHSaN7/yxRNjXUg7kRD9A6bte+rV/8yXNo7F3UMoStYztR
ZQE496QyAd69ZLGMQ30SE2ik4VKENulpwfg7B7w2/xdN2u5agCUQMTbNOcNNGHe2
T5VNoX3z2fPAEMgpiLjQ6VGCW/qO+9dkZ0Tof6AyuI90pmopi3JIj/K/YXzbjma2
oyBj/M026z4kdM3dZlzmLsO3W2uxHTMQ7UZyIc/k4dtvR/LAO8OdwkQQswDnaKTo
1pS4YbnJfDkxSzihLE59lrIhmhk3fq0DfFXzOaaVT8tTaLNr8QERdG1ErUqPwaba
7y6DDuc4SJatGwgzs561Li4Vp8ktFypUB5AvsDY5eTzcHazgGadnRIE9GM9KNSN2
oCNHnycsC5XHWsUcaNAflfeliP5J3t9f9+WtZUek4UEPJ/ODGvF6T+nWpPgsmK6t
F9g4ENZnllNdpbYycIB0piweBUQdXNNs1NHpBtUERjqCWiVIDzoYIu/V/RpbrDCf
XS/55tzXaiV+tictFCGbosb+EaWKCvNruRwW8F30AmOU8emmbS6g4vc0RlCkIIBA
NepRM2b+M6Bd0rmmNcESpcSgsH/guxcBPykksTYpeLSxhNZMkDhKTiZBHmOO/I3T
Iw6h6C8PpABOv4B1G/6sxSdl2byn08sd3YNyxD2RYptx3KQxpLWgZ/JU+rXHUBup
uknI/A3AaAvWw2jlsKt2dYnQjflENe5L1pjRRhzUL5ASLv2X4meBQb7xydaz6mvx
A4Ugq1IqZMXI98/g8vzrQqZ5py2oHMvqQMXA5f1qtDlpMg8uN0o+7yDyo/qkKEDp
EgyIKyPDKmNu6Fpcg+s4vLVNiAIIMnuIDKBNjiMC1a8jsfPUFa1ByUTxD+Y/NSJV
hoauMe+Nwwb094XFkPvDLj+oq5nZW3ZjBC9lD4iRmsA65CnjJhZR6imb3RiAU5pN
gKYYAs5BWSnk5OvgXXIOuReAG9qXOXY5QvmM8ggYAKB7SVc6e6g9NrVrWnJjHEem
vjrZLcZDX2dKridGgzue/75Of2B5hAVHUVeZRT1EFvEbNc5k2KaPaArato1yvmsY
Fx2UjrBFP+q/9bzzZ0ddp/3+FDw+Ubg/xhhH/tT8VhVBDk+zG0awx3SAQ1qv8NHs
mcrPc85mqvWNjZf1Vp7gnH90JMsxUNGZrbOf/5kG5dWEjsVz/hJWPJ+IaH4VyQgf
9KQYgNN2Fl0oedhJRAjWY0YG1aIFNliT4aODxa4DrX3iZw8dNvICRF5zEtude7r0
7lxR0Eb1bjrOV+bc9rJ1CIQNg94+ehI/H582x81VEHyAfP7oGE1odBXUOJ+/Nhng
FRuh97EYa66up16pvRpwrFy6hz0pIVz17Dx/dJFglSYkg0xrQyi1T6OZM5QesmoL
soO7Pl5+ulpllQ2zXXO/Y/x4j+sqGvWCMjdbyXZJdHeWf9CEEjP+GiLLPKybJxLP
h2HZEdaM6vxn32Ftu1LInTZXNIZNQRcc+AqbMrrYqAfhyCmxP/83jgSBY8P539wz
LDi/5lHivmTX2NfeXLaabRJZrbVEhPSE66lF3qiJvAj5Te153xO3Fbk8dcffnHhy
JKMDr55UOrkN29pR4nnwjf/rwpGsJvf9mL5/g6cSVZxLSdB2lpm3XEKaZNoRVwyo
hF7rQK5smBgPh38Npl5/fFKqqMdsusQ05Oi7NBlgD2tULONIWoVOJgELIS/z8hl4
q3F/juqkaiHWICAPv/VMsq8k63RD9sm1KOuiMoxWJ2idSSdldt4kFGzcrXzzs+ST
PiLAn2qB6TCVxx2ww/bBFd2COtCC4tMVkZmxF8khh1oplTpluZ3tgQ3zdthx2rNm
dFyWQa594x8r12euLQxcWC6ICNQbCgMh5blLy/rnUVHQgWoxbpWoeS4qT7+SqoiI
QWTHUueLb/2a2V4Pjl05kK9SG9Cy26rj8NdLYmle0gnAT120y2yL1kJXTgiEr89F
T2nKsqHtQJE9VJKZEutyplKcs42UUeYAJuitiVVD3XkeX+IWSJQHhP8wnHS6IAcW
/Uy02wXc2alD+drQVcUJqCHQ1bhTRa4Jiz9c93nLxC2FsXMR56Jgf/3+grnWuZWm
ise688nxKl0ntR6tCxbjNSVA251RRMN2QGiRqww3f7E9FIaUifgfiGBQS5gPAtDH
fgMoaEs88F0U20I4UQWKvZE9GQGg/9m08HuzfPFGYqXWcdwahzEBEgZaxdJOesM7
NMd7qxj/KJEbGAQt5Ok8X0tbBuo2To+T+fj0f0Hxn2S5zaZbh4I6h6k7uyjxnoK8
YN8G8d6dEjGvhyv1lkgoHNJd1WKAQ8tMnJuAjEQjS1YNly9k/fW4wNmchpqYQCXy
WPIA43f0XoEsg/prmkFQM9Ms929IceCe/dqzE9jJotrjuOjuyGM4WvMWme+M8lAW
ZtzaIg1OqiZVKBZbu8hEo/mWoG4ZPPI7RIWjZZ3jtfNHtPRHA29RLR9YsNkmM62f
dOGvsechQyNwXGTUddKRHTPqPvkNmJyQEedTMhC2xl5jTKEvYa9CAMWOYLLZRB8K
/JU4f51UGmloLuRHhKwrYxnL5/+ItZ1z6dpOMObQkUhq8ty1Stgk584qGeZlxXEb
IplKiaCMPbcl+NnaSRwi5FwSujjsuH2uw8969Aaj1W9lPkAp7iXUSmc9vrOKImA0
nUHafHCvJhEu9Ddb79cOOIL+rnka0Tu/Zh3HHExZb9/XPBTlB6eTRfPkVP4nTddu
5wnSsPM4N9aet26/VYbY+ak0F8fSAUmuuUBNjGOn0ggfnkhbshq4yAnSMfDPJ3pg
7eyU9PASNTQBVOVumCcirNP3gLge1Kix3mbpPsorugYqzNCFeVwHpMRjdo/5FYjC
nv8DvcT2xJI58TPcGDvsXkHyNDIsIT5AfimlLiElUDVRXpvXL/juRmvyXh7W5SjY
QYbpIg+GyJZFr+69UaQLb7RP+bSu6WPrZRhtKrJ4r3IGhcZ0iz0hAzMO/BoTRQsj
hbvFZXY3yxf9HSp00w/Z0lw+aMJ0+uzaA+/JSOt8WJ0m4de4xriu6CFsMLSdu7BH
BuumM97wORpyTgojCb/5YKC5izOxLYKb3dhyRxe2Xg55fhkAfn88M1NEsDHnDwOi
mOlDaUOUhubQlRyd5elC2GfFO65t4hLhNQOvEHGVWwowJV4+LY9vVk7pTYULBBeo
+ZeoFr1TbGbQg0whh1s7Veg/U7ai/W8XdC6UEten6VS71iHss7DnDz3jD5CXlM+N
R+/ZSAUmrglhfhzOCChFrUm5wyIATUJpC9ONcue24lcr8ZV8Q9OZP9U7x5rOtZwB
kiA60H6aO+0239zF2aqa/+XKjNxmzQtlLOQoqVbQzvLXuEV3Tu9ZDRECEbFvAPpu
9lXAB+Z+3cGiIakarAzEl5E8oTgrgrzyUJfqGZkyCJGvnDROe8X7qiV4OxeH1wyT
9xunENkw9umRHdFbq47eYjn9K+31f6Px7zE3JyPhiUvTRxwL/nqGRkkejD6wuv+p
gzD5mhGZieOknXkReDFF4cm7aPp8rHgF2LjBdDvgaNwmJM91qUvXbRuO193ptKup
OlM/MGtyboYQPv7POvhRzTuZeDNOoc/fErw37/KMFfPe4uI3HDgQgjoELXVbzMCI
JJtqVhEEdt//B3qbM7i3IsfMpTsiUCsRfW6yIBvY4xK0GzbmFgwg1bFJXATGOPG/
mdp2RJgITWhLMjtNuvu6Y/xODfvsXNsaKbZbLsUMcFI2ZogxvotUVPDxp3Ho4kya
ezmzZfaMewUNwVNcaZs3uapitbP7SyXOl2mjIbPrRmWrsI95E+UIsYPvlJO3tG9Z
hhRy0VjV+1dn3W7IUXXHj8/P6yt8hNV3Fcs0tZt/UXTcNlhSiw5tBJFjXRLOUhsy
z8cLRYpS1OVpQy6i2BTWwfGJbwkhb1L8Q4AzyiaEJ5HdvcALd6m1ADVxm7MfUd//
RoJOJypQjKfWT1BekAURqCZo6Hq26KaPOeBGvn5i0DG29nVAMw35MSDMmlvCOLOq
aKiphZm+wPinrS+m5TuF4wCnkmcws1WoP+s9bZiXPrx3ylSMbPfEBuhSnBluKUPm
mhbDTDy8IB0HWdU/XnCgeLvY+YTa1Ue1cISvjpMIe9ZuH7FTypyC2kKXP+UK6ImW
/585kqTbjkg1Wxr9/dmxccqSSULmNs0aOP4L8QESNAKJH6G6It1EEM1hT0/rmxsI
LqKY/4tmYMA6gTuvksc315nKOgKQysKIT+UiswmzoMV3W9xTcIOjWz3tq3hfMaBW
7sb33ZvJLI9FyhOGiszs6r6zcO/tajAwwmMHhFUOCdbErEMoUm0IzV98xXUmwkmi
bYaDO2Rt4nhtf28PtjpCzHyZjMb+UAafQo43ItKv26rqHhprB+RpyGObQ8LkxAv0
J3fIYxF1e37NNGInb4NCOQGA21bQZcNiIkW3lSQ4VGcvLIBybtWQNj1R5WqCb0YH
aN7Ts/EVMs0Uo5h6ynaEuVWdQsnq46rlcr1S63OyQ1FvXME+cIapWDU1dG19EN9y
xU987eTLWwrdMQXE1ugbZY6PpCkP41P+yxZx8eT5MIFGf28majwjE3TszE6m5Jol
Iur+SPAWjuDlGdaGcBFycsmq6SFWrx330rwYKYohXGpPDRaaCsoQBq9aybMg5wxf
l5s426MvyfOIGgHh55uvhXdMPeRwz+IcTtu8MRSCK1kjOy18t+8sM2gLqqgJg4KP
6XOqdWw+xuIVA65MSYXzDv/Mqj7K0G/dUoqRNT0j0U6PkCDgfklDygbRu3B6iEfB
DP1hlJ/vRdjxd5uOmE5tVOPeQl6bQ6yhmvR8jofatJoVWMmgP/WBYuq67Qhguri8
TuW5WZBQxHqcANu00u+R5y/xlIOWl5dFryS/kPmt/t5EXcJW98tcDp8HeWn8d2ug
ZqK4d5fCTL0T2ZPYaHO+b9TV2BfOfmV37eNoO0+pllkEZgIm+9okIfK6a7INtG6s
4tFnR5SWgl0e6gbY+Y64lP5Ut8SgzTV8/R1hEjjsIVGEx9d937YrMrLD6AOnylge
vCR4xQBKTpviRKid8jCAPr/+Jh+7EHo7JZ6Ya95E5Hf+B5YEfKiIwcyZxq3pXYiy
MwUVDmBdXO6o9X3ezJfdidFtjIqowOfgHZQOF6LHHxftRpBh7dulgjlcmO1m96Ob
6aG7vYYQ4dYASs3N9jSGf8k8byeTyY6FYdDd5awzJCgPUoSuJ3Rh0Y5OIlhhXLGX
uoZ9f9WxplsoNLUvzs0/gZzJugH988/MEbTDqDWNizSCauarSl5txJ4mquuPacaP
kaea3FcgPjSrgThyC2Vej7jkVeduLsl6wWtrca3h/Iwl2W/lYFsek9aK6uiXZvwi
72+dwyNs14OlyG+t9YWr0bAU6uylOVOPTvwvkQNH42WbelrfcsSFcXRgVe2k8yt7
fJe3kd+I3G2V1sxNw4w7GSJJEh7Y0hSC5kh5wOvXTXD7ob9Oe1SllmGAy1XytKNe
WI6xQqtaMguzE9P0S+k9E5QJUDK2QVAEWLN7C4Pv0za2lr+BkLsmpXWVGiHHdvy6
OLRl8LRJ48n9u+4yNn6J+8iJw0Jf7UgTPRIF10HWXjYwHJghtpRu3rRO6jEiV5K8
XQ2iueq+ZXeA/A4bRiJmSP2tDXWNLpzrpVkxTociGMcrUOee+acf4YWZis1y9fnW
Nvkl//kadB+UdRPH5THQwSpDWx3dwkER5okWkkYgIVhl0c5tkaNlTm71SuQXdHkG
ITpJ0sQLjpp+ju04f3LiIcdoWsk7I1l/ohJEhhhevFMO8s58ZL+DG5LITipOXh0z
MVJkX/BwuGTqS7BkRqX0IYvPUlG0eELD88x6f8Yt651pD+UITr+hs8NCHDBCsgpw
3CJXfWmgzagJWyU2yLyry/WVP0cpjxdF1Yki/iy15DOZU/kPGnpN7djaHemf0o/i
06wNLkb6jmQyOXv8k7CPIOJ1Aw4mhMPCOTtAXzVODWHFOkH76CSbN5V8dfLJtJWM
uk05qXyA+s67mtt8oRolu4Ful9v2Y0grycy+2dgfgroQrt2P8dWUHtJUpIvseTg4
Zd0w5Atx9X2IZEgZGp7qNNZ8ollFHaBws3zNAbTZypoZhnkpB9UFBQLm7r9OdIQm
0q/rX/oEtFxFvBRboMpUwK8QESU2f2Dy8/Tt0SVL8zF7CgwkWMm6/gJBWKq7mJZJ
YYGVigS8XmipwCYuaKcgEHGqdoldiBlUkvNh51XuEpPLsCdXIBjgcul8TEDhTLIl
/sO0SrT7NaBkv8lPXolf7X/FrNTcksLcDwzxBEQfJCp449GWtTpMqyfJzq1w5AGK
a1eXsJb6pol9dcUCsTVyRo+FCX0zGjnyQ1UQF7kWACECZCfM41+x9dEeIcBK5gVh
/CqO47oX+yhrjsknZUzSEZWB/RnhleO8xDuvurRu5Wv7waAxC/mvudQsyHOaNY9s
Ng36iv165l+TwvJXpDmF9MCLISKBzgWSUbXvAVpCHpntoAGTI+RtD5QdTc5sXLZG
NadNBzJqQ+s8gebmGBgSIio35JFBNQdJd7Qqpn2LTTeGsHIFJZ728sWffWzNqs75
QmNL3dPyGYWTkej3AnfHRbEowF4PKQYu1peQQddvWk8BVy9seFpLIg8g62cgSOqj
5J6NnWcAYgAQC9L9UPQkN8nJl6xJVGV3mRncaKnbrIJrqT1G1GKXmxfXhq6UoRHW
IE/1XgA89aa6LjOMR7Q99XjkHWIek+cTSUAgRR6jceA8lak28kGq6w0wukAwKJYP
q0FxrGBJ5Nf1Ucb2V3QvnkpRTWZyfHPwgwTdE3vlZJrgkuM2xJ3NpkLFqnl/kNPq
AQy+ifhOJTckLPIPfCgwiF17SIWqOtMc0i1+vM93MQBIe+kGjboeB2i0V6180I9+
CjMWC6LxEQ7BH3/CkyaD8cf03ihvjnjW7+Wn5m92kgnriT7Eszdk+TicSgr+aRfp
mC6zZk/gOrcphlDyakgn8uZ0AFS8qGwqYXKpmrDpUs2JnS/tQR71jc/lOPvF7X0r
xUOfRC1mhJcLHII57nsKmXNIt+EV6AdnsVLkqAN9pTdIgkGH8l7BFYyRPRQn7REg
XbFXTh/8xItU/zYl68iy1jpQbXc7eBK/V9KiyvdKpwBHRmC1DXAiFMCoKQrqHDCD
ypBcqAJnGtcmzq31rWk2KiDAw6UHNcSO5KCmp1/UAvXFp7nEW4h4d5XctQ2mRx0J
MwYbMw2flEPPFkcyXqqfleB+vwulMYzzZxXW+zyaVsQZSsrB8WeTKR3NhDPZMHpi
5ZO0bcMlv0goKOu9h0ueFAoNUngxR05/VlGEhsXUQzh6fLPD4WpquJ5WOhHkDTsT
TM62SCQp46v5vaRNX1MXxsfsbPYqS/DqFujs7IDbiE6iKAT+2EO9xdjNpNrRPfGy
6Gu21xjBk3hdE8F9c+JgyHum9Zeic6POuB902MPbdTaWbjOnZGqgJXIFDHM8Vh9T
d8nexS1hHwPWYA2kYSQEufnGesDS3g1LWYCtcVNe4Xf3A/37qwKHo6XF/8fbcYcL
yfKxBLO8l4E+B1KVit7i97vR3YuzUYWtTIIajV288j/TGs+ucMYWgeRbgzRVs8GE
xVb+Ivqs0p6bE4XydKOWuIPK9QdujyR0/6PcAjmyfQuF7UpeSSqJNAhNtGMrg33N
tcwuM0Ng2DcnqugzizZXd87NAF0PLTVt4lPU1COqTETCHv7FLKZL7YHX+o7FwmBj
b70Lhoxs0Es7u2z0/nwKrVsy9M8bHAVIlmqsGvJfZ3KyvjbpvBIDFIs5MqtMge9l
cLMlozulfQLzmQkkPC6fPeJmSm7pmzZ6s3s5nWhlU3cYnc2DGdcD5Uv2RMRbOJsC
uq29MyZsPaKSYFdqtQ5S2cqff2ZxKtQ/pwlnxig0Cb5W9S6C1lyiOJT5ijDK3tSt
/tadmmWPPD7I3R3RC7ESknBjDmZHTNFOgvQjvtYyivn5RxIzTlXSwP+ebVm28c43
79pwaaoicuBjgi6T3ZhhZrl5Rqe/24+L9/oOrIaY9S5WGPiRbdBcsqNgk/0qy28S
m2EvIhbzIlZ9nGax1s9EJb9UEKfXk0WxbsnqG5dc/RlCAPlF9AXVXb4D8BKuwI51
7CMMvngLrTphCIPRd5z++YySHOpzpk/k/J6lT/mMgo66igZZ5ILiPHX1bjbS0RGP
PJuR2/ucA96jJbzFwSC/uFFNUpSqQtjP2xLaN1qqkA48NyOv5WefoMbTUL69hxPR
RYfLGzV4+SHlvJz+TfTiPct7EoP9IEywVw8ruWuGVFNfRMBuF8M5TiOZrVw8BmqD
nEMDe1BGMUgGcf6Q1uXMvCh178afcbjiOAZuoDpy1sY7tCeyGlSKlS7PiPgM4sEc
L5ApZqiESUdrGw5nrHdWdqbuJhaR9pCMVlTVhMpmgt2q1Z403XmQ+rAqbCYTQgOO
1/o5V65lqUcpxQ/Jg1OdoYoXFq8om3P25PxpJuO7ilCJwdVO/dCJraVn3qZBxdyF
Xz1BZkE7x6Z8qQjwu08aRdGcv60kzkZj3v20cWHCHx/rxtvNIGHvqEA3+zWiLBi6
23VddT5blTFuJHprD5UCgDWIsXuwGGW10iIKlrtVJVY9EjAXVk2hqhQ5sAzfDX5e
aIDAIJK5BPG8xl3qaUS4Cx9mAoeHpkH56nAXoqZY/X/9Pn+xdZmdMXEky+eyPeiB
XR4NlrIaTA1Dy9YdR7T+bE6dqbamEqAYx9LIHIUgssWiga7wK20KmjmBhF/Zn5cA
JcWKXbOhxVbfKh5qpQlSTV/IOwv85pyw0LF2afZHTM6Rtjax3BszbRC8i00Be6jC
PYxHqS8n6svJCYBy2nthLVkbSPLoFf6fgJwUm5aaDQaHHMnSxB7GaZXQDm2CRyMd
rw9OqhIa/HWfNz/D/pmUjlWRH/CjYqrf85If6+WN0Weo21OfPi/TH8CuvcUzMJxn
3RGy7GA3BTUuakRCRyIHesAAi6idbIOgsBImQnJvUa2VVcNH8gtwZ6x5WuADy+6x
EXkGCnt4gRGzBwROBbNVjn2dIlbQoJ5O2mLdT7v/x7Biog8smtWFEeX1dUZtsZmb
ycb5JvwaEU//jIbvf8FAk4gXUKffyd/RkFzmI8k6kLWWR00mEPwvXAM6ja1Fn6Lj
3ZVvz5ACcgnWWfadLWx7gd2N4IXTgNcMsotyPewXbVUGoBLBpoTrOe36ELJBAJSc
qfwyLwhPXNG3m68veCi13/i3Ujd3pVGc5LA9ONfEZKaiV9lDnKBM9tBtziTB3Ahg
7KyD8GYv+wgmkUUPxjS42ASz/UIxUmgdVevUSjotM9COVB88lQOQkT3lPpsXAbi5
3nxUu38N3g8calOF/2o4bXlx8/H7fAzJTlGjEWS6oyGYgrFRcDZcRwYD1JKVpoMn
xV72B77lDQ+/XqLktb+5Hp+asufIwJhu5Cr92LOKQeCStLxbHUeNVjGkxdJPO2zH
zdxb5p8y9XQYwmYf/2kl2unHi4ULz0wwXP7PeRUJAFxqj72g0riz9IKaYbtyC8Ut
EIXTpP87Iow8XolOa5F+JbrwwK/g9YKQSoduWAfrrNEEsH2P72WqPBoh8W9D6J5t
BX9FeC7IpV0I9qTWjS2NNqaHC/92jX3d4VlZIQeIyglbg0C0EAue+HJpOvLyYBiG
NUat28YiMw/yTWB/zUimIpHS6IZ63bFUm12pHA/DC/ml4NKOa9pop8VEIq+qOtf1
Ivo8RCLUrVhZbsrxw0XIxmn4DzKjGiI+Sg6mKx4tdUBbBTNM36dQk7OCOoDizxbB
+oCvKYs6Uwy5RqXhYjbpNCUk3n949GAY/Pq6DXEZqP1JDzgg3yQxsKffRdwlztB5
IPMM3ab8EXsaXZXFqhwOGOS8WHM7ReA25wbYyCQNoL4wKwU88dRyVReDgBRz4PcK
VhUVvqSrKIR2mVrRsrW3m+4QmGmkhXGM3A5YIoYwhIWiGo6eRZM5zh6mNcP/eF4E
tWVmt5WKY5B+5kit9375lLVeEjAa4G+TGVq2cMcfwAuTkhzD9HGdliGcXHI4xHZL
J+C3C9VN1tZeNDUufPqvKyReZYXdYOKI5Fmbs6mSq46cqMOyPdNdA09iA8ZuAQPh
3r2g2jaR/MhUBgu1ojSatOw2W6mS5qLFHcwe9gRIHyUL9GTDBoTo6hDe8J5BlCNk
uuWRbhqOx3UF5iapfuFVytbTyIbMDI0LmjFcDF7vRMYpMKYcf6D9fZk/nZxwmqWQ
2k8IQ/iBCPmuE88XVgDogeC8HIP6bFboGI4f/LExfS/D6CXvBHnOcGUrcH7m8eCf
M3Kyvbj/Kv7mMJxI/1weXNHcFudAFgnuvoZTE9+kR8eKLw2TIOikOf8fT/OeYXPu
MnMBi1BaMp3fhVQU0tiG0blcdTNqSms1mA/o0x17r8fMv6TywodzXBaG8Z+/iV78
NTi4pBPxZzaF19hmKaMGp0Vu/j7FKNCuN5hyfiNd0wMvINNKo25XgG+3ec7QmDSX
rhOWs8xj/zXqMWW6spkffE5VdrmjYuxaqT1hh4pOPEaPGuHJ8MYuaJgSgf0PEa5w
IONmV7hVhHhcD/4qskvxTIgj37LNbwuZqdrhVWAvL7VgmHil7tNBDmXl/+U3aPyY
Z9JKrBWCO3znbtDfY9FjJol5a2iUPgypr3Mh7CEH/4A+IjXcjeLjPmldUBVa2Stb
MWNCXq7Ss3ubAMZDmwEYOf0unYvFEGx+yd9SjS6Zl4hJvI+xC6GU5HnafVGTU3VM
hiEyyIX6HgUVSrBTN1o++VN1KUllCVs0Pdb7qZd5rgb4gZ8lqdnqpFZx7lwMalnS
2lB6hXVMwBuBbKF26ugdFEocSQTmGwyW+VKEv9oJvjDwrHdOEyfzKk+uszTOCeMK
225ZkOcsDvEaBVR0kOsb83BbSwm1MYOsBMY+SMDz2BcwpjOR6GhUhDjJdYg2vD9U
Jhf6VGDiwAyvIJybDbBOFj23UxZSuEu+z1lI1wuyjY37iT03F7j6ccZbIlHebm4T
/SFo2ARFUUYD8jiQcdugRQEOywQZ+3EeWN4SUHHalKqbHx4lZIXpr9UXYggxW1PB
0Hxqufg6W4FhIhB/KOVM4UJbvAt5QqNl2Bi6cktBx/+ldrly7QNHq9w4i3722F15
kuwGOgICx7NThksOlyLeazXruaWxamF2v3HQ5MtQuxTyufGq8xg8DmaFv/kJX3hR
4GUuUGmuDpayG1RisJbyS+o+aQ1PF2gEpWbwdj0wCGof8vSerFNkHafvLXI7RJ2u
AF46QyIaYXo7r3B6dxIgzv2wixrrSe3MASKlKAh6RZDsTrIgydCAKqvsN2FLdnaF
9Y1XLqePXsQblsxGjruMuX6WxHvIqtlA1z0PLAsRd8pFq8f2UdBnUvMTUtPEVFqP
+3x0WH0KafKKP8/Aji/ReXL8G1m/LLYRqcPZ68YXVVHsx73cMoVjVt8XVNnMRbVU
eWKhT0Cub18Ifvg71Htk/lRCSCp8r5H5I2YVoNBfcKr5a4vgSLYaNu/1r9G1KoYQ
w1PKv7a8xYn1b5coI6lGTo7OVxr2srn3H17Gwj4013Bz+iV4PaZ6fRJTUnBgr8Vh
`pragma protect end_protected
