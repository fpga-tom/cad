// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ow/lZ6QSsFFS7aVq5ELKsJLJtwlzajeounpdSmzQK3RHAD8p86STQf+okOrsMNgl
/scy6s4nLYaWW5xXIylU5gyuazxPUXc/zav3YWuyxK84s7FzX5Jc8UJmtIyvi3er
/uczXwSvbrVQOx00eiUyCinoO5FI5rh86xJeeFqSnqQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21920)
CRxAmZY4pGKjphrhlJiNVfOtAgNzNhuGiFFHHjVTgFt+17t9uRhzHiSIYjBMO3/t
kyOa3Mhr7ZTabdMRDHDBX81wqpDIYqADIwPle6XkcwksBe1gUEClFpRSH43izmuf
dMyENzmD85gZ+QoKqbTyuBsuBJcIu0L9TEhxMAb26VBqacJs00zrg7BSx9RlHjof
u0kWStGFT5USoI1/7xMn5QDWgHVJOVzbJD5jLchUFUbjYxwUpgbcqIUusZe3deBR
53sU/2asUJE04ftPg/5CGglVWnJIncNyb4X88F4GUMzAKV/OlwDPsoUCgJt3FNfm
MpzseDMEHKDvbvsu7Ia3pUTlpCF/W8d9IRrvZjtY86Wsj7PR6JZOR1WiJe+tHi7Z
ScDAvX7Jox5kRgqoR2PuBuMnl0Bl7L6rgzx4Wqx8XLu11irPf2Y1/ERxrcmPh/h+
wHY2JQQvhe12ixQvB/eU/eG9bOwVWNzFP+eqUM5z4Kj/AIkQ/etoSsGMYrDTM+lo
/H1+sWRRRhTIipzi+iJaCVXKEdIB3syf+MdVYWkxr0W0EyAfKVQFrLj6WYc/GT+Y
09lwobxbBNMURFqXNIwUzyXWsESARpS2ohPJAjkHUjHj8z667ABXnmiWVCFd3NHB
aHwvEm/4TZJ/TrOunWNAvR6tMcAeOyDP3z1N9Pm6b+qAT8Cpom0xT0BsZCQoz2Ei
jgeoXC/sOlmRFJn1eoVRZ8/exuxHnWqV74e9ium8B0LtBI3Gnz2Mlvhyd2IvIcDh
FttRotAYyvcPrSFTrjHL6T9JbUN7nd5S3sCIpXBKUGeHWeUEULCBH9zMvLIapgD4
fhnaiiQEzup4+38DrakWNQ5kiDQAK9d5H5hf99etH1sws+PR6ii4FcFngSxqX2xU
IDcnr5N8uJjYu/ALUESeAEg88PCg61jeTt4ZEF+Wi8jTq9Qy+mZj/e1cBzPjfVJf
s2cMPxHV9BAmcONtwuD536rCWXhP0OSF3tdcwEnYybriAqjzW1zf6DjMY315WU+9
LqNLSn54Ja7i/RNvEbqxgqinKfeDvRARIxGxqjZqGq6m3b4i5uKBMD+rll6jcEDW
D7wrTdPVbLaYEQ6pLvJEWBUy5EDJCEJDN8/V/z6ev1c6bK5Kn3QC0NB6eM3A2TOp
ffwkJdfudRuQyAZB30WxDlCxE7ZoVgecuzeUKCziLVgb3z50RbEOboQCFMHLGTYY
iuoltz/UZ0DLvwhxKOzhCul/0FgR+YD5k2Tw2O8hHffQSJfJkg/246uCV4Dh9kHR
u9WLj5a0oMH7UY2v6ByxuDeJdhByvG7UAmo9O/uTQyBG0Xaz3fb1BmELljdtu2x5
mZP1Q5U3IQc+zpDnrwO4KVYgS9GJK7iBxLyK3ngyMOzKkmsejUtCcA3pxmfHTRad
aFNhPoS1bccpL2hNGCo8tMCIXoNzd5DYjRsAAsbaAr+k3BkpZrbKBdQuv7y5tmXH
vJgBe1AWWZuP24OkJwC4swxT6y5VhQSUOuKKddRpV/0eKr9r9bITZ2IF6D4XXdNG
90gWjJX1d83g20bSvjioGZeXGzDDznL6xDp0DJJ6uhWdAzhhBgrWPTGvkNP+2zer
jtkTS4P/c4+92WyphMzKXY8nLF7Oi4VWF0RFWu2kju5sl/KscDqirrQYmSATbHxD
qkqovFjUphBVdFhalpMotegooNQfQGjOk0BCVnaJvrN3fHNgG0agn8ELepTSWp+V
dZqrxo/4bU7FSz2dvOHzhT2UOXu47+HlbCf/bDxOBqoZMwzmtT34uCUpdswA//KJ
eVMIz39wXGiRM0BTVHYu5uRUFHePU0xCIDtttFeAxXOpLSWawgfd3p5ZjloBKUwX
b4A5MWbOu2ZXquHccmTUapoZU8SA+DgE1cqzQnwzRuoh6lmOMRGjA1H/K9mLRdZe
EohT1k2LpCdwHKqjKPJ84bBrYv8DF28j/cQlpWLQ4HVXIWtdCg67EBDbtNDIjsGr
/P9FRDDmUpX6AffG28nJGkH1zIt8vcQVV50TJ5xYQx1t1tb4IpSpyJSoxOPVN7pw
H5uD6fxdZP90M8MDJL8TmayhKT5ntOk+SC7GABHWmO+nYDt5lEIDZ3EmGtA6Y7x1
nWBKOt2pDZhEouVpQypZzGllt0s6YM7zr8rPtEFqEWs+8FYkek1abOiL3m0VdqfE
sB8sKRD1eSFHu7BYVj4RJjb1rgNVkjCpuNFvy/8NVEpdPv2VQYLwQkSi9A2Nawh4
4DE4nGdbUsKCAe3NzIipp0xMKmQt9Vi106rsiiuddakDCVu9vst8bC4Guw2qH0w/
iGO7NHkrsjlCjinqkURi+Be73uQqAPRFMbT0IqFp5CRNnruT2THyPv3P96AO1Q9I
HkvrzYgy3PN3Zh3SgHstFEK5sLKkofE6I1Gp3T/DtN2ONj8vpHOQLphAEDy8VcuM
k+v0CZnZihqlFmA2NKtqoO2n1DysCBKJiuKzy0nvInyhQQNdRHMS/9qXOp3CnWkc
o+fLjxzMaHMY5v7IQxUw8xjZEC36NeNoI7vJDU63DGsoiekEaIug3rs4sio9t1bK
+fV4c54IePC+syCIHKCmYFWvDryJg8bsqU1jDW0Fcx45IrSakAvdviJEmZb7LF9U
WQS/jNW9jg1VYHMu8BZaKUAhjwxvQcJ7DWVy9lLxdlSpB+v7VWsMqLhhLjCBjNQ6
Fglbfi8bSpfL2GDBg+NJgHKdepNV911+EE0xctCbcy2BpkfSC5QW0C4CUx2tslBs
zTPW020L+QzyaNf766VjRAtY92EsogDpBrpyYzaUDQ2zXWwTz3r2GClWS6KYfRMM
FxpTp3/j7UFo0xfMLxCR9VyA0h0YdKyFQtfakArQqrd2HoWWEf2sMiGAQmH3pRWx
8vfFS4nNHdUBH7m1IKjwuWMwI1ae0WtUmzFIq24DU3kJdS+B/zdbqnzxqptUSSYl
Dm2xOgya+So9O8PCr3V5q2xUqNiWiXbMFt3kTgPS6TkLbccqNWdsu/mwMo2s6VqN
wpunz0Y6XM+ZZnHCrW/th8fh0Ts3wz3L3m7xZ0BGEkkHbz4s3XV4gXYdhu8sGBha
aHlSfIbAe+OBCUxZhk7V+FLs+sGiKhLofWvCsC9cNeF/3tgI5idH7QTaA4oa0FT6
xhcuieDpxxxWz+3pKwk+CpNQrPPzOYKvKTIrfkRBNWRnf51Xn9C8FIaZN8q8QT1p
hrLNjgOgwCGx6lZXjd/yogFPV+dhGKBAmnHAQlOoeMvAi8PeFUR5MC85h9NugKHe
1HmfeZVGlmE55rEUOatz1acVtfnTmnL3Ezn4GvTq2LKsJHXmKxyAVa8yGNev96MH
IUT69fl32RriEP+bQAzUoYgRQGQzilp/Mn5ppP14sydtYEW+774XyHNucYpM5woI
3cmzWixzeKQhPHIx5vTd6NmELIegL8GQmGXsSLWO86sGeHF6DcxVZYaDamA1ErHo
2FTR6Y4eYcLIgkO/w3NBY8AOdXcMKr6MxTp9NCpL4j5Pb+ycLNPT6LgeJMgLzGFj
U6IUKVkR9/txZRGnJKbSkevkpM/00bSE6zZx7QzYKMV0UpEOjfUrNwAwkOy6MMJ1
3ATKyUlPexT6Va3P8UV5l2TRwVhI80OSHQGX4eO1mN8oj1quJkfPdB7izyQa1dIH
c6+6dFm4SzwEmD3f9x2xDD+fyLnjnZqvilt9CVP7/+j4c/h1TXQiUUCV8Zg4IK6M
Jg0un+EhpsCpcGK8DnNhlXl71LxaD730BOy7qwI1D0R9Phpym1AV0fTm06vDRxLp
oTMolbKEIHtXVGDvXhN+BZtLVX3f9gWjJU/8oRLkKX6vnHN7Ea55aU0aK/tT22WR
isWZxIwjSKVQRQFOOvT2LutTZ3dcvjiKzRSOMIH+eSUTVPyQ8lo7EBQIcpyEqlCG
vRxwr8/e0YO1Xzh9LT6OSlto/evvYeKLK08CzGbjhvzaYW8ctDfRGlA+j5U9U0xS
Jyyeu7rrc42HfxvfzfzaHCJcPpQo/VibN3/e6PEp7fZGHPvKIZRiAmCzk4/ggZ8X
41bRlpJ7axukxnEvRO9/X/vwhJYSOmWeLhPl2CBCOSNp7Jhgf1zArsSVaHP6q69w
+EO5ogHorVWGfSVY2AJfwLpY+cYC9nfwom7AKVcVd0hCNGhabo3ytIS+jrIAcwlN
0DMNNaFByAtxTd5AmsV21zDVm8rhPWnLwh8mhJRCbSIfo7W+n5lEBNKApsMjBVro
Xa2s4p1X8E1VmxUKYxP23ySvXK+q2u6qJ/4gWp1VgOl9i+kKSxX9743XIrRCYoo1
wFvuDWb5sF08JkE/pH6pH+rdkQnpkbs7CktTzzrhESsltbICtvlneZIaz+i8UKF6
psXsjlZYaJ0TYZliFlbXx540o9IVapBSJY6fS6EQx5JiXFd7aNM1l8PaHdeWAf4B
O9ptLULZNIndpFdO31nr3uyR7mxjaLLXlrrd8e+kXdHV+yAyV0IFFLUeHKNRDobM
ALpXetWpGVDwQfCetW/VwsGGypWGCJ6dPUjLvqDfXB/8lsmAVgy8TkOojzUiM5NK
s7rfGqnHw4mpnMJ+uiNK/c1FLVyXQnE0yYNIwmeFBjixVojuQQ0Sips5OkySXllc
HmnFX/iX/GiPG+M4R7zeEoXplomP8dkKIZFTeXK70RrTHLgz40IA0GqPYepOBjgD
Rvt9iZGMifqLmPGF0kzdymP6+8rDNOL7jFKNUAFPcdXpGnqKDbjs+zZ/v0UGgnR3
9HCNpHsUA3lWoD4i12roMKYe1xUSjXf1n9qp488nZvURDvGaxphRhqeZMQvZmOo/
yb8d9nMG7YHTp8F1JALOylgGz9gQsjAPWZnGErNZIoSVbp1qm0JvNbtHw7VRbggG
DND+vzDPXBRY/MS1SYrMS5/3odUNNelfwZ4XjV7Gbs/SByRZtqRwBHeAbNyW3kf3
44Cu4s6sxmEV8qfDvPrRv7cS5ab0K1uvR3nXr3M4gPZ93rCKaKAtpUuwIJfWTj86
uJH0coXKOim3zMmalDQl/9O29eHr5nla/KNUXi9DYSjfXXfGR08HDB7AmyXlXd3Z
USzDKrWlpLequJTT6+EMQg4PX7iDbGZgG84PneREJZkJ6VrgV1W2bfd+pHHrys4u
ZHFSDPO0zQ+Skt7wYntGr6719UerZ9aolxD5G6HCEX5n1Cfy2EAhaRghmV10GqZW
R8QxTeX26mghhd6rRdnuRx4Z//Cvy8mqZ4i/7ef4IpA296/d1TTXx9WZOHRMcznd
ifINftBCHUU7q/Ealtu5SvZP1pzNubWzMmgM7o6PAw/gQ3fFgKbswPbU9+w1malY
qgynYlerb5rUWII7fsbuimyNtLv2y9iItrozy6fUiO69kM0532BFAtlG2CqCj2MX
S2WE/QaNpKd01rCyFeZqZEE2J9rtbORY5H0kfM0qn2Mg+mrrYIxte8Ug6N61+enm
szJwmCXqAygDUp4e5EgaTP9ihyxGjIvVkuBZ2elLdZANzrtExSiqUyXN5X7Mij7u
MQFcUTp5UrKSYJ5N3NlgfKjPOeWDTNmc58y55mORrlVc2jDKjfvdd/266spyF7CM
lMX6+Bkc6FAVcjGV3mkPhA8LQaDK22auU0FzA/srCVEtkO+qTLmpipzY/BWmbMYV
ZwIAja3kAVgKmsuSBctOEB8YdqmGU2wBKmm81Rqi1uYviuKPKiQULWsehoiOvbyN
NrPC0CbKcez1SG1x5VeGqAQIZvTNd1athhvK/b2VDry7zFruVasVQxtX7jW2Pnwp
fdOr3DitGxogGwYeRGwyBvhiTBndnILJ+4e1c/JQaYRuDQBhgPHX5j5noy6StRmR
BNXBL3QdpVXbmQYhgCXRw+Z1eh/E6aA2EJDKuyOLQKGzbVdz4K420aOfA/dHNdkH
fmEDGygYydkYBVkWy7bdftlEID+G5XvGvPMwPLQO+/2IW6q01/yElWOSBj2cjwgq
mOIDtSEdRfG6mM3cveWPON8JdpT1OiLXxNYowIlcoR0xbt6bpMLhY+StxBrFdXQe
48KLfgyZDRaKWEQheC1OKheZiN+7VF+C1pplR88tXdvL2c3GU+775i2l5lDppiRO
me3A97vFCIDkNMO5LipkayBg+dWq8GJicLN++Z7beKalDVjsW3asi5g3MUaBNuxY
Ay6GC4nuKXu6LtDGwEYSGGrw8QAIOScTtzNn3qAwvdLGva+nwU15nNZoCg5NWXlz
vVyPEcV6Mj23uT8hNptICwVS14DT6h2WzvXaukqz8t/QR+oeNFWGUa0nXYDc27cz
/VvvMoVHnJBVw3VsaNTX0xDGeR19EB7uNG/mQrxcyUoZJr/LqQ3eoPehJ1+ldE3f
2NA2H2W9qjJe1MYgTBvMeNow9pmhA6K38HxCbjHXcsczJWJwpgbrE9Cdv1xrNSWH
am3fe9Evfe1I7KtDxKen8CM/Qyz3gteNYVF6vdJBllfJ3ft9fI2ZvlxJnGQnxmOy
s965l+WwhS4s7+CDipXWghos25MlxrtTwG/Ag9VFt/6NYxZgnHiyvUBQaboHcGTO
lzB6ZFPl7JAx+QhURHn6q+T79qwkvsibvXW463l0AkXIdb9b1Qd31k6qTmOHLhnZ
Oji3CPmJLCr6nJneTyshZQVKCTxPXtrjHOVHk/kB4FJl9EgkYkpXEt0M6Y956VEb
tre+dplM7/lvkqNRT4JnH7YYbCdb1xavbA1kahLRersiVhXDif33TOwC7iOu20Kr
URrCfeiN0kbp/tHk9iD9VDTuIk3Q3Zm/QhYwmNJSqmkDM2b5HteSz7NuQe8OlNOr
DSZZOf3yi/31mdXFWBjrvEZgSCeJCrXIojg2Ij4dbNqIkY9FzYhpsTb9LbSM8UKs
tKfuOuRmvm3whMJmzkoe86MLc97YbnSaa+K2AdX27LrHG4Ozn/4DBhHQTmLkJMk5
l+bt4BpAH03nG/qFjg9Tk8kJ3qumKG9UzlpdAJV3pW5GBeGJ5ZdPL3VIN4h84RxJ
7VSDCNwSxz84YQn8pLXosbnt4vMgQNeugke0WFBSSfdrjAKZ9YYv6vtL5EyUHP5z
UbN23BiCErZgk/kMB8G0ZWRlj0NwY/yMJa6RhxIWFisdIJElgrTT9/E89PZX6qYa
fcdQfjDVuWZxULbx2dKh/XkYEbqnzRfkshpKxsnlk6+efZw9DpP0W9MpiOyKB4QX
+RpRK9kl07LsX9cxsXQ/eHrIPOyAg375i6WSbdBAD5S07Ye2fCBE6vL6tkqQbZxy
gngx+OeCa8F6JOkMJHaqU3/5ymVCAAuaf/HqAVgTSNzXHYxStP5/I3Dc366CMzrC
2xEieyTeyjytfY3AW9yToIJTCEPYxK14Lk7FLSSTcB2cjJ/TbyCF2Khul39PCFc5
vvPzI0cowYjDUxY1tBHZtTnbRqCTc0LBz75CXaMB1cS+9wdouFXN+5jZSHyIbhKI
DpUWZv9NkmGxP37isZK7ZuTu1EmbyMCFnsmiQ7e+Qg4omSrQVBoa4e4oq5eeGeMA
qY8I7rl2Q6v0dqeuLLjkrVbx0I49Rkd/rikUNnCGZjjcPk+YQ95aOyl3IzVw52G5
nETmId4toZeFt+JMj2Q3ZN2RnXagXQHwvCS1g427Gjo+4lGSgqtxhlBwYgpYcQ9f
leIb1CHeGONsbFdQeoOCI6JCSPAKifRkFGLjs6eXEwbhflXe3OnX3TzAMOsbRc/M
OvTIVG4TQF2OlIB4JqLAEzOohPXPVT0s2d385zWabMCB6ChPQnGoy64GhiwsCbWO
ex5CroIpsAr91/piXxt3tWH9Zc3nkTDApgxrGeYa9KdY+gUZKnVRkRMOQ45h88U/
x6iDGuAaUK0TeI/1TCQ4yTr+t9o/q9RjBGDgR6EtCJtdGOct9Hw1LDlSjx2IQqhb
ZXw27J2m2q3AWobRcbI1Xo1is1qdNP861Q7CdagXtTRnqfOGFK17XBFOzfAcVtb8
fsGyyLcwuMT05YM+KgkU4xOwlH+ujXH4QjexnoetuNje16A561rUQPUnOEmvDiER
l25trQkdabasILzqmq/vp+PxveBdOOJUZYPALDJZ/R6ywrLvb8Xi54YePu2tNcvK
hCHtSxxoG4p8w9EHL83CokQ0CSNeGWcW2OEMm1iUZo7vMTq3iwz3proZShN3hY0n
FUMI3+VOluroLZgZ5Nf5CSJ0h1/jg9cQobpiUPuKvQD5QAxYY2uw2TBA6Ad/UMiu
qRgp5jSw0RwbfHKq5XJzJLUqFW/84EFSMeHFMS/KAWIGRtZ56kYv0CZduiIcdvW0
WCAMoIgr8Id4GekH9oZPxmcY9V3nxeZE04ZxdryYM0hCkVI+C4Y0Mn3D0k5Qe0OO
gU1EUrHAdsoriqLdPA12yo9/o/jjBR+c2oE7OJAIc1/Jeu5Oq5p8W0aSFsidJ138
iYBUDKacf0N37iMpA+4wRrSneWDYDepW39+hz/5okov4r77MWs8VzwB5bCLt6oEw
8j58zLU4gqhzg40LZnLZ7t3ZN0CImbRXdw5PpXqMcDElNWT2yFtyuD1nC6f+Fx23
iyggYiUqtRobONIuSR0gJFyPt416xSY5WS8kao5RmCJ73O9log91ot4/dQS1X21t
wTcuheUThPbvYv7D18l6s3t7hyEJeHtCMfsjcQzuoxhxkaAGJ66tjaBRc722J34G
52zynA56UI1l2aTVHMzoN20imNDp8Bx0tbzN7M6WZUkc5oNxEhxGoCDS7Ivn7Mg0
CAsAU0E0IdQCvuXsA1rwhvz7d5XeaMtax0ojeDo9yybeb5CRcgmpId/4TPY4tyzc
ZSioO+iG0v8EhfMFwd9NYA0r4PrfwK3Ygi7v2hKY9AkDxY/rmjTt+4CSCNH2o2Dq
nJgeAWubt7GmaPnQKPjVqeaf3xmB2RpResDCqkVx5gATmAxy/3qVFKr/ZPqfTDFC
65r9jWnvta65AUu1VGLb3TgTJ2SnE980x0G2i2x6cuDPGeTOSRt8YVgKYjohHuGd
c8+TXZLGEi36Mqr7/wDqkhreZM2J6YfzsMcRvFU3zN6lPF36AhFrkDW27KJ3B6A7
NXr5hIrTF4x5/NB0KzqFop5waGrsYPct57XaLtPHDyHOV0h/c0QqYIfMUDkrXqq6
2DHkyseV3HVdRGIH+vPOp5iaZCFpWtj9OWhCVPA7ilmAE9biPOOfJQ9gQD0+3/FW
NWFGckjEgb6cywOo7Ao16YnDPynnouvLlCW5fbMphLUtbkPr0MTQjt0JILzAoFyA
B3DYzQKlRQU0gyRetZcUqMQV+Hrq0EEiVw6ooD52AryRqZ5PrG/XBRXVYgJ2fqsy
0N+8cz8h/y2jJNuhzV3XQpVrEF0yrijJXDx+puWlxpFii/u2Qnz+UIw1njhjvRd7
2G131aUncKYNAdU+erBElgMG7ECgHtoOukAuKYWP2vdQDLCJAUQDaZI5IJxvx+Io
vztH7PNZ/ADNkfkHVEb6i+xVhhwuPF2/SpH84pHaM4ys8pN71jd2E2gLsegOV5gl
a1z57OG3IbSy73aFtGqUGjEQoRGRAO5FQugC/HiUVehp483ByNLSD5Mb07pnkFBq
z+Cj1PyGeoGY/iWbfvir5sI03FleRdpNnfJ76uId6CYwpep8K1dEn2GNssLHjdym
ugqAZkurPP1Q7m+BDKZwBuEa/UVSrmpoEhQdN+uLT2x5tgx769DOgBqcSry3MdHz
TNTXfMd7XCrr7d6YY5CYUITkPB5uD6T80aFb0hxCvRpVRskwnz9AQJhztdr0Qn4i
m10MUOIpUoVHR9ZftpeB6tvo1bqEKYj4jMSCweVcDDNjyn5GGG4FXcEnmhdFr+3H
iyTvN/QXjPseCreT6X/OZRDXUlFX7yXuXx6U0vqbNfqqsdGogwuJmE4NdzRAVfzR
Y4cS9tiJEjnhAdSG4A3xU2SxdlnaB68z71R/GH421v1mm8artO6Xy/QSmxT67a6b
8eyYs91zkQ3ktGaiZV+SqKof+n9x0BeBXf0yO/zqaO65wkrS2qtbb/Vm65YJVMXn
r4SgEetaiVmBerR2MeZubjAHwSrRBFgzF1eQpWJuBPdvdhEmYHE355zA0+AJosuz
u6/ob/uwZyeUmdKGTBF7olP6N+5zWPsXiBZ+kF3zFv7w27rY4J1fR9MQ49cjqnuE
+b7ETOLuJWNjkTfToeVzDH9N4o9FcECY5CPCr/hzHVPGuSA84iicD5fBD/0J2LMn
Mz0eENFcc9rbCxZZPP4lx6ZAomo5ueioQik9U8T6XgAtUYWKIOYLnPCJDTV2ZsP9
N5bP/a01mUtonVI6T0zd2AYzYpYrI+ABopCiTIpNyHy8ondd8i7Phwup0Y3ml+PG
4aPUxsOvYuHvvkBADINgw0RtGEnoSZprmopW67hF/El0Vzgv7Bq94ski9KmufqK5
oCADtjQpbUrwvkzM2U4LZzaqrU0zc+BZPzq51jTDGQY3dC2g/U8pCPyjleNdvp6N
sDYfjSWjl0HIs52OZVjp1FTGWCe5/nakLfFNSUSh7uFMOBB05ZWmigsxIrKcjiIz
nAcQBjmg99fdS6vo8cd8TsxdK2vg0hYYjzZ/ClhFP18H/1nX1WYakqN+AYxJkB2P
PiX9ZZcXYSz4upLcn6epBr3EaefDgsiwZ5GI6WbNLmD/WiS/RwLQFMOY6GE8N4ll
nkdNQDWVAQOmtpI/znFOBIbTMNVcXbjV0fJggvaSGZq1Ifx/iNOTmQWFkgqCt3/H
x7YStmlYqGTictZy/ka/atDxaOSkAJRTFUdkAYyguRaeLqNH9Y2wrZ1TNOL9hssm
EfSDs+mkIV98ocRhOBl5BpDGd04BnuKy21DEy1Q4lO0kYzlTTh/v5lTaM0Bn7LDj
yJ/PIJnJKyeVW5Wvja82H5h9Rvy9CHJKsaX584Z/8MeWcEa3Ucnyg0bIv2DKYfEX
Utfb9250y6puLtOsT0YOD/SQNFAUSbznijrhdiZ9gsPaEiPxYhfM50qXVsOPjYtI
F2o130VYqRJsO6UdmDZRfrGCqXd9D1WaIib7qKZtTYFWcP///gKbIjDgqfjN0oGi
Z301bEWSvZFOPvYLA6Ah2y3TJ7O96CLqoxjsSo4fteJrnvw+mxOdJeW/N96kILyQ
vFkBLZ0dGKy18Sf5HHQdJ9oLOOLUTFHr43BY/1oxpPOZyb+w2GiOTFUvQyh67Ocv
IcNKONL17gHQzqxccHiwShcp69zR4RVa4gzHaVU+IhbKAyjsPwo3H35jhwaFn/jk
2dRAgZ0tgaYap+uxoB8PyNgZDcHt6eLrMLAYQvGukKrwbwtg/R+1+FMPCELWRo+y
s0rMW88uZUkwGa1ZGeGTwpuwrLspT9PyQuR0Pz3jUHAnflI2ygVo3PVHABSX+zZK
4TzKPOLeNLEkrTvBQhnlfqvxl+VjeTsaM4OWyrz3w2ipMfvOP9meAINZbFmwt8je
GFegB/YNp4zBSqG8MV+w903yZ1INCz5LsGKI30aFcolSP50AKINa7KMlEpSjEC++
IKFSXGSOXVExrjcyOoLXJG2Jc3plHVZ8JET6qPPXfxRErAkCk4LpF9nKA7l4LFkM
9XoWVguIRbNUNioCSZvwmWcgTnnOWmJYsjQkGDAaRNTF3Xj2BVNw7iz9J8rofbwf
4xjz4BczJW3cMrPIN9Q3xkLKttKqh6eaUhbdoFPKH46z34WliKHa79IAWCXoo21V
X/5iHykE+ub61+t1sTf2ktImUUetRIJmpXWmvuUTybwy8SsNJ+UgfGrp/0kfnsyj
V40EdBJAneeL+f3uvuM+6Ny19gQEIaSiTtFooUugrieraedGcJ5jSyKXyh1m7TVj
da2NRXECRvHYhn9DRzRMvCAYyG68qUNCfJ9nSavotfoAUy/QMZl8Tz1WKboGw5cR
gHT4v6YVoWkTA10K8Kl7roM9uuwXH7GtSLI95gP1WosMlV+QIPtnXprh+QICwBDT
zk0JnaTNhILeoCIijwkF6UkLGr/D7u1dLCauVR4aqxNsVmLHHUuW23e81mzWwJ55
6bMc0l0+eLp7wntZmqJc/tlK2B+CJpPkttsJ87M2UwwAEbb4+VHS8xEDUmL2vxcS
66TbMc2VSoQ6rKWiBwQYytJ74mLtszYOEZuzfuHehjBRATkamGcDYlbEgHzv/Q2p
AFo4s1BMOoptxnDfl2HNjdIb2/juwU+B3sH2GQUGgjY8TdIy9AozvccyVtVTsYrg
IJnCf2HwbaLFzFfq8SFlxcTnFpW2kcZt4w7hIZa7NZfNJ4axBrSYAgT5IX0Vag9t
e7INdTCnwU6dlN4bruXTv9qyOgFt2tTS7CITAibOpS/IKUQG7YQ0+6bZiimS4CGE
6C0ebl7gDuqcei4SlxPRdSRe9fCzynf1brudTkjld4g1yMcp22oReEFrZfdEIh1V
9GZfgjV/eMoiJ7adofJ9uHNqW8BVuxtAt7LI3bJaWddcwAvVctWJZNcV68QbzTEr
1cRrjIRBf/1x6j33zEvm+eG6ft2pB+3d56bOYS4Q8bPb92BQ1THqCdfDJhUUx8Gs
Xp7no0hmGKwEyfWtZyTM4hb4myniY/RJcTdLEaTWl5P7zLE/gQRz/ZqiWuuHJHf5
qupexNIw/XjLPXWSSTe3KLXpI9OKQGGuC+t8Q42JInbhXMRrgsF9pHxVfRDR+lH2
emmJLCJSj0Rx+ZkkcGJDGUi7ynfWmN0pmAqfhoiy/T1AcR4TisxCKGGIc+3p60a9
eCCQIuRRucNX0WivRYK43I3TeualLMEzH7nP/uDs0LKZF3AE95mlWOQVOdeFjIC9
ofnvOBg83AxTl/kRLPXEmI7W/xqfmXEJqryWf+rUuFN+ItRGecM6rLecW5cNrFnv
kd9UJ5Rtr1vPp6zlzXKSWzJXl30XHbF6DFzm1clN2uErrkRkoSYdRcQ4kWp0+eoX
g7U1Q1v3aVnPzpeUFnPBC4/lLDNYKEciKUZVzYZv71CA6yJNuUKhQ5iiP9UFvETp
p5sdATMfilD1aAcnvOe4rZdClgocm4b0bMww7UG3tvQ11vVRnUycUoOtfqz2NKhR
XdCKB2IheCyJxhBEyQY/xOPLhH9K9UdZGdKqfUl5RljS8OW3Vq6BBCLerF+Y/TWM
6sE/fZsIT9wVff+qFY9AvIq8JX8PISPBoslAHfQnQIOLGQuX6mE9xm+LBG05+a13
xTQyzqpcir+Q0OMfvas1T2wCcw2/JJ8G9oaiVCRT+PwUpWEc7bguzZI8sC2mrV74
18w16sMzDZSWjWP4iMJT+V9ew+jIaL+RzzzvOJVV2DEFSoRDaE2hfBaJvWqaEiWq
h7Cxbp04o53uyuES3ALGmAt+QgzXpAzp8Cbdw934lb/9wwHEbSu6N8yu3JT8IHDG
huI0XMxDighWysurFppJlr8HWYqsY8rjm1YO5Q9GcVH1t5+dyt4NJ/6XJrCHfYre
qG4jmx5cd9cHwTuCF8GspX//SiE5k0SbDGMUopNC0z0/YDtj/5woYBIp66bfn5IZ
PSUhG3DHKjerEfoG2lHThaweWEsu3brrTkwE/XsTDqvk7N/EM2HYNTne3w3nKylZ
slimPQyrwFhWGWxOznd2GvLhDvaKFGf10+N9rAbFGORr5AfQ/2rZEyfo05QXCkeI
7gP239mx+V+LWEfrgNmqZ/fqlUJAigcaAXaCHmH1aNCJpSpmMkUnoV74u+hdMQei
2OF4VB2k7Az39CRHk6PdQH2N+gZGvZj9eqnAB3iQ91Y6Wng9cXORweQlOOL5SCbZ
A/EH1GC12hJDAGokWfZeXUIMZWriwaWDwjndAwyVjUKtAFCNiUdMDn1PjQwzk2RA
R2IMP7CWXEwy6mrerYPJV+hUsauE5Irm4CFJzNy5vz5Kzars2LHMWeMo9Ldl03rn
0oc/J+X8PoK7op2l99zyLXBgWd8phHh4PmiCunyZD6tD04o/peRfqHfnSu+B51W9
+r56loiq/pdquP5V635gfbGw5rouDe6xmKneoNaGETuUTp2DQ7IW+hzFB8B4WDH9
siLNtjBxKWRNCFPqygeC3AU+o+eGcu2VoZDd/N4J5yvk89+LbOF2egME4JNZYUO6
ES98pZpgaW9Efcmg+yc6EQGduMlfJ5bUCYLe2uuVs3doaTpqtEkvjrNZqR92NObB
OUNv5oYEoZVFWzctfPLiKihq0HbvuUFuk9K+ZlMDXb4xPSGOJur6dlK3SbR2A+nR
5ooHVkV/lwU3Y79TGlOsAue6oooYnFdkHV8ZFScQ/ydf/85uCgETpgiKdnsy6Um0
Y9zNnQXoWnT++mWB6RaOF+9o803siK917Vpbr7xBwRqOYZBFPVDTIAe/x/PGqI35
DsYGRL2f47nnGyIJSkBqENwb7y8F/SQYFS/eKUg5ix0uCYSjlJJ83gGLJsSPjxmN
dT4TIsNtusyEvjuyubqa6+MTlI/M4xK7e+ijMrNLdLZOLxnN/IhgjM7aFkVBMVOx
yycYet8pFh5lPwGPVwdvIEEkZf0ifcuNJ6oQQbYkE86jNEi2egj18T5VBAGoMtCY
h5E0yv+tkvodZbTPcxtoEAPC7S1d6EFgJsWsbDBwaifOhVcCtw58tNv0l59xAgDi
7y9XIFkH+P2ivu7jSzbm+h4eVHbdMB3a1HhNwccmtGV2FyFt237HZtfyZQniai7Z
kTeeNmV+7OiYWoGjJ6LhAzpd23s748uJ98upHfG4XBv4fBh5bu5+35dIIrLbZYDF
TJHbofOCnfzFnJ/JJMWTJefgYn7PmbdBGAI2OmmoI9QiYj/6s+urDO9JEGD9iykA
9lafuZSp1aEhv7uGa6wM2tkQnqaLgu4aWRSzzJr9JajUSsOSaxGzRZCmP2ZUeUQ2
7AMnwmM/OWj9DNHAsaHcXARDUhO+DywDzWuBnquXZtFqu3Y6c+llxilTUH8h3NHB
IDkIryJCXEaF1eQREZyJYOpCxmKJVbpA3NefG6R0xLUNm+s8bH6lMnhw5uOkGWFR
lyOb5I8y/XjH6aSvc7erVwGvSBHizXghZzKQUMWy/q2EvFJt//Zw0901+MzPApF4
jAeVs1h3SIK5y8xWfRxAifY6XiEsXy0RoeUsniKk5zHaRb6a8yO6ln6UpnJDllvM
Y8peeyE9FRgkhVLR7R5j5t7sxUVMxwlgN7wbV6OllVQEHgqjGtNEXZhKeFjm1lqM
g52etSOYNc5mmhIG7TBivGhBPVLPNVCHIdEhQhZUdiFp2/G0LXy6KdnEfJ1HOOic
eR+C3JZDYVyxTnM+4WMFzptcsWjz2Yy8Rx8AAiNYMeKku3N93M6ah8h9vnhXWlEu
24fYk4sDQZ1xiBSP6eYDBlETgp2vSmVkn/A4ueWcgwrcwA5gczuAbUBzXkMKrVBW
bt/z/SBOa+89Qxnd+5BQguOZ/88co8ruD9KKHrPhwn/KZdVtHXJebH2GbnA76VUf
sx3kdi5jtZPa/Q9TeqSue33/qVX8jmrn+6ZJGsrHZMYRcOTU2e47iGLvXHzyDGwO
MQ7edxORq0UUEa/GpVv4YxbADK/P9KNW3jx8GnuBf3whAs5+Ua8a5GUDtXfoddcc
M5dJaQdERzSF2E2zAuTVTS8p8h4JkGw1Rk8t1YvqY0LjPNeW+XXrlTT9s0O2iEqk
qf/3RMH8jV7huiRPqbZljWd5FfkMcQC++5Thy26k4b2pbPAPkfdJb0Hqn6VVI+WP
6sJmJBTPMhNTGKEJvoQPQegh7PDgElFXrMi03kmaoyj+I5P8hvpJblHw1MYvNmQh
sqbBoX74YLJFp7Mev046I2tx9hrcNA2qkGWKBAs8Rfp8C4uUTdYASQT+smnNBP4q
nHHeQwp2Ehz9RFKga0c7qdB8TgIFbHCj59JIRxsJi7ViUdJUdfy2S13nktQgiXZC
9JUMdMLSaPouG0Gx5YaKr7zdglxhAe2pHmq6RjKVvxxf76SfOn7b/xsyf/vmUVfQ
wcQR61BJ4LKc7B52WJ76gYll5lyYEjC5vzJrQYudFeg+a+TzsTt/iV8Gtl/JArX6
WIlBDJI6cSZ0vW493Mn+UP6l3lHl12g8RmxC2ZFdpM6k2SPYDZYG7mIws9ZEWAwU
MBQloujinGjnGMnmFnh0CtTlywRRXMrN4e/yMSR9wNz5O+77lMsS5tJAwj3qpoqf
TlwusBTGVKjR4nUvx0019HeXePLGfnALNMa0zFD0+f02VDcTA89e5mZQNZ5JkR6P
vlQ7widzpONxM8O4fWLR+jCY/fSudDZaNrXmnjmYeRGyqtdfe+zPi92z74dGme2Z
zy5nvsZJZX8J1nBgpF6fiyxXJePVNBgmn+LyJaLQOPH+R1iMEG+/lWcnmdjZTsSi
541NiGMuzLqtHiXTxs6DgzbbnvinP9qi9ldGGcV7rSciPCHjLmBmOWGcBnAIRahD
22d9ZOhmmyztHgsLLxK4OVzB6JHmdHbqCJRug40I2VtgTccITls7HswRVe3qMHeH
dw+gEe3KAPeXV//xUIJarCggCuNgFZtZnkV0c/0Ew1+/HyX1AAxS0Yi7p8MwSOxJ
IHZUxMcLgJGTMbrdwxR4Ww9WF30H+4ssP2KH9J5jX4GDe4aKy/Xi6+bMqbsXOL1Y
0R4B1qBKgF0fCFg4VEJ3jqtflmIHX4cIRDO7KsxT7Xw/wrJJipUmBmSFdlZj7wFV
g/rHCEgI+1bqSwJrByQTJyIhrWBAheLmDFcdZ0pdLD6+Aaj2gnTQuIIvNAeYw6Xg
CZpp98FynlBmXs9/iZmD1u6VR8x3pD7jfEuj5yJviBx8YbvyQn2vrAiUyjn5BIn7
VzpdyjyVCfsBUCRE8zMBqGZss5KpKpHXC82cO2iZTWimzXu5+FsFRw6nfYI4P4+K
hA3e+Q8dw48bhL3QaMY92gJsvqpH2TyMeD+jJeYQUjCG0t6QHGsdA0wlAAtJsYr3
B5IZQTJppx0p5NwNquqff0Xkp0vePXzRBQV1xnFGAR6V/MnapPIbh+VBIV0ECqX/
wN6n+2fwkS7xTYKZsno3yBwAirRJ8RyN3nOSYmvvlV9wsH4SMp/c6oIomEilcBpc
mHlAERPazyuhdathGLkXmoFVezHnrfThiLY8PqX8wiN1zohVXGEyt5IS2N+CUhkG
zXLGP3O3cpekoDVfO/S8681YM44KDGODTPazJ8YfoGPwqIaSIw2D9QImc7pjfdLW
BTxnbyytCcydfBPEZbv1eAZgxAbEZVPTgFDE2UkUK9r350aXzGcn4EbXPvubVrxT
A6EppQSkK0n8s8mvbnms4O39zPJcAr4xbNcxobrE0G7+jaJFhqL6c2FHkd+Orzyv
nmhP709BO0FhnmDxsorqw/oHDma9SgrELp17d6OthK1xEs8DuoragtN8B+HSn3Hj
xmgnPQMwXYl9Y7qVSJVWjTM8PAQNbxM/xDZm9dhEigdaAZE7GSE5XoiSD0Jwsvsl
RIyuh6IvJXMabtAPGAixZ3a2S7+Ev2tbmheNZyhvtK8zRZzZ8Esug6fyRZLTeCN+
9ESoyiqxgtaqooiehzsDyUOrBpUVaQEBNrXqUz9R1EMarW3jWGE9mnth0v82kFo3
HZsxkwPi7ULTglmzTqWDqhiMeyJfZiyp1Zb3XOMqBDl4O9v0wHIZpkLwoV1iGSdT
T1ccdDfLBLGxGEyCNel1FjmlV5kJaXpix3CAy31MGeodmhrl4HcjFHhvhuZZanvB
O5qsIB5ZQ/Q68WwdVf1uixGLf8qLzIPQ+FgbEj467WwrdzyQLwXs5GfII02gwgtW
8THcf8289Co4E0Eb6rediwnf2QNqcwVuZCbxS3HTuhiKf7iEPNjQp5EkIZcAxcoO
n1mgUhvd8W9stVc3lmTRJ1cPMITS+suRvdf2cSHA+nzTiWxJS/ZUEe3EI/jeKXwC
BHZT3VZuXCeaOLqS83ahP8/cMcgMbq6NlP0REbJuK9hGYsNMs3mdT7fKcuBTW0qV
iY4yOz7EEzfE9b52l+IdIcrFFi6Tg+goszaGfvUTJW5sOObw8VEqCXcPeJvk6qZ8
0A3alrPNV2LvDfzcQ4E0MYepMBTG5KsuwdleZxKVTXOZU3dGohhLtgSoDqm3qRfS
hMT6zLIN8iJbQ/4J419rBxhk3KumsC4GHalRD2VLmG6AxlZytkGlzXhLyvCyDneX
THyIP2kJuRzNHUHW+0+3p2tcPWnsRMGRuI27GAYlRvnpnvc9IL+iwoSzm9Jzy6Pr
Hckp0Og4H8meWH/JwkcwVDFMontgqPURCYmPjKB161XZrakToPpDkaNODtTJPZF9
KK3sdCdtIIqYvP9mvC31MZtvTmGR78RtwuIHa0Nn4w9h+meq3Efj21s+wQbFVAAG
LCYbuyVpmoir2Tt1gqtBkXLVhFI6GcDF62aHNqHgBuGp0vD0RWFl7/PXfTZA9Tyd
RFv+XX0V+8UpMaibT/UQyS3Ra9eF4rXgL3xSQBESLGbcVWtk1ZqsuzvTD22ebcbP
9/8wFCFu46U8uy79B1BZTNFg1ERyzZPyBxN97HWIeCgqTkBoYuNFQ7TXVJfNRgHK
jgjUhzUt0SWJwSxMA0hvFjKQo4PifIfZSM4PVigUWnAYUClPPD283hk3RsyaEjZ4
FEsUNvUUSojJDuFSofIUy35n+dtv7nCtqvFFgsrz8tZvmPDmVVDfyG7d1tYii9ss
QNVBuVWHPgTs4wkUFqdWK0LoIlKJpeUd6mFUjeEG0CYVQOOlq3gVH7+COYxLvsgt
SEqXLf7aob/RfWzzNMwOHOYAqE5v74GfIUWUPrKYxbJ1vpqddpj7fAdD8k4BFyde
hl1NE7eLWYn4+SmZHH1ud478WUEu3TYmFujHeetmiEurvKcKLHpsYy6J1cFGQNcJ
GwW/mkiD1Vdzj9r5tsolCVX/peBGviBLabQXMnX15XLAgvUYIOP7ArQz74Pj0Xsr
IRJ20vO4VlIYPzpwCaACnEAoqXknfVEDFQGyo1V0ZphO7ODyTqymSapvIkhwTybS
PlD+Y1Cw4wq4cuEjEPzM+J9Mgug7fdgFo/TH/aEXeT29/rWUnm6rjNbqoNLBez50
Vfl0IVQGPZ/+NQqyzZ+EzvionNNth/j1WMkDjFb6xKUi8Wnr4Ohp9t5JJW8wvdQA
zdgZR0oDkZT3Oq6jLVxJLR+UnTdgFcvUJtT9+R0BXrMhvRIagBC04NVGteVDa+kr
J++u66zkbUHHesDAzLVfJcxVgVMIWRg9ixPnph0Ox2xkjK2XbJTcbRu8lItbfL+Q
Lj65HuxADJ8/fF83I+fOf8YrWwCZFH6pKcMsZwYVbGcI2FAwZ48bb02QjRbDvPsm
xx6kPJ5uYLXDUylNViyFBotcN78DKOp9q4inY3XXqnlFxP+3cvtP9uei5363uLBg
SMlZdbsWf4keE2Rkejt0RFbvKkqU6JqJP4ohRobYxciQ3dhOLFdqP0iNx7A3rGEq
GdhBXkWA0vXeiIZ+u8A59geR8Hz24zIXQ3+Q7yiqWDjT+v29YsKXknqLa7BQCeLq
QkuAX9/qr5ve4q2t+guEDv8kpBkD6QPPuXL1mt11AG/NJi07RIIqzctHCJ9qz3GQ
vgXZrpU9ycKEFL9+3Yo1SJr7uHF8G9+Vf6CrbhD0227BD24KiTWCxgEm98I8dsHZ
OHbQyaaeTgqEx36KaL3ZuYz61wQtPoCwRpobmhX0hsALVNvzmC5Kv9y76oOT67as
LPm1XykOvzvyD18++Y7eIHvIg/PehUfIWiIsM8/7EatVuq+3CjkmLZtLgOC3WwGP
lJB8/cwGYlLhexpftpJW3ihYHB5i8C16KAdCQu52HyFZY5hhq4HapvIZA5/XdYmn
uWutf310K5nUoThtqmh0UtLSsJfFSgK8aCLtogYMruQBdeQVWnZJSLkJhV0SkwlR
XQRjMa/Cs34ZGfE2gJ5CFqdqUnGyKGrzaWFuICh4O9pj80uicKxD9rf5dV2sxCRX
JfcIhlqjlLJ4b11NikR8hJ55UUOvSQNNlcJjlb2peCI+HlyZMRYGrxsHCf4AMkbY
9oM5s78UypPcTnuxUGFWVsVvXNjFAhqLwuIlHxOptuGP/9Z+hTRLX9rIVfTpvxEn
uCdVrSk2IXV3+GpQq75CV2K9FvHVbC2sZD8VhJk2dw+qgAa7Re2YoXyYol8+9anV
ljTkqp9TrFhouW337kxREmMW3t2AAKC6TCCvPIz6uObvpr02VNk2BDvu3P3gJpCL
k/7AEe2ire7ZpvDxjBKzvcbyAIQK00ilMVpYIIgyn9ANTLFO8jFPBYl06mhuEJX+
bLvVuHO08VryWXaOjnYIECkTFD4GeOgnF5WvAw2ulId0YxDn3s1mmaF0G4N7ls8t
ZbUfBLPJBQ3LKwAvnj+Zrwxnr/Ek2RPP2aUwNsrQwpZXJuUA2eR09eFUVVflhpxu
zAYYjvcPBVZ32ljz4JFGJYnnTjjdxSK0TPPVLF52MMYKqfP1y5cKdCRd+SkckvyI
2nzDNvCSNaKSa83sjcgtacgTQPaGWPArVN1mNU2CPTXrhQk4S6nmO7xOePKTZhEv
PCLwjD17tIXNTujNG0UrWK2tk4m9zdXQ0pa9wizMNzy3IJaPK72MtPTQ1rRENR3f
GJVtPMwMk5PAvQI87MAzHys5hfUKe6zrActKZTCgS7CjqmWmmw2ivk3SnagUM+0q
IxlL8+pIIXAFwD9hanrR+9K3Qb1Xo2l7UGYJTmZYf/EZxRekggXaiv+kfliU4hrK
xpG9NcTssyb609J4YtijS5M4QERGLawp9Ru02xGsaWXlODxSq9zzHhQ8j/Hc+H1l
T3Xj5l4WXE/8T8rgZBNY1+8qS6sWHqguVZde9bvWOwN6INDFrbV7JOzr+xu9e5H4
5iIr1Tb+PqX7z9wWl42L8/AiS47cdA2zZ0CsIzYm5uLmHlkf4SFrjtSTOOTqPuji
6ENi4Hv8QDaLBgV0KqiBAgfUiTsEIMHp0pSPbKYxgRevfegxhojNBgRMciZjyGO3
3n4p4Z6tsHS/BHknmWumbq0ZbHQZ5dor7svF50C/J84nlhcB0BK3Dy7tXzDlKfnK
415p9p2cMO0z0iTrxFZkLmdslwIxM4m26Jw2VchHx6NzMokr9N+KnYeO2zvacAF/
f0Y+LlMpjkxUF9Xlsc8P5GQ345ExTtYtmIR9MRFZqLRNPLsVsfOLBXoMdzfsH6Kb
+xQoD+ygW5i45fA5NYqhSIEadR6xQKV36hML9oFK3TH8bWhxcr/QMQWa/hi/hENT
QSJPWlPUrzTjE7ADcsh7uV5pxiNSvt5Ao4GaROxsuHxmKeMKyUIM7p5dNZhuC3Mh
t8dpgU+JclZbUv5ThRswvWQRm9oeLShcoRXaV3rANn7kZRVlLZV2Zx7wQbwscSM9
G0vnJjeDmCdPPU0cMkqx4mF50qPBA4dLKWul6rbD0SdK490+CV/PO8OM8Anhr0wu
X3pR4D1is/+egA7rfFcQ5Yh/NuQjulNhgSyFnVqe+pdzoll7ELUFVKsBU2kn5min
wrT8mmng2jmMXZsppgjFVBDJoUy+1YD1tcLhrpwAEr8kAToJVNhLZ2KP4pG+zVcp
iPKQfqhfkZ5h9VKtDY0ceWThbgk9qVPlRUXjxDd90J6suEj/aaZaPE8nEXjbOvgn
QHD8JEVEaJUIPivqNwhPaFSRzhTJeHSOSy0oyclNXmkd66hmGcDywFoj3Dlzbeif
gsmmuVIpHMKGXuBG39E8A2GraI4GM46wZK4umLFMQ0AvJ/CkR2+YLtIGBv53egcI
LP3kodfSs73LJG0uqgKP3YYFQtx43RCHB1S9/CTfWN/Ipn3rrdNjw4nsGBWAS83+
a2ZrwcjiBiaQ7h4eQEIK0HN4MbIMXI1yGRhvnu6eHA4CFVp2r8OcrDA7UTTpmIR9
296BMIVSrJG+0e1fehfMvVqN6naujaAzfFQAh46vPB6tEmeDGbsdq6nQYDse4sGm
1YkbuWrIV5Tod/qO+FxtV4b4T0qSVHe/OUZkDgB7Us7lsVXUncxnyLjk3OgbbpDJ
hYvXttTyiLbifR12w+eojFqOdJqq4CqpWFoxG9K86nVr52CLxx1rWCAQDEmxVVRr
mCmmkRntE1DdD8xbiO7yENqGCiNzhDSnUItauX9AMLE0EgBR4E4JxVKpj4hELfVD
v3kHR9NNjUY+L7xvgPROevmZXVF6W599gNs2GKCUX3GGmBw+JQlMvjUDfH8Pp5nC
tkPQuCMgAK3Bl2ALRpYq5kKsWeRQwlVCrkQ6V47R4XhIpATVSaCM85ziW9kCXdeY
BsjQg3cj+dlOl/jI6njhrPjOGrXBL2bBtRsRTdLE5Od89S/8kI+lXkUkbLP8fU56
TuTY3KqE5a52vUv3CRTAw1udy3PPGmrUWQs5JMHINWIWCACkponYaaSuTy2aqP3A
Q/dHns5XlTf87JrtX3+1PKCmYrWNnaNyxC67VKch74Vg9NbJhxuTZyGFlWqE5ROd
0oGF69UidNKCMyiuAU3p5te2AkrKWIm8cQtBEv3X8H+NJCe0lqL7Xo6lmssK2GiW
XxG0vyBtvi7bDb14OK39EOuIE89dNgXlIGmR+A+VW9sSIQu8jFAKtyLEHjr86ouW
yRVZXqf8Os4FgfuetVp4ppWoRmDFpDut560/pUlr308ouMwmxXWafRqSdNRJ134Z
Q0fFPwH6QjJeHnUBSgv+/DWekA+rsnG8RSkIqI9G9myLunWfj8SbHDy5tpqmXupn
e3UyCWyjUsBoLm9o516T4M2GS8Hdc3pb4mP4LPW3k4bGlOfr994uNs/fCicH6Gy6
TZryqfT36MqykpoW7JhvtB+cr+h1Skm9ZDYnbRYVZ/lFkAqPe6srC2X/889sPedA
QjD3qLa2IsU3UWx6vTQWJQsSTehv2dxd4eKDFpZeT9yAOimhmJVkIDKParyuAehc
Wcs3POKZ7GDzJuXmZAxdRzygkhAugTLGeM4u1Rhafe9NR3kzYnqwo7cbk5AcqoJk
MdpYms9OZbr1bC+QdAiNVXGHVpDl85DdDMvY4HJlnMaBszRRux7ytzDM7NG/ngNY
yIBvd46MxB5g7UlUYcoFu0GihRCamKWFIDXbC8DpMRkfSkKaVm0AtgINmOMcCuJb
qUsI3kZnRDNDTjcU1+KKt0aIr4YEwSNRFhKhl41hwUI3gq3it1a7lB+Pl6+YwROv
0LszVtZLWvdhpp1FW4h9kuG+5jHIP83C692rmvngMy82P7SzAnXCtgjgTWzCl39P
Kkzr/gx6JgukdL69s7zLZtmUVN1KN5PkQQL1cX+5zlsSyT6NpGVHt37TEh/pgfjR
2HjyTpRbKopL3Sg5MI601acDDGJQdQTHfTBZS8KriOYW4rB+KP0xNZVerQpV1NpL
DNV+HTyMJzvct4yEicaO/5RnR2nxhiVoF+iByQij/wMopM1CVJL0F3SLj6/rbNhT
TT5ToxLB+iq6iP0x6IBSyS/QbENe+DJazyPPPRjHjBlipKZR4rp/UMXg70E3JiLm
HNeu8ZtR3+fp+zGT17v7PO4+cjJmzmje5qETAgJE3tyqp28I0HxFI4LpBqkdNFAu
/VlCX/Nayyz+92pCKtt/+gj1XRxzd4DL9xDO4aAfGwnD3Y3RRLjGEwlEk84NSGbc
IEm6tnrChNRi0sKbgtCqZd3SnI5Y+2GeV63jwiyp4eoelxLzbmBUHXetLs3eQVPX
2LFPY7UMqngp0bRR9LWnb5ilxE0vTGGAOVPxp5Al6PE4t2Vxho+GdJOAiY2a29oB
sPL3Z4ld3lC4bX8u/bEHDLJr1ET4QdUXI4PclNfndGETlagG7k6j85VS9x3NSvX5
1jvsMFMET0zazp6B38uhtquob1TVJUSfFtqAEyCkTkjV3Vjbxk9GcxmN/MlNU2Vm
C+gLhrljk1igYe7W5wJKTwqBRe5pt6lE8MJdIpsdzgDgGNviO2cOdfoDzvsTy91o
+jMNM/gNVvv00lsGhXK4sTlQs+tEag9bqtTwgpeQzoBffWoBQzvYY7MAgrvKuke4
dF8xTDdC69XMIQiuedmP8k4F7xsN/y2HQBPuTKLZaFi0/qcCy04lrgAg7oJLGy/w
QS5ZDf0Jfy/eHD6bMNalxuL2ffCy4PWq/RvjOW99zb2jPgaRnQkT9JWu+KIRwNqR
lNWzOQ+PhdClesRB4ggdQZ79Yv2AZyp4AkJsPLVXo8NoASXIK2Hd26ztlMXdyTxt
OLuXcTDj2c7rqLPOvXX4S1a6gt1pWx1QBAq1hDv6ManShO5Mq1rLqqdCgXSY3fkO
izhEMWUq47CAGcRrWdwV07KYE57LQG/e9Hk9JhG0+oiE6HdwLKDosPRuUGmaRO0/
un585+3BHutDuvxMLdSgnzsU+URb+/N0mVu70/x4ksTPQAxRRqlMIzBSQ78RcZLi
w3FBCKhdWc2wJp6/xbZbZr4eDTLaAXeErOqXdkJ20Kzi/7POAj5UKZ8uXk9hsfqF
/3a7uasoYaldfQA6sSngDArBNCfnYGJNs51dfjnKZ+G61dBwxf/tzQ/MujGej+M8
KTv/5OctfEZlODN6akTgaSltY98x3S/niTn5ZsRMV4ZyJMaJZEn3t4+Qg1S8NzWM
8OJrJKYOjvlFJ4QNjyW5iwqZY9pYsz3a+KUU/JJb+JAT9oYAoQqzMHTejtLT9S8X
BdhCx6RPR4V0zt3YK0+BZBL7anAjlcFyqsPS2Mvx9t5/Gvz9i1LpUjNSb6PwhdHy
Zx4Yb696j5MV5zbBtTT96iL2NeVnI5x2V22sjBto+FR60J9M/bT2lUsIG5b6N7mL
0gEp7vb9hkozDMFiSzSMls4cUHq8kZK0yIDxzlkdrmV3umHhkQk7ih0YSEPIryzV
H6z7k3nyFuY2vsvgrryaG8OFRigZ5qucfh12LFZRO1AD8wc3FOVxFmL+67ETgeqG
Y1+hJXrVazzCNSZjLXLVprQnAw4LD0zkdOnzhienyXxmvw0EBNhIGIKBwsz4qPar
YSrobrBxbr4hF/AXJZipBZUCbKJ5gtERPnUgffql8sniAODLiXh+0YNGJw9ftPdc
WMSyfSQkInAK6AMYL9aqbu7uQ/vWmOTLtW0jswQVsIcRxvUhGsm1wHYfQ9U4KBa3
BVg+QSM9Vu6nkfc7qaq7X2ne1ZaUdvWW7S6btAkS+PXcalNYDoXoEwJE4lX1xwjL
ZlHjkn0i1HhWknTXq6XZvqvCVr7z0lvqX8I6IYeAyQ/uQU47FzITk2ZgtowIUKY7
2i1qwFSc55TNdFUWnwzwSV35lU7SujDEDptABLXUZ4aVMjA8Y+iJsCgWRq/ffk47
NXZqwWi4aspJtyeJtrny6zASlZD/u4zlh6U1RrIOYkwYZC/l4EFbK8McxY23h6sX
x6v93zIOUVhiOlfDHCCruMlxaljrDvSzReUkatdquQD/wHhZyyRzD52+aOAw0OTw
+J8o5i/x9kUjHwPTGjx3AhJiT+COeDW4QNyrpeN6muLUQi3N6+bbJOj/sOCOtCDi
9Rt/MGF8ZYgYIxa/ihaSTKqWrFgME2QOIkxeHNiCO1dm52P1MdKahRan+5aALDiK
wIW97uT6bnaIktZIHfsn2NkiPexHwMRKLcwu/SWtSIRERVjk2ALusmXjhb2Xnjnu
rCfW/kDgj+GZZaK9N9K6sbp3NoqPx08UWKRRARI+wOGL/6EvxBjrSzdGa2UDeLhC
B3kNyLZRny68V+rMC72rK8hK9lxUWqHxIQ/Uby0d6HL1IE12O4IKa0H2i7aXB6Aa
rVAMbHIHEFEfccc1wt0p+YQXEBJtKLAxchpPqVoiU8n4+gIP1Frm8g0gl6iMOoZh
Fkq5juBR5/zZwj+gQzWOBN0ZzLz0v5Ou70c5UA0VR2ZEIT2QfuMyfHwx3eQSlTqj
CczhXY/VcFkb8ML/U3XLBY9wxY6SkrXgYB0fU/+cR7q5evWd1Kxr1/esFmpGDb5Z
iw1z1yBM4ZmtNuPHyHBADkWssnNB8xiNTdThYVk1FNS9Y6Dl3fRbMl8sHtXiEeZW
1Ity6gepPylKTmB8UyrHCvjE9ssaDB30Lcbe82vJh2we2ZZxMikSmI1dksB0zuIf
RSDMqjpQzTDW/mRfpB/CWNnWGzbAfO9by72jg1ol74WU/9Sy0buRwPJWw2Y3KK7G
z3QTNoaCKqDoD6+p89eSORvUylzEtNOWb/LPIKscYqsCWmFM0h3UDHSaUCVtwej0
7Rqo1YcxXH3i59/uVlriAAO6fq1oENTe3fEbveujFUg8dA6FDr+vzQjFbNvD9WrF
eEi3BJeCBhTOM+kk60nVv6ENGKFt4eICQG7lRCbwc7vgEAXMi+8PyOXSk/gXvmV4
kw7TdUHrusB88wMfo80BmqPZ/ZS3N7QF9oY0E4UaP3LlvokfPLw4JA6i8jqCrQqy
jTV3jAdkj32hG/D2Ez6EM3fJhyKRwp/glzdTctRLStutbFZ67zqUGkZiAFh45rcm
tGqdN/RHB3+5xFLKzqQlaluxaBNHk4PjRCv2wtuTmbbnJzoqvnK9P9x1/EAdcoDd
NzsdS9HsZcHoIt+/EQ2t6Bygc8vBMgQO0OGgr/rkh1YM0fC7DyFqHR7cxdrpx0St
dskuPxjkEFtHeuOtCZL55LmPiuafPpQ304FXHwgXfOuo1vhf18j2y+eO5ScHn/+B
L4maHWkBmIRu+tNY6QVpjlMtgy5y9Yzadrjj+/N13SgfzIqE/cTNnIVkHTT3RPj1
arE0ZQUW1mWta99uHcXGR5uG/w4GPglE0r9idHCaSwGmfMgkGtybGnCzHhcXgWnd
Ru0D6vFyAS5EX/WZyoKJvNcYE2eJyPk78HMWJbyxsrz0WS48uw8YJpobRo7IrdMH
WdRrfYALFrQWP1prd4tvnifBtp4r+wak/XtyZucLmxbgaBZ6Ja9CZM+PinKfou0f
v1oXy8VCBBuJZ3HHsoK/NYaIjBaOd/rWconE9IZ7cJpuZOHfuDFXmB1S0hRWtDNW
JlpBFIPIoe2fRpo4qciFBE2DkLJIBls1IfRMxvsY42uwGJHEeZTXRf9m4DyGeUil
DSkhn47Vh4Nfq+misUciyhmADmqKUw3YuNgZH/nBiyYBC5OTB0SkDnZRBVzTnMBh
KE0/XSFMQdFmJ5dUsaroPNrQdz1TTeuzWNXwKHc9BpGIy1N0969kslB+o+nsv6FW
kXBhqKV1NUFb85rw5PEOiGVRp4K7IZkqTyDLP3nQvFDKOpFiAfeo7Wqmd1sb29L2
aYUfWFz/QUzJ+ejvSI2WYoPERd1w5jZechcNfu2GrxjAGeiXvoy49jQrsYGoZk/m
T8zREP/2CQj8Sb9hjskja9adX59ZB5IqdGX7aKhKYkUJcOLjWNAMR8IcJYCPWZHF
D7TApCqTFEdg9KgOCxrSKGCfEQb6EPAQzI9vVxqHVcqIr3UC5cFdW90F3+VvlCec
6wqVtAWY3WURmhdXBfycyakcQ0q4Oca52U2zB+UVRQreWub5H1QULJocAdeRANh3
a7z36RD8dmdeu/j+A6FMFhs8GNaEFHdKsxGQqRKtEW4+Nk/YEwHEYmTxvqvF5ZnG
Z88DIQ/vyXiuE7L35C7bxv/ZtMtPn6b0yzo/i6uX2thjhXW7hvlLIce9YbiDmgfq
pgxsgSiGeMcXQBXzu/+RyXWYYOPf2ALFU/Qa2yobFCa3dgsC1JqXnBfsdMBy/VSf
eKjWdVZiiCx0nvqSyOJVxzMcTLcmpMh0zqm/tl15IHagAmFPbsdDSAbGHBsTqKvq
Hf73PQNLjlxSGn/2pgikPKaZdLhlS28joBBuIfVpM5q360d73zmiKeOcrhBm5ZnP
Okx/3F0IPkh19kIcmEzR7bWZTIb3DUMr1KGbojNK07ODbY1BE6e27VehDH9OIq/6
4iRzjQbVvPY/ElyFfetdSjsS0jadhloKneUeSOgj/hdsLNjR38+AIv+nFLgl6wKJ
VxV6wNz8kcfn8H+xmYaNRttBfB0Mp8t6VvPqVZWKwHGsawuHzNZx0779jErqM9Gk
FhzU6md1NxgHUlbGDYepLoo8cR1BUOu5GORjbD0iFHdlYHix8sonpXlqLjaoK+C6
+r7XvNt/KOWNtL2wCdJu629+Uqn+hOZfDRUBeQaYw3uKW+SjJ12XlBzK4K47Xmt7
PphFcje1c1b29PCiens6xYPV1i8uhN1OSQIMHgqH5oYeJ+/YMpz0SWdOHrnF7POF
I08ARBn51VhK7Laki7xIuEgi13l+lznB3nvD8ziRB4T2rdOP1/YJxIZHSBVknlbn
n+WCjDMWvc66Cs3G28IzuxcMz6HcNavMf5tp0YdRQLYZL19nk87b6OIKRqp/5Z2N
Q0zDWbJ6TbaOPl5IduygNnEY5/isH4pcWZA4l14Z6wJiQbB77KC5tK+zc79MfwaO
ElpyZzIAPsk6v/Dk3Emr0ufSFhXNl/eDqC8vX/r0iV7jtIQsBjJ9tuW67ecT5qOQ
XsSH+hEQAKcaQ/vijCf6BI2C9k/81Sr4KqXxFwDgkttlaBhCIwyneu5ga8Hx5BIk
HxZ9bd52D/j4S0JlIJh4NINnyMFeLK3dI4HT32pytEBhx1yldmPghljm8mVR5njq
aVCkSXJlKZGzMd8gEt9xNeOdhkpQ5k9GhVqvm1k7nFksAZGw12nqPwvrAo4Pv+bY
lj85C3E4JycjeV3MzZjvuLpVytXw9s68kLvmSp6wG58BKnfK4pOir7P6J8dUoeI0
F7VjD6T5fhCXhC0nuckUNfsBFaEcx7EA7eXIJpljADZLlRSZ6xdaSDiRkqmaWNRm
zECgFLEBxsgp6SqYqCAlcLsKboCSBuqNvg7srjWdDyJKOMv7ED+atJCT0qYhJAMW
1kiC52VkqMeRxT5MNJCM2ATKQqHpGSy77EJOmJCepywoQvVcWNKw9KqrTUhdg/LJ
INkpY7X4PGIuvrtwr2bPmTTUeYH7g54ai541+mWqQEBHo50E3IlbC6+lQlegRm61
17Owuw+bgrl5Y2w50GOMW9KNcDFGGJQG2kfd3nHvTuCs8ri7J2aaHdDTIhF/+IxM
mMJW+p73gP9C7TBvWQyXnaXb6HAwZqQaFrRsL08MZckc9sHlHGmzxuosqi2da7lz
LpPlqGzA6pcf26GGukyYkTxDxxb5e1URXhKsWCR633byAO5nbXQbNxgMpoxoomoa
9NV9Z6A/MFUEdG05c3S4xN4k+Ov0q2aF5BD8tdsiJRRf8sldNRQOShrcc8kbagLw
wMHtBDVCc20OdnOMLz4cFT+OnBUjw/BwMLlLg+KjCmR5ONrQf+pxhzvJNpLhSKR1
gFHsQz7tB6eeIDRZJzuVrTUX+D/p+TRroWxlqEhLFxzebUWUurmpvEpF6pWih7wm
okGBuJ5OHhrj7cS85RSsBQoOSXMJaFjEsTGQMSGENWc=
`pragma protect end_protected
