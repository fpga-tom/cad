// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EMKaKWDDo8G/DXFNOyKrlBnSkHdNI/ZKeZ1kBHT8TKHExrQ5FN3m8eY1WlkZuXDV
C9Ym99H5tOQ60ZhaQ+tT8nOqvgUyUj8CXNHIrafcXBSdilWRyJfUy6LLsu8V7jQA
yuvIdULR4+8VET0tjinDeu9sMs/VHq5oFLJiCl9Hy9Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21680)
Zx5yzDyLuztGCpkSSqR1et7MsIWm2guRpoqjHzEMDJj9P2UU1usCbutiaGyuFerU
RkW4zVCuYF2fSDyyesQ8iLLhrNAFu280MspHeWo4s9baoNRiSPMGWw8vWYmVTZM2
0pXIEZ+sOKtuIJCMegh5g7fxpzfnXQCr8iFXraEuRGjHh4ue7/Oy3dlLbj9oMpO2
6aZjg2IKVhharHcH7WbYzNm+9Ui3/oDY0OT7WFd0hx9PaHTmHzI0qOUbg6YXMxWK
t5KQgljbTBeAg3Olb4oCCrzd+LnQQJc8pf0mjoFFsiQELZVJw8eU0xCx9Ge0o0+y
LYUQRClC3Td3+nM9MzeKr99paXHXkNyIoDNp2C06BP97xk/vp2ZFk5D7g7JW3WB9
5kTXC7Bq3yDfSgfj59OKoNizEnu5kteL6ds++4bdxzs5LIE8uh0VwH3gWFPluYKw
pEvssN3SgIpOkrqjkAGw+SWnilY4YH4u9ZCCmSCMY6EbmHIlXzlqvnrO/ENDt0AU
rj/p61vWkF/3nEJX7yMAR+9tdRP9o99hNiqjCUXZ23kpQi6D55qOsGNFLHelSQk7
CcHKiozlEwaoYkzA5KbkrNUUFfA7C5K63mMKB5m0DvuiKxT5NmiTvXOpZqdLIfoo
cXcEne2DLLSpPlcT9bxTu6NH3oz31NlHKwmj+WvPmjbVVHAWKFSrkod/ognTzHST
/Npii+p0yECLt29d3arwLTDnsq0JNVjB1DxIe4aDcwRoIj060Nt74xMkDVPhcap5
ZB54/sJyPPSJhXLerVjeLMhK/wRCpLLj2jYKNTHMkM8FIELLnQWVgqmgjTYi0Xi4
Rs2553CmBYIz/R32lL9yIQgQsMvHWiwyso3+5FBS7ebHKQWEZHSiaq1EjPFC/FWy
4PdPipQt08S+URzX+JMMZzcvORjXEJfRz7iu+A/HxP58beh3JkJAliTCJrKa+ROy
Fz6fBLMPXE6jIe9t4berBmCNJR4nz6d9Rq4GXPIS4G7S+tK3vzqbumf3Nh6fyCRc
m8nnTJeBrsEehPgM3tV18F4fOqUlFFtT9fdJrpjxQaUI/nt2A+NXKCaISrMfAebf
xFfyMZzNHpHykri5colIjfc/ItExbdVUyucIptmGuCte/ZdVEMtvrdYLzBDC9ZXX
+xht+nuppUizMzC3zUkuuTmimrRyc7GKiL/hU2L8u5Rwz4i/qAuoJjmBFS0DeyDc
LUS5NzgjlXPe37Z+Y6T8z9tnkmnz9cj1F6z7rzqEdFoy2XG2wPX/Dhi3Y9IZLK9J
jSuBKu3D8ES+swwUMqUjt7bVlTDu3dhm/2f0vKAvsIbJNPYdfbbXmYSWny8EcFjA
12UsY8R+i5Zp87wSfTkwVBpQw/GZnOcdJ7YqVs6UG9x63dWrnrzr2d6xWzf40CWt
uM4gkKMHZ+t9O+nOzfrD8hZouSPqrVvJTmu4xGtPDXrDSX7DJy6tuMrgkvbznI+n
zLgXHA3aTISlgv2VUsOkcjE762bDW3qbCVtxG7I2T/D0Q6B5KyepjZ4WGjliNOor
cpujo57d5x0bC7Bikb+3qon2dYRep94kV/fIh44v4DOdi8yZY/GI0EDcEVsPFt1F
fBXVSXG56d+VBg7dS3W17WDOG3XmKK1u9dWQDkXcP/vYYDdyi+59OR8igGLhTQSf
BbDtDtzfHCgDT35AMzCpn+7FHDwTrZBjCiYp19c2wkW+nyC17e3CrmM/jBq9g38k
uul8xsdZ23W+5jOIImkINuDEIqlj42gVxai3k29ssntI5DJT59W7e6Qz/ER3ZyE4
NGCTp9xefzCnhUlhm6soiSiWNE0tvPIhYFaBzD0570od7waLgpO/gOKMh9YqHNuT
2B17k0DI/2IaYI4KCZqZhh5eFwAFX8pIZqKZP5AgQLQOf87bplkp0JMwUmsfQxfW
zhtSdq540g6FxccZoE8jWjyAhzEDou9tQ4ZYnrZCu9rQkRZeaZYTHVNtDzn/LAxA
FLlb1xRIy6W5MZBZZI1ScZLfJH3mQ7vG/0vW/aRELs1cHHnHavMC8VkJB2eFSJ5n
xvzO/+49XpNf+fanZsCgvEw7eTWBa7DRxPGQEv045JLQ5Vs1MR/7+GbRnH3Paydj
nwih7RgyHOCjFd7yrhnRI2iqmsPjRvHx4dOabAXA0gBOA7UARWQ1/ttscT3JyTj6
fMG2IC9EFPIWIaPqFzXJHDMN/R7BEcAEFSd49TKMZNYZO8Me/+TFkhJHVFTZVCmh
BFoF4MNN5TSu2thg7XxEr9R6ZTMIHzWJ2zMes3j1KxMtcnOsQqISuru9C49YfZWm
9TTDX68uiXQMWkZGMnmjE29uzEP5ocwl7ekUVZpwoxQl1gjLhAY/48P1i3z2h+62
gGyumCgYEn4z7T7ipCR5imqvTnv/kH0xjLiHR+EZ9xP28jfNsTKngN4xq0KOiD/f
LRsFoU/oOJp0GXV1Rx5xUNbgjEIE5aELHcLMk5CondLrCFOK7DWmZ9z+3MDVxzeE
LJeJCnQtewwi3KYgEUyGOF+Ihv4lhSNCc1pDET+lY850IC3YjbNN+CSXPyE3rXuT
YyelCU7O1WqLcH3gMfvURoV3wz3qHvoQ+Y89Cf+0quFHgll0yuMl7P1MIS6SvgcQ
cj5Z9XjaWgAXrCE5fz82MikCxNXmT4HV1dc/uT4CxkkaP4W99VI0skkfItiiovXp
NwP1w9n0fjx5unIwXUKgmpDaE4IZVBxOb4WHalqtEGEt2Xme3kmbcUxRcilvKcIG
GzauBVWpv/yueASIcwZ9gYaoVduIzeVxLMCMr8lftdKaXoLEtRVh9d1GSoIZxqzS
D002TQP71Xb8q1FYBZor7//cDsdhKebWKlGJrrzBPR+05wENDShuxAsc2NBr05Zd
DgdoYlF5TKzQyPdTEq56Q6dZuw07cGadcrOZ5G3oCJuWrxSexcGIK+VvXbYvgwFw
gCD68sBr07acZdk2T1V3QZ00+k8iqVufyUXYHD4riGPbu447CRfzsfWEiL4cfKII
wGecVBdy4Heb/drsYCTYDMYbcEjaKVuibV5Sj8edE6s0tVuWrAGD4f0NK+jTbQZR
GowjKNICntwXj7qv3rQdnhHDiQNH98GEapdo/INGcEVZYlC26+Uv4+U3plTaOKvg
VyB+W+D2XhJvE5lPk8IF/YgOsaDGh/tNmzLc3ssZlR15mdaMzqmp/tw4LbF4T9Mn
AOfC9aZbhpSJu9fow5bfD5qMpuIO1MxZiSZSNPceo6nt9pfcuHbj2OxGdpy54T0k
uIvTJ02DbQTTgs2VaRgEPL7jr4bc6Le4vTefZwES9OK8OpdzwoOebPRpNZxSWFPs
XKanur1tCBeZTDITaPT1qNoF1Q5qxU1enLfBontKmv2sE/8GA/ISE8kJrM295DNJ
x1ArniLpx31RJZwnL8N9BQ3OAGTKnegELoaLJgecGthWLrRbL4WfmpObPxBMh7ss
xWvpH+V3i/ZV0ISdsu5VRAoJK2CUavKxm8/yMeIQcASYpouAvQEPya/swEQj+uuL
I/KehM8dQ7dfLt6tIk9x0tWQvtifl9Osh4REZJLnixhL1B6lLsRsGOgu7I8ikPH3
+tuz/2ZvHpulXQXrZ1V6Jd4PBdZctDA0DHG/7+UIRfAtLw0cyepRf6IATc0O98UK
u7KmBX6K/Li/uuqEBn+jjNI3kDD5i49lllvN0Vf1MFXs5PgkAh/rkaUOkA/owXE3
oUHTLUj5aVrvMjJ4K41l7csNgse88HDsXJEhRyJbMG9N4wCz/YbAM4DbSgb25sKE
Op6YCipypgdilOcPHIcGPjwx4iTaTn1VZevWJlS0+v1yQv7CzvzdZrGyvmYUj4q3
7iqNZmnZ6IyhbQmsh2MJguYRjTnwrC/cLrhirYEbtDImCAYczvd15a5Sk5+RH1OB
SQnFNgqcWgns8R/CuBJ3BNxtxQ+jnL5Jm5cJrTM0TkOVLcswADMwldlAJGLYF/gq
xma9KAuZDttJPaALeK9pngNe/bOeg/7dV3IGoxyMh1DuJu2mNTptcvSFr5hWawu/
Yxm9+dBp2oobFkPKwwsxJG1/iko4H6mXgVpXU/N2xkVrk2OSQd1v07wGTRjWo/qw
h571oVaTPowqP26ufyEBu+0qgWf59he747sLZCsfAiLjv/WllMdh1tLJgR83pK/4
P+vCAKLzBBkfHlRdqTLCrZ31dH7m/ttfrskLr7EhbBkV5m4n51kRdowipUs0U8zZ
n4eShZNQkIOQUwuIKnKeT80YnynIVvGzGXX7zIETNaXI/Vuw8ZWuK4V8basOXYuY
bQd5ROPgPoa0dkSass/IAPlxlb21mrtQxSJ1KvAAu7c3c8OvO7pIIf/bWDNcBS7q
JhV+QSSyuIBwfkz3KVbpiYDveoB/IfNWvNca4JDvq+N83qj3eBvczw+JSAyfrGye
hNLDZN/4BFewvwAkXH1tC8I2fXkS/1sW/uQFBJjtMOPIRi6zD27WZProozpFJ/Rw
c30vfn4fUHd9/LCf79BqMXRQc1J2dc4bSww7BYgMktei9/bquz5RFc7Hy/83lzgZ
TqtqVcBq+g4l7wP+e7LMyRUUbgQ2gR0L0ZzGVh6VR4uQfeZMVIEsq1iDQLD+HWTs
1404oo0LDs9Agm3phPMc4Gu6A4BLMKdFKRxcp6fzWfgkOY7eCJIUQvRgf3KYFjCD
x7TdOX4l/cczwF1iFt9oNLtpHk8kwO4Yn2WFfHwFCPtFctRgz0RmkoPTjn8xmg8r
Qu6fh9yQEJiHdti9llg4jPdLUJbbmuUanrBZGuex/JFA+2yppgwSx+cFpmX4VV0l
eTADY+jG9fzCVr3DkOkKT8fu4WxpAUg4vnvXKj8fL27xYo3iu83Zts5dC914dANv
4Olh+fzPrwlAmmIACdAaoqeJZ5qibkJRmeJAX9aB5EHYtrOtOf33woto+ZnhoY/a
EjF6eBGH6K5YMB1p/fhzs552ShcVNW6ZjIH5S+WEsYGCo/+crKY6meGDp3ofCDua
If2waawsOu/BIPyDBpzmkqMVAg0C2lEmv0RrbNXfTcvKmijiMGfQ0h+51Ld2I4/x
QvtIl5l20jfVrjxsrFKU14DnmJW3knSXBbR77SKYw1vU0b0+bs/zDSGon2O3jTKn
N/EdTdNekoXilev+JkHQnNxaUU5w42ZFbsJrHW9YYk9KSyEun31CaClmR69NtOJ0
aF71fdWpPwuIfGBR6u+QvAyuCr8RmSAlRmIHTItATKb1/93x3sTJiBsMAOrRffaW
KaXld897yb4GpwxckVn2Vwb4AujA4WJv/fLjLGWD2bYi83gYf+BJP7h8O4ZAwfdf
AXYFDV7bd8iKgLhNrPoVjMvkzitQ9R8grC9x1Uc6ZW0CWkYlGTVy9YcvPm8uL1Vm
GqZFmQARS7uu8ENkD6b8hQ+/QM3hXwNBPjDBSveWypZcKFhXzQ83KA342ksCZ4m4
JyaPydOu2UFKuQ3VEsgIRf1hA2CI/1N7a05rEuX1frKxNZCGwiA9S/YuWTDLX4tF
ectfU8aqJBmALM4084WADopfrfiiAES1GS1CB39mSzU9XdgaV7Q0f+iiMRbkndEL
tINz6vcb/OVACQoXHGYgqa7z7p2PGANJ/M4i6/awXc7z7LjtHMADW3pURwFSRSJW
861mY3leWxR6JZAfM3mg82bwEwAM6yH0LMV+GQnmZ6ZSRu0f09YaDqfL0pmB6uWv
D91SbbA0Cal5f0kiVdPulupxqA8xL3+zMswZCxfgpZd26EIVm78vUoKct0OkoiPi
ENMaCLPWUoNSqbtxeYntQinb4hiV6s9NknEpS14M3+2MO8AwAtlfvFGUW/GeQi/8
tUqGl+j1bgsxxffoZaRJhr226+qOQGuXsmqZTa8nJm3UHY1SfLJ8KkJuIuA4rcve
gis2ncvcNbCOrlZhQQcccOymrss+FHGHw6dQ8snaPBfP0twPoFb/GI8ZACPBSAmW
/WgbB+mdugto/geE5jT7wVm3wMq085iV4Y3DNev+893MM9/lHJJF3S9En8WJ8Yr+
xSZ3IlNp4Sa0Rp8SrTXZ5XKfI9ZCtPxez8RoTIc6XHq0ltV7WdZWapMF43Zs+MHn
AQuK7/Bj6f/sRTYusq/0EbwO7424O+6gXqBBDd4J3q8HDZ6Jm1RjBkWFjOg1BtHm
Fbh3UArE/mIn1SDG3m+MmE8UXPUZRkniz9zXpyZynGvE1aXB7Tpk0AjzIDDMh6as
qBtdQ7gXQnq5V7Or2edA89LgEb2B2Zf0sxBf6N2+jc7mCPBP3lSTJCr0qrfXUXxL
JJVbT3uzMbCaI1i5pxh54EU6MOqaUuzyYXxX2CiC1+/VUglGZy4GdowQzYO4VOob
HcOOzqKLymP/BQR0YK0Qyxz9TROEt6lxvz3hlWztyGa5uqIBAw+idsHGCaINM/Tx
pXqaY32Ip3XNG0E7BFvGB9o/fr6uqhsPTs71/9YRyQi+45sGSkEyY3GZAuW5pG7s
12xYmJM1AagJ8eR9ulVoWAlZ9Lyp+dXdxSYdM8eLqJMuWqfWe2BNUBxvsaG+9JE3
rWuwl+3ASiVS0JSvBaes7/81JqKmtBzuj/HgC2+c97nZzNusas0OY4iWiY6ihF2U
MOha2VFLqMY7IEttdGVle5BCxXwoKtwDz3KI6v3CO51OPXYzoyJT6Ha2IB9IekSD
Zza1MIKlwhuPNWX7bHU5zCqqMuhcfD3xZdxnGAqK7nbTxXtw3BI5CPp0AoN+vnhn
Lei5IgB5LU8lCpRSeGjnVxm+VX5792rIMBJZ9s8QeysxwugS4uy24rMw7fCwUGm4
MMLnVN9O75W3jWNLavGqeRd+vVjePzo+eQwmT0FA1wioKdKCJ1olyTYNnZ3tBiHk
+G6KXZNeLkQQbEE40+u0Iz8ZwiNjwmRCA6NL5knaJbcU30kELOav188SHzhb4vJ0
XfDRUuIkFvG4Tr++ipwj88BRgSICmoieDNsfmCK+2wzKjN1I85fA2SiMCd/0mH15
AA3WVTxsBTDyy8ZZI70q2mSSoWfN8yN6xEK97fVHNiVShOY5LEQyXpHaiD8PF7QW
Pm8MKSmtBfmEeEwsJxgh4HBdiY/CG+cwuArRmdoBxSo34aVioWSSKhFbHiVROqkv
jJxVQF3Z2SKaowFSEaKfetvCv7gWLKfhI7gZmdKoZ02fRENeZP2wHDpT0dFvcdWJ
61GsQZ/OEYX5v4hzGkgAAdXvcYp34mNNVcewI9m/fY1jBvBJhrQHqhp8d+R8InEh
4gnUxHNyls2lpvd61t/YMANa1Bn/KmBEshacWXcOiFJLWVW2hmCq6u6OyxtCr/9V
ICVJp5O8NqQnPyZzZU4J+5D8DIeLyQQ9zadQYzHKDnFTIEF0a2w1odpyE9BtMF8J
3+xViGmMIrKJ2VSIzd27+otx9aP8iN5SBDlpOkhFA4s0jjDN01j+ZSryDAbFNy1f
bgwyj3JSKUxpxXDKPzRCbLx3VdLZWvoHg/ObOq82kkUMEi8x5SQ4hRRSrGfXap/6
vUV3O/2v15iWkfn/mxORJu5dor9dAi31SNE7zISdGahimv/VIGlYfqJ6N4jegFOW
MLHHLCXf14a+JYuLGonF0O/DRrptbwQJWqvFfAUytznv1t5GJ0uf6vYj0DbkpbMT
DgwP2uAf4SULnY9vJZvXSpbArFYqGlnolVBkLQx861UBQuYzi2yVIPhKZaLVJlPg
0F7ayaT1Jb1LhYhdqnmJXUpzBzglCWJX+PrIDftmkbJB2+098S1qx1LP+kj9m42v
dJ/L8n54DYG23R8Nmi/jLaiG8Tu1v71WfVA/VgwzDz/wt2AXsZFHFJ/V9E4x5IRQ
lYNIrNSW55dSILSQ8VZU1g/BXYYGdqvK8tqMKutVj0L0QyAWklB+AnENgjx2SU6l
zK29v+xAbfC/Lx7E3s5RnNwfMWA/9wsmx7wh+Y7s0gcWJXZRaoRfTIF2NheXyuBD
6g3af5tvBUjMaCOUywD941R7EzUnUqoUMwtaiSyLgyM1yl6t8aomRxByonI85E3+
BiYDIQINHwHho7eItz8VKexSMTx2ULFtuqlEog4mvLjvNJCLWor4RI+yGd3bY6Z2
TmkOtxcvpEF6o+QlH+2a8k4FdqQTi5rYTkpV9LwGpnhrQBNCgfvIfYzkHOsKAS3f
ndsD4TFeciWc6W1ZuVrtJ2TF7jMNnjNokW8VbCCX8Xzz+05FWu+mEKRvLIVhSZgl
Nvph5btmAx3Ok64OofLuTM8NHkwdKFh2DEfHo54AjyN7gJx9n2R1hFagBhj3V050
dCrzqlKVoss2KKO2WMCIKU0DgL2J+560R4flkbGeoGlCr1I0BCpm/iJNp6jU24sM
VKXw1zt1lVKK/x8yx0cO+86fLR1B0FzI0JnubSkTr80p8QS1uKDi0fZpvLm0KY0R
3NK+dnJQHe7kbPl3/z/oG1eIubYUvfqL17mm9il6XILsG/2BdKCF2cz0LTwEKbjF
EysD/AdDlQSfzXsgybNCfYIBoBO8lB3lOddvyjkIt5uzCKaNErn8Zb3Dy08G0Xnh
13yjDWPQIQzLiIcdLw9a65CMJwPvkzylMxaAEuYG0HZXvO1a0IEl5V81gPSZ13sc
Jmpu5vCRjLsIUK3BtCIeb2VVEQqZMQ9huoxm/c1H2swlkUVeb0nV/lFvxaxQ4HYa
B8HTM1EuofQE1zVIj1dQt8ocpyuYtjS5JyqWBYC6/bK0bo2biuKvbyU/FQSG3VG6
155p0KprUgYU4uNDnGwdQvh03biT/N282bOJ9ryrldROC4nozCSn9MECYNEapySb
dcnARo+vRLRtU2T74WZSYFvSGvy5LWsDlaFoMaQZXp1ct/EyMY9yBhpeAa26TXuE
FikpN//6uQzcgnsMiDk7ytEFzLbxEW06dJumMu6bHPQRKzc4/YPgJPLn7RMCbuEQ
KZfx5sZv9wq8HlJWEhdLVT9/7CV75WBEUz6kZSj9D8XiyuKWXRxvRRncSY55oirH
WZcD9I9qGYrsPA0sHIDxUSVrZD/uNOwS4sXUvzTGXnfHhnmNRChf+qD9O3iHDSMo
37Dxc9R0I3nYb/pyqz5+3FH75hPUJYpa6VtxrbBKKlEmz5GhyiJS1E0nFG5UqHA/
UoIx9amF+2fQWYgdWbsHptXmU/kyqzzrkH4eY4mlxXMOtCIO6s14RfiikTzFnKpI
o5GNOg6KvhvPh/fqY/jIV2vlfhGBxWVyAX9d+urXRInvDOQ0FGrbRuvI4Nqm+FF6
nwsTBwS/0a45qEw7GBusexK5VH0IhjZRjvvlJSPdz1EHEdy/yvXdX2vKlCSXQCUy
KO5QDp43xrBEJFn+5+xO7aSnO/h4i41efaUDT8BRGgtJIO4nbAD3rhKs30npl8bY
9S982OVfFnf76FwKR0fAMuF8K7GwbXhXMAfZJCIJjy0zVHSW5hpBAMi5mZ/8fWN9
0PSnFdg6TAiTYNmOHz7xeeKYic20fxl91HS43XaMSIzlq5ac/iq/0rIcP2k/trua
zlGTwD/IlzQ0TN+F1x60qbY7al9Sl1Ky41+txlCl4/lgdG3MGO0A8QEfPPWOfgHr
gErts3+LEKc8pwHvBpyOyAF5eFS0ntuKjNwV3v8QmrTT3AwAoSw4sVhq7kcA2dGU
xWKe2kYc6QIPdMw+WEY3PdoGGc3lp85UW/tQ55okf644JOIYExSvSpXF7FRsj+b7
lELhy84Uoo6/q5g4tc2NCCtFRWw5gneWoP6LVlQgyPFUoHrksOlJbYdhABCGEjct
yByMFTSptrvfN3eq0ub40KjvXSOKFrymxjYjqF4E1QD3rhKnHPZ6vAONteJ6u30b
Q01udnbcJW8RjV4Juw8EBuA/EC+9mR/TPgSsyQX9HPGhy98EZQ/AZgKhS4K4A2JT
B3Xjsouv4ymL7OzoXnkpmAj9YOm4dBeKTDwBwZ0oWxztvF6MbUE48pVQNf8xXqzY
W7Mk1sV+XR4fK0waHMSq0lAfUs1WdWE/F9JANCEv1sSQ7Rioa5IYBp+tfo3dZb9/
ZvLmOxe1yBfjVk1YCXJVd22MbPzyvr2vfhCBy4gcxHMYGW8y+kLe6th3iNf66vJC
ofFy1aYMm0ymKkCyHDsQara7PGuB0hfri13EFFoUtLJnaoIM4+PNBmgRynbCguw6
MPnpfFeA3A0rdcgkRM5PzUWwHn6qriRPQph9/suSl9WILqHL/oMjoyJhh0s1VPQi
/dclzyYeOIT7zQJKdlkTTbnDbgpwQCJCoyNcs4uIw2wumWFzI3/ugy6fz1STXuH8
QtNPTE4qV9UQL708X032svgjOqac0nh1IBV+9qeX+RHKYKFnm9MYJzQF/kj8NhkS
dpCs9UivToRAE3/wNbiKxYaPakUg70LAdtVy5wiGNVU9DD0RuiTyIcdnhHgGIQWc
ZJnSVpYBLp6Ur3a/6XtkLduCgvSz/KQCipVsOGwCiPZcd8E6Xv0BYag8qhj8g0aA
i7Ky+fBZgeqnBC5ns+IiaBjJtE6P+O0G6iHKgczZia9S8Q10oUOQ4lmWN7qXrUvk
x36XRwgu5HFZNYJNfd5y94+NePA9tiWV/O7UxGtzitEb69ZGD/R8FUhOP35hmmah
taqzE/QOEINgrr0XrfESqIt/saLg5lDK+P05VkFc2gH2DOCtjnEofZydkNkjnhE1
jhohlgPHhZWosfUUMP0lGTO/jDZ+e+5YzLiCjgcR+xvalwZbY8i+p8CJeM8qx2JK
XJbp8PoeH1JYEt1i0feXR2Yo8gxyEEIuwFZ/WecEHfwYXBknwFwLIK0gjznRFLqU
WAYd69El1xP1dMPTtjLzuhsjUl5STkmbI/HS/cVGr0+cPP5dbBNZ210ZnVWbGC5B
SXAYlafaL8pk9Lw6T8S/Q58vnpNYIqxlhuTHjHa7Oi2YUbwCyCfXHrmbH4vUzLsz
h5eGSUTirWQMNB8iCHpUE9syJjkoNr9lT2AMwz9HROIy1hwbHMC6S0/7NS/Pw0GS
RvPfZd6TPK6YViTbN+enKw3vfVxI71FKJJZNyx2qgQkPyAvMw51junZF0GMrtOGd
KVpxjDjNdPNaDL38GtXZB0shaGkKzuGzRJmFcQqU00fcpZYegPNdhOn4MV5ivs4e
sFPfmugYqL9KlwaEcKJfKWkyu2GqraTP1mTHrIfIw+E4S4xAGKSkW45F8HhaUuyh
B1kwFEi6TcC3YmobSIX9n1wQUgWDpdAi2qq8Ktj1MU27XyXDDbQXplRaVfqic/9b
CrQIOJpueR2wjcQHeLak+lW0NK3phRmkqKWIpbFrdUeWIrx1OJxv9/bWXPpWfQM+
u4BB8GDlbvJUhlKrcmkGkoyI0R7LrZT4NOkOKAPl+zVLzboD0RMDNTnKlY3TZrJR
2oa8VUVWEO05uGxuaChC0P+ui76QXtTz83+ml8ewp42pM0zvv4TD6/uk4Cd7btTk
6rzHTfHHfQl0VG3BjGULDpp43cbDpcmXO/B3zlxkTGlk9i1EJpKPHIkgkQtPvPUg
8AKpgp+a16Hzcxg9gnFZ30KS2GNR+Ds/vo/NGWlTzXriayor6okc7FqdiewJBlXg
stiJ9ybBae8WPfv16TlU2qAPAzdmzfSY/RMEqC5MR6GOCAmN7vR0VAoqWuWugjkl
0iCVG4M42K9QRwxM8fxN2YECojiMJq5aTLei1Mjk6Ja8/07UJxgXipE6KgdeTjFI
21FEnY1Anihsq3DjSelSWBt6UuEGOEJYbpt6Z+6o305qIZ0PV76+xse2FiQo4MNR
2t+CjvjObEUPokPemi5o3c3Qd+oQ1UN7S0AfeQnJTnDXWgaGxRD2pLnHt1AUG6nE
nzoZyTkTsRij97svm3yk21XERkh5PRq+6tzVwl9E8g4RunSi8tp36jXo7xioujjW
jlfZgRlsnxbuLKrUCg1pgJ2uGFYo24CLtuPCltIjaQlNEHvC+N3HzelXASSYUKuz
/VW4rH2go+DQV6NEMc30TEV9ZIxfeE9goRn/f62MA57rTRL+GoebrUpzt8haQ3pK
dt3jRTi0N/w+rx+sB9CUjGyPZRnmhjLcBWOdYp155qP54CNVhyl+I/RkuMK3eEkt
LIRgrAMWtNK8HTPXwdllcN4DEII9bCS4Oc9cxUCldl52I9VW7VMWTzCNjKuDiKwC
JSekg7Z3vq98guVUaNq4IH1+n2GcE7sKwqGw7Hf8qcfanpo9jfUxpL2a9HmYyBB4
LwLwYBrDNIkJhqPCUc7BmkZ1YDh/pxbajh64y3zmtmBb0kbmJ4ZWNCepylcagaWp
8OAYncKAkeqvBJe7H/LjwYjRjdsAOXS0o74esQJcAgKn5Ewa5keLlbZkINhQMate
GO1pyvTyXx94L7OshWvgPb2mCZHcGPil4HO1ntk/lBRES/YYYFmE2Tea9YZAEHgo
X08i7lWoReKUio8gj4eO/n6pXrzSWFQHm25yC7jpwvbx2Lf3aAQCOofJ/Rq69jZF
c1obL1HE5L3Sk5Jp1ERsedUvuP6UKi50wwUma/UYZ5LOfKemcOoxL4R3TnZzS0Va
NqrXaLw/yt8hgjsDQ/RfW5xKX+mT/0FnL4jaLNZoyrmEH/1eS3laZK5E+KaI+F7/
dbpG7m7/f3YjeOd67CMPpqd03IEVTXETdi+vX78zqQVakIwxngBw8qfTyWOklekL
vDUsBa1V/n7GZQ0UMhRiZ2m41yL6nkW6BB/tKwVKACr8b0pbhdJA+njcBG0WlW69
9YEbD6HVWMG1TFD9GeMXfhzPp29TMQapT1TOEapMqao0ScJLU2fmB7eVLKLM74mr
wW6MBeWSorcf8w3chMDQPehaMMh2tirXpd7hqXSGKkGEn/OHygky3kWo6p7SaLVm
40uPHDuDBdNHWwxiHjgbE6wbKfaTn/Ts0okiTAS9tY0zBWKlz/fs13BkD/X2RK6t
VAnFv4X7qt6PlIvIjYVi77sPZzHgKH/5su9Xuuu9O6E+KvtwOvIWCXgTAL2v+z8i
dmeMM46B6jX5+TJzC9Gf56oHYC7pJzaK7oKvv3xm7vm5wX4rrRE5pDjZX9p0dWmj
nfEOguX24zUKMEvUDH7QXZ4dpkJW/GIcdDnHan9HEPp4Xhm6SgpmSRXkjd2cuSqD
GQCJdHJScoTB00KTpHSLOPWyTrCi9YP2v6Rs2rHpiRiXpsIvZhTXGqZPaLyuWSor
cZbBl92W7MN8PuBPSiOoX2B6j/cEfU9x3Hw1mi4ImOdE9ndbecSciSDQCH5Kml9Q
Z/KnGxW5OZpn5o7mXzIF/IKkcfLQQGNE5gM4E5qfJwqnlUksIlawKseLVJzGGNsT
34KOHBCp51nzHsL0GIygHDRxjqZZqJ0s4Mqhfem5W+Cp8JDB7a0iEITPRkibEBR9
E3GAemSJZ5nH9tv+/ultbvP6KF61fflwmGugcoLufBZS5PfQdG+HD9JV/qvhqiIL
yy1zcMIp7Ablihb4gG1nd/X59NaWND1SyOfG1RNhe/K4U0uCEN3RQdCDBG6sWPNM
ZomRSaZVRPC1Y7lSMbSgISVU/QiYXdFpLXQ4SoiH8nj7lTmleFBfPkpW2JjdCfxH
Lr2680bPv3ojXyOF8UV85rDGH0JgpmmwHl4tHO7R0CrdoiObLqkEwGiS/ULawzds
kHF+oaL9heeiH768yFaZA+1Zj4o99KaJw0kBtHe3U0m2JGpDIjZZUTjmcFjjMCBv
OqsSRRIzvftVhuS/vlMLdg0Kra7NbB5CesDum6cquwR/KYqqMoGMGoUZ1WJCqw7E
CXyP4mZNCfzh9chtsU7bIcKgwr0oaeyPHpy9kXtvvUBXoXcqec5pBr7GG8rx09se
rVAxKo0MKkrvpH3SN6UrQYjJREz2U1sWGq8+Mbc7NpzQfxZXQgTml6JrsG21Ee+J
PdBB/BWpcuUTOOOWmdfM/UuG6K52M2ZWlxlVMxMiAcsarIvIhQjaeN61jEfrzgzN
gSyT0i6ZPHDi1vaknQTEOfjtFoJRvk8XojeK82XeT9SJHxQNXTcHKaUMc5oHmyaK
0hCNlHSZ0aoLz8ZkG92u+26u8J4+ntkX7DZlQgRO4z89BA9Xq2ee+SJgA64wNYtF
1HrDZRXI+1uFSeXwdvZ2IMD1JGaOQCsmSOs+AbsFp7XxBhZcAueXWFj/9kQJIbUh
mdG3mS+4pMXG/HNeuEkcGt85FVlCnUZgU08yDgrOxdj+xCP0QUgZZ8hM6bu3IL6J
6hXik3YBaW7l5Rk++pmf+4llbaKkJyGPgpMv4jz8RS6ct+fOrJ/t2o/c3YDXzABJ
4Zs1SQIe2JPyi7M4ce/uxG2JYfj0WEgBOYcWAW4ZUpx27TC7u59pmY5dFFd/SqQd
SDdSdJ2oi9sgAwrVZY4q+IEO8EPr/OYMb2DjGWfci3qZvT6MGRiI3mvq+5lWaYBj
3qq1GsyrIUUBoKw6vO2Om39DQzRLz0BFvODCxfjdzqFQc73KBE7EXJeyD2qBFxZ6
PfivUr7EDkZ6QVV3C00OEUZ0ItF0q/zoBzzuvCeqD8gsoZ5QDo1zhuUII+0kHIo4
yvWcHgt2lraiVw+iMmezmcJO+WgCf5HcZSZUpPKrZ57Y9TYODhNHktFlSoBUlkky
udIiCa27WBO+RIofZOxpNVhPWqj0lvuNAn7Y9YqZeB1JCS5Vt6kxMQ3RtpFKgFfj
vaZ2kIvYEqJwCLAg99c25+rqaIfItdN7JNnSI2SSEsEftnn1+KGe6fxGMWwWA1jp
b/9ip+ih5/oDNKnGdQKo+H6nd6NnMRq1M3uEAFbIDJVA8m5kp/wIEti+HDfsiXC/
9vsQ2rDdNJKs/tL7UC/PFUF7vaUFjbgzaf7gjlWJO2RdpqrfEboOQwU2tZZ0EC9g
DjDpcYNeH0aFnrd/kt3E6gjfS83nj9qda8VaRFS0Day81Rv4OMQboVCjmC8puOxi
nD+k5u75dbmo73cxWEl/v0FJYhC8YvXgY2mggKrz5sqxAj960eEDpC1vIPGXYQR2
aSEfjREQLxSa/8WlBMWi5T54i0HUDudubdz0a3Nng/OfghAnbdf3I9cbum09w+Mw
3FRt0Tn34a9iASJikPKEN09b8//pUV0BXIGyQKUrzh6tLwcrz6cT3SXmI5/MkUCM
RIxHyBdO650NVLZU7EWbl1i5lGI3irHYRzYT+9QW981L/4naJdfDCiqXPSPKF2e5
ARhlOpxP6LrZ2HYBabq0pYtklfZniExBmumtvTy0yE4sXmpCpVtaGLMcLKURwzlx
d/mj0N+uXh1TDJARXpkfxLO2FGDqsdyD4LaN5ppRra87mHVtW8n834W9a5QUuUuv
Rsn9YDaYYTRTMV4UQV2nNGCUIWMFsmDA5796ofz5ekPek4CF1IT4Hj1zavuquBWb
uU1WhOkg2oqF89L+pr94epwK1FL94+XvAENkQ8PdeXRLiCTiFyLxYNYTos4ictDJ
DcHydnYvdcdB+gGa44/LFr7Mj+Jpen+CaEeo8OKuJRv+zTvjBZIOvkh8UiKe8BNl
QXYNvXFULNaupsMTxwUM2mG86Gw3nZTiBBwnyIFiSCvnMfoGDqhteIuyV3FyDuyY
IiDLwG0MihcScR2XxUDQDyhLrjWCun5x/XOf+g+kgp+yBp3M9ZCu3kzDjNgfxqUL
BfGNiM54CGGc/E3OBrFzr/5czA9Nvef8CvKgrDekh6cb/leFw4Jds4GwnU/C4pN3
U0lsCVaTLMtVUoFmwe7KSLh/P0cLhh4KDc9/pDgEUcbtmAFY5veLqJHjrgMYE3Te
wkqnIEnc+JQ5DFypPAN++j8aoUL76O5wWqojrtnm/NMj8U7v8DqpT+mvmh0OcRC0
ml9I/58uKtjiMZw51MsO1hFF/2f5OhQO8FLUWqjy3yZz0UBJP3y+tkA5CO2ZCyIA
dgLpLV7+SRkjJA0YowwTdUVquGBYxjnkGQXO1gH9hdaQnUUDowPyi/EMq5pq104h
zBEkXukHG2tUMRxLaWtr0R6J1vKxeTvzjtrMGtOSXLZcUFIMEJ7h7DxEQHGwmu/M
m5KtqGD4oj8NSZNXVQx4IRqjwn/tilCQ7o9JBif9p+YGCXGJkhFwk8LjHU6uyj+j
ZuVmRBQFBDKYTtRNKZbICOa8Bm6bGQEjl9GQUhWWLEGw6/KEHlfJJt+RS3faJbn0
6pHe7ds454XjMsEBNm/lD77hfjR7wzo7Ab4Rw4NzgmqrgDIgjvcySjFgoLv70BOY
MFG7z+XV0y/R6J8P4ASiHjtM1JuwVVFexktWqshMLfAv+6QFdN6nyChZDdKMrbgk
gP5lpsFY/UsFHVB8LXzeDzRKzybVGe3lse4m2X4hd25x9/wmm5vxODaldGPTWl5z
M4nYttDFRC06tfbnAzkwiouAtebvLg0yzoQNDysV0A8Fio9XDUSNw06+wF+8s+Fj
eIsvKGBSkaO9ID6Y8F3mcgzCMV/RcMs9hDrcoytays+OEDuExno40sCAqss/X87S
nRLeHBov7vMo0QjUfdg8Z3Mh8or0dAK+KYT5O7qFOlyqO3pFWWybHe4erh2BJy+R
/jAfMoJ8ezBpHngbAK9LotNSEyvFrjOskIWVBfLjLkpZfMlahh85wIoAX8fkoacz
uTwdSQXFTX/TlEiUc4oYaIT9FCTJMGc4iz5J8twO7kaRucIwoIIq+pth8CdSLAwy
pHt4WmbvscYEDqCi5qrr+Uufe6TDT6Kgg1ySbkStv1isaH0OpC0toTs7KEL2ZROf
Ilj+GmRxw5d9YpEBh9YomfdEJiaZnThqId1dJepFGFFGsFMHA7WouGMVG923zpBM
ngqfDCvBP9fiiimWpQfV37zbFn5Fo8TPxbGbfTccp64hqY8GSjqc0LK2hORHQP4w
MdV4JTIzfRnhbkDbjCOBqKwF0ovJ3PnkwZfg3HSnVfvoLEFiqwvGW57v/LdUY65c
YwhW4H75ND7fV89PmrNaFHnf4Iq+q4iJtHAJ9un1f9auHI6iN1VqErV68UF4p1jW
avyyKuVUooYvaZheaNV/PJMQ/7LSp7St0UAv5keiycqjid1Hh+CXsU7P8GqLlJER
/fAs2lltHjKD5VqucumhGjwL6GzF2AG3ys0Tqn+nciti6aFFXIeQferloxjb3UJY
tvOWGd9E6NRiY7oQHIpa8Mfp6CDDt3Rma3bKVyfkTZ/iuUd3XRZ75VTHHrh7+Dd+
vK1LD2GCguV9lLQlomifMGRP4OhNFEe3h3CT2aJhLU8y6pjsT1TsJCQ8FqTg8QI/
Hkc4gYXgugTf2b0hjvAG4aolE2vkaFmTi+eeIFb2C6n5JxhPMve70xHU1y70cSDs
YRHhilS9YuyXffH0CaqelDS4WU7CFJpfxMOUy3vkKwu4ksQWkTCPzX94SQDPrvGj
CFLUhjG7wWLn6pmyL8XSd6EeJFDewSLqC7npQA3RKZdX91btyV66Sl0yvK9rgONc
jEmucRL8S/IDPEjgbFfZUHlSreeR8I7nRqGvnAl+FuTWLA5UKulYhI86iCcHS+dW
HlZikYO/qdy5dN4bRDpxiPUyuX7MRpJsUlGoe8G57bN+YaDoEC1ucdXo4neUgUNO
vRWfXNYYkbei9KeMWJP+xYTZJxVzdPK/bynKM9IbAiqbmB47AuberGpIfodx/UV2
bkNQiHvY5gk2JbNO/OhLGzNNBECU2X95lcAPuDMPAF9e4ynSmdZRiFIVQ7PeyF6t
3CC41c9h6+3B4UO/RHvrAXb99rJNYt2CTNbVFUlowEDt+Ckm0CFW5Hbo61O1cksj
3sIaPQxeOoLkrvChXYi6qsdvOyZlR/bUiIEJnj7N1svVq862wa3wI+nY7lX9RORM
ei9uO7P1VyExoGdVIOAwJeYqFdVS1dutX68nLwJfRqAI1NYtOM0YEYEwFvxVwfCh
OXfOGnK2I/XzHs3HjBdaIR3WFAfxy8IGeBkWKR743U1McFwiCosUG5C6Juw2DrwI
HhZ/eu+Io1cN6+BcQWVDbcAVd6nScn3vwK9lxk11v2oqVWfuts0N+VQnj/Oa7e7Y
TiuvRwX1VPsUfZSBjGbHxR58y9gn6603cDkOEenAQ6hRw66lN/rkJxhGUe+h37Xm
DmBjibYW/YkQjJPpTeUmDwEIJ0taH1pEkZLGBmdYzQ47VyvIjkwaPYjUOMs6OjVT
YdV+vKAYYXcFEUgwAtkrZoU2o39J+I2gtlF2SMsKeJeifa+oHJuudZNMHwkteh9d
T/woMDLjA0yaTQLoHnzHo/7e1IfcMmreb2W/AIfNOH8wFiNNOJvhS9aQp0bwa3My
XIDqNtoByKNizVOOLpSIJOwP43xfryMYsmJfjb3r/o0rzzKf9x+xoGdSaUwQMxTG
xoq9me5pJPc6HGlDYyf1gBaR/a5OkOHvPwcfhfHwaCHrgXGJtqIQFIEQUkUH3wK/
T9LHbrFubTkHx49rsELkPzkonPbjhyOVwW7oe5RIj1k+Gmb8PjryFA3fUavpQ+ZG
HLJ/oZ5qpG3cY0gPMjiFl3ZF/kqqmXn1gSHBOxGZoI8OYLy9WgBTIcwzWxgzLC3Y
Y/NIeWqKERRG5vyigU7sBq1uEkl2c3g6HLRv5oPn7IQHt1WSqEJ5f9s89eI73OhN
GOYtNHJGgt7OYaD0EF4vSpKZf2Z+NlySh6SkftPXHcg1UIWG9kYoZcUnIPntcFOY
LJNh9oVf7Cy+sqs6UZhOrH6mWx+BWo4JPG8o5jf6xhroMK9P/u5wpG0qRqalXxd7
ja2/zHGA4kSRNSrGmBH3VwZHnK0RpBDii4riZYj5ICI9xwltn6tqwwVC9zXMY//A
XeB4DrhccjCs6KosJe67+NEIGp/33UWeba4Uq5n4aIV4BY/u008YmSY7lGXHlb51
mjfeNXCrB5U2KpD2NJ+sZHRX1ZkUk3/wuIGAdREqVb56sZgVJGihRb+1Gk9OMWW/
AZVBC5cJkiW4XuTTvzs75TwM3G8tJIw6cSWpUFhVEBnffKrS5YOBd+Cr/TLctZZa
ine27/esWR4uxcaGVAtfaNdww2DhdrfdsMLt3sJwxckwKJy7e6wJ6xmviEPqiHv+
epKG1LYal3BruXfkkxDq7dHsvfLSO6ONI5TTmgj02hPHSQJhMQGZGF6lzPAcAcRN
Rb+5Z+36xIbOiVgIyAwDo/bRXXfUbI8F36hjgwEI7NKQZXv89y6rUQ2P0EaV3OKS
0sRF/32Yz7wPVXAiQsw8mL9z1agEFQiW4PwIWa/nLOBEUEFI8Deju1oNCQZ7HELX
ihWb6UWRy2gqqLM+rG+vk9fptobFC4fqznpRE5GzdV352Zofpltno88/fmo5w31I
u+7pgPzswqY/OlnXp+TBr61eycRG3/2eDH3dkXSEk+JlMKwsCZnSoSHJpECjWncm
Qfmf/rl80q6Lu4oIFon9CBC5uioyr0b+1h0DKw6WeOdjt6v62WbAPtXNvJDNFUQc
ZtBxXH7VhQf7admB+zrIY7s/iyH68zgNPYN9TOByZr7I9omdkjE39c/45N77KmqF
EYjrHwGBt34cZZiAqMhMYQXoPHZ9DhV5MuDIA67P85seaG+X1Fp8rGydOMaO5Eli
UXYrcVt87LqE1rTvNErGc8ez21aCbgEdwrjDCaXNXqkRpreUxnAUH0aiLIIZyvJr
ToKUeITPgD9UssV4GCeH61fnFYPT84FhBMuJc0O17cP0xoB3En6libuJl7c6JbXQ
rczyRULSKDj+AiSPu2YRqVuJS7Uw3m6vebPErxTfrd2cUPwEs+2F4J8RTYIMUS4B
jQAoMDyeVTus+J8t3X9ueR72yp6W2hkT7Tk5SbBfCbNvISxY9J05yqMQJaMIfA3C
EyOGTboPdqu/xnTOny2Nfe48YGlH222kqKHWtKARzeiKlCigQCnRkN9xZ1U870UV
GMaJJkwlV27LNnBubDDTFbgQya6T75SME8fOc+rzBK5Jm1lqflEyz6HoykGtXfZi
+h3xDgWU7xtBVRDsEGjZdm6FOBRpv32CVdvhMV8luBQvfzgJ3NtupRvQG/KmYQ5n
Q6TUMYmMF8aDzLYxBzh7NkdIaM/B21FGw3QwmvbOIAmggDrBDd6OLtMG+FfEXwwl
DtSGoyTv2fEW+GkQAGXNRqWWeRGXT+tu6POyco3TTvDKXRL6GM0UCmeoSsehb5Vv
jQJskqQDX7e1igf10m+yRP7qBUH6TJhY3Y6Y718v/u6/3Q2YrOik7ODHURjuPcaw
xDl+6MjS0R+6xBo9+q0QCrC5WiLfqpWiFNdprqL/MvRytb7rl8IT44cJuSFea1fs
HX8qWXWDI9Sc5guigaXENCWIq2NRcClDIzQC/RK+vpArGu2lplkKse3GJMBDLqBh
7/i7RUDq0XFA8UvP+Bx83eFCIV44YsQMoe6pL6kxsU04+97SV2gdFNCjd7vE6+zJ
qkbTQQqrkC/jd/1V2FpgD/u7G2aQFZTTc3vpjdAzQiae/rTGMqKKzZoG1yJzugtE
2/bcanleHvSITkN/44fe0PlO8nyYTButSXSJJqxl1f3YrA1Ed98b2D0T+H4rcFBU
Ol2alAtnG5zBVTIgWAgpfFy7MhjgRI7qBvHAoXTbJS+nZLTIWza/wC4cbXKeecgu
9BSmCQWqkPg0kHSiXqB2TAXugkT78x7CY0LGWPEQgLCYvs71onap/EfBV8lzweID
UNNXxAaqIiwgLankE7hG6MbA3I4ILWXnbYYE4AbTJ99OR0xBFyYRHEu/DTsnTp41
HKmpI0gjeDemFjRUrL6BrvsiM+iaKNBvg05lP3pJ5NftOJEASST6zczVHH7gCMw1
mIstFKRfih5YhNOdfezvlgIdZg46dcwbNzsEtl8d/KrRn7Oxl6tZPKaZNPVkD9Jv
Fvihzjrii6Lid9EJjrdzhvy3ox0/8E24wE433t3UJfJnjcQC3QU8Gj04lkcQWmDe
kOq07+ERF3eLupEM/Shw5Gxzgla5ajGFTpn8OIbeaEycTwoJfj5xdlplRVfh/u5B
uF73lqffvrvctC1stsvswocvXYSnYubWe580y9MInb/9x7J92JXO83wg2uOb6ipy
FO0eoHfskYBWsjHFoXMxMmkRx8h+c4Yqgi8yVAL5QH8HXxECaZzPAad7DAiGWXOY
dYOo5x7+lfXJIUiSJypvT33TcZKtlzQXRsWwShWV8vMmv+K7IVIrJeGPu/vR8KiN
luJp3r8bUJH+FlutH9ldVqboKLPaFipBrW1n26y1eJ1miEpKUQ12PdP4lhXJ070O
XhWtoauBA0PrNRjxvL86M+oR9/sd9Ly670HJYT56PGG+s4xhzEkGPnYhX9VuGYew
hsj4DGciX/tbMvIxPAHGHrLgYPUEAEfgF/K5NB15zmF3/RtOjLWq4icyWVJDUotB
9IBROu4V8DHRjZtiMMdVZHca5mQxxSkvjz2YgTTbL5fGKrPasiikr9fRUNr5qjj2
7Nfsn3caSUTdx+xeC/IXPb9vXcHeNpTSAh5ywyT5379eBPdUXs5Qp3wO37Zwhv4V
7tdFZItv4RMso2qg15hi1HXUz91I4Rgt8jTPP4gBgmjjW9rn7EaubGRuztVbgf3Z
JdfF2JC9DZh0RyN3WN3Tp8/OqCjnD7amBCJDYJZXby/YC6OnCpijNtHBzDXF5ISg
OYmh4KQ/KDs8OKVRjz4WMgjVj60kIs00riHRCVkWl2T7UbY+QaJUebaFWD1kX45F
OIMieF9U0ICh7DOgmFoQZA0iJFdHA0H1Lwxu9obJjk9xrD05xaFBjbdwOI+nyazW
xbuGtsG1fDaDi2XJbTSAVAtHPzTPq2voNWC+9xxOVvvDrE6pBDVgmm2AJuGBpTas
Cspo1q/3MgB/TWBLOBnilQPnKMOzUrCGHFZ93vLZBDzHPzJkZOj7ZlsQksNmkrex
3eImjbAGKHglDerwxeLZ9Hd+zWLGl+jUQx1zNJftKWWPXepXj0WXfq2Pf/lsFYUS
HkbHvuo0Bot9DcmxdSQ2Be5BmtHWvVRVupcFN+/UDgqZcYojCJMm0CQeMKlXyKmq
YOIPbWfk/reONVikwb8hbfGl3KjBKEyOET9RGOXgTfFoqp/TBedb2jn4vyF5LbfV
R8zor35Q/jnNYlw2KkXlNyrqo+LNwrnBCJv4YkoMegDxL+3QiMFNZpG+VZlwIuoh
emAOSV8yNJp27jrJFMsylPFx/EalCeneevcuKjZN0DkxeqsTrCdplPPjprLlEDfz
wO6R28FRw+bF118vOZBhJQ3I4zoRVsOeYUx7dKHKYYMUHuDmX5VAjLNYpPj1kmxQ
4U4owY2wajVbN8IHDzmWv3JE8IhOjd4B0DSlq3UHR/mXmsfHqDhWDjcWiX1s8Ad+
kKk1xRPnvIUg0YEIRsvq8Kac42K3e4rTY8Xsd5iGbFPkBym61l35eSfnuwMS/cYZ
Sfjlh9Jk30Ar7uTiDK/aouoJm/LkJGcVfmKVTgWNO5AbdcMZTH2SJXY+lzQoeiXZ
JPRokW2McFJoPhYEiPCNgwgvvuprPZLmqOfBtYMeKZy6I0MszS4uG3UEShRJ66YX
w6+g8EOAxap86GL0LTFibwAyHoFGirFEwA8OJlwfZAAnfblirfHRdKWN1UcGRBmI
tLx0/rtU0M1r1VxNv00+h+QoTPrgtHF4nsXsfUPslRHjLMbIofh8kPFYApRAvtpZ
aQk631qau0DWnqNbb2OqVrxjzSekcXr300iyk8xd0ETbF03raBvMyI0sMbbacoM+
otribwSnI6AleAjx/ri4TsFh9+EYyMpB2agpje1nhH7Fe5X6pma6frjV22i056kB
JCxguQMynyheZMcSri9AJVR6No1WK8O2RakWMe5bRdpRAiQ9g75DsqF7J2x87vBm
LegYaIJtW5l2JIxoYE3xWgFKZbZyZr22zEcKxJHwpNbeoKkqlD7xInm5F9VXklHU
7s7GnV/HJaTE3Dct1SHf1gYNwOtIrj4nlomtdoRPSzob96Z5OUpsV8mgEV+4NTKC
Njd0me3AbgFUNiOx5jj9bg6tplYrIfosmCNeKW6tZmHRWzshEejRSsU9YXqzCSaX
Qjdgxo/JO/tQmyfQ+DXDWrWWjS4ft/518s41S7FmeBLporOFu4ZrrB55JowM2UwS
+aU+p9VIUD08eILMDEB1qnKN52fKIznumvhht/uz9C7vI2Lg86BWHRcy7J7G1BnF
XyOptjFGvu+0Z5JBe3I87tP33u5do2ffQOdyfOkE89NwWI9FPSgXGxUheZe6BbeV
skRusfp33wRmi+0GPnr4jjfwvVQxrpSoDZJ8oriff0QIsHT2dlDzC5hgLVQPSnTz
4ARazicZyQ0qkQQ6GlT1DjsZcviMtP6H5BkaPiyqnTdOqsZ2MLZ6j14OGg1630aH
EAwTZWPOjdOLoGpjiSm2uMmrarl8tcPN2OWTI0HOP6PCD6xsUyKQzYr8fdTw9Kt6
+zhA8hNFnGGHsDIvkPs90KQ/y0vmCvIah3C69noea0ecyxBfk3h3AwNcae4IzO7m
7qg6CtIdQ6ioysQgaWlykfKWChFfwXWYGugIrjZ1rYPatgQxqlZL92drGLRlwbPo
CnH7luP2Fs5ixVjAcmcM7/vrggE970wXrYMeRFb2BLltVccR9zQ/Y22FX3J5XyGt
YaiKAJ7ngLuAFFimCH3LJu5rKhcv4ewz1vOePEgUsXAPhWnPcfM1aDxtOkD/aDhR
i3+cbESqSLF1Yfj5YTqjYBMwKuCO2FaS44OxqoQwscD+SYDTx/eEgx2N8yzsHnjj
+gUMgbh6jjPmJKmKSW2apK0wXZ2N++wh2isjRPzh9ti14hg32FdgeMN3+/2A6h8y
bhzufCAIpEXyIBgio6SsyCgrklErO56ap+NwwT+VeiJIp502RHb6BfwR+YsUggXc
74gn7TpHwzIMtX5rvejO4ZqQhCzdd49Ta4kc1zdfsOkg7aWLCU7Phs2e+E4XvI6O
ej7TFCW5kh1LHnHemRbAWtnsiIHwTNFck69d+h2IYp6m5ASd8GnuwzX54tYUd/Qm
BO1rd00+fxyAgFEkRa3dQOFgFNEQk+7+Hh91ZocNsCPYCuaJbIWCgEiVZJyBeEc6
wQqda/ao2rpve5m+EcE8DJIkWd8s7+EkEXkxYnGUeoy4+cSy02EYc3hVgImbre4u
R6WOb4VI1oflIRfCvTXzhQrpvK9x64EmHQrobBvDElGtR1BjBZrZ+9bEjtkYV72o
4wvlNEV8WCDXxO9HFI3Es9ZpuwHqj3mITZ1fBbB60esyrdNp5W0nQaw13eQbgzAZ
YXiH06sto5Eev2ToqFZbt2dXhjqB3lVN0FxfZyKDusES8eqaE0qJBBVZKB+Gqtn/
+UelAkR3b/BCPT/hLjBZPLlaTOIhclHSrClPtTNQlRKXUZN8BbaIZi+8EofQVXWf
XxB8ZucOypgIU+gBEBIZ6jdSLqHxyRUZdzDIPROm1nvfCmdykwa4hB3POYibd+cm
AwxzpKnG/0LezuBmMonAjH4EP8MOghJ5MR86Ag312hmWbgrtWktv207FgVbcXjzi
uXyFkhLYn60CPx1ND9hOv7eJr6iUh8EsZkfTIAIsLs6NZ5jInrhYL3FxF+AEFWE+
q8Np1V88uS2uXkyMDolg27XsE9VoDr3PySp9LXa3yQO0uCVWo6bnYXPszDpUaR6F
XW9xFsIu7kFiKRBpvamt0XTEpYr77EnpKO7n9qn1N6cu5JpJZdJuHrbjuEIKKkhD
Hgkc5IFVs0nI8QXTavW+VV+BKplPz74g2KwwoWP3BEVZrxXCX23kYB4n8jzCENL4
1UGgu03hNJ8A4HWY+shh/VPrHZN3iKTTwDpc/SbJeF8zxcacwEU8OZYvcDCNPn4Z
MJOHKUbiskPvYkxmMM0SYXFdsUGO8aYKpDv3M35sf9K0LeKojisdlI2eHhfdn4n3
+AZfCIBYAlpvm4AB/jl7Eds5TRbBrd1+YqJ7O1/PUk174tok7KGr7ecCs2DgeO9R
ySrD2X7XiQ4gTHOUiduA4S7p3KZpxW7UctwMbXEU8vjeVsNsyNaKKiYm5js3pRc/
prPdeANh5HnLDCwCGq96c8PL6K5Twmf0c2zNgcJSUWSd7q1GcmqTC8Vye7xDp30W
dEX7WgrZMbMCWlXEC2OjjQzT2xjAQ+/VRYbIvIg3qzTZR2FGSM7wC3jmYIOIvzix
WorNk1nbYTBCRyaGorTV0Ht8IGC+UqlDOyJWPgVY57tSlY+Efs3LnT/XRd7puY3q
xSAT7Iqv4fYwBO10Ug/H05iklNKkpUqp/i/WlGf4omEmrUM8+GAV3niky0qYTNnG
ayMXxq+rqUn0fNdCN0N5wv7wZMw7C7UGb8zp8/HWuYItxyMN9mXmCunwcHmIkDof
VbDYFZQxuemFc3CTKYEhsP00nhAww4aprAlgWRU7ycymz6LcMzjMYb5BQZbifgA1
tbDzTaD3UtWiZb0rWdj//TLftyufqID0VMPDw8/v86r21KeGuMS5v15x6ZX74yZS
EukmaMkiqWrPrt2LoWRUp/pqZTxzkfvXXPzB/1v+Baun1iGQ0mmcWn+TpnIp80sB
0O7/smOx0R1o1va8EbDCzRlPc8uW3zTWYOvKfA6Oi7O+CX/9ITz6hTt6DwQQx7gk
+1XxxDayFDfzcE3+uY6bPMzFEKPPbTXklQ0lvX1FFtk09qOCbLoUiyaodYiHWfqF
aYOyIbAj9wkasqM2MDDlVdwjcbehdpII6xTJpIDeA2/6ymYWcNgjk81yFbaAlGac
Qn+Lz4idaJFEqfEnc5KHh2qFysyoNXlTOCmUgIAIJ0gRNR3Iv57cUG2jIlajdSoj
SvuCYxEHjVIe7iQGdKmDTvZLCIQSNnY8wtmT24DVyT6BoyVePEKVU0Z5aWn/iG/e
mgHcVxiEXsBQ/YgiyFbPdbOlsBsByufOF/U7P1YVdU6/JagSc2zoaBjIue8cLtS2
U6IcK5NebMHGct7gyTQtLmOdawwSRFP7ECatV8U4PPOGTdtRzalJkbG5eOSMSw0U
W5/vCTefi2b5PuVjxhOSjWKF1IGwJnk1qLgZc+l2tFVSJ0mzj9rknKIysxj6qxr/
U+EnnOijsGsqiLlZodAr/AYdaukBpLXfPDooOWtnA5tzVhBai4+lYy9FQQ9P07a6
lwzbHYvVynHnP4yLhd8OyeIiCrHQ/2Pjl1he0phpPOhxJnJMvVgZyquNnDBuuUhi
KmSLxRj5KZ7TiWetpPZDawJKTsTU48d8LpeBeJ3bns2stdM1UFuQLyFnXcxO7bXj
5g/aoqWWj0n1SJ2QFHGdisDuADUCv9WsmYaquoiaiCZihsnibqpYhg0ZCUpUvNph
zLuM4wk2G5gKNqTsI3cA4Cf3Z2Ve4fUkpQv/JfAdOelHBjd5T+CcRVXJfnNDjCKb
irTK2AIRM10mLJeqGyYhUAHVRjzhJa+G/UXrEXD0AISX1E2lNmaF81o2cj1TS+NP
PidWLoYpkF7Ta1Fy5O4UkPUEdYuBs86DvdEUcEitaN9Rd5dR14zM72czGZygLgqZ
3LVYEtYhaU6yQ9YZC5jwxcoylCkVP4JUUkRyHltZHhFfm6r2lG2bf4xNV+LG3L+d
oahTWoNHjwIFD4SsKklW4JQiBX0OaasqTkDMN5wygCYOxGKDinR6ZS3p2ZVA17QF
5sUBlmGTyjRMe1Z4ALlLniGmrttsghclWf15eyFIsOC6dNTcr2jIN7IZ6s/9FRL9
4DSkBzwF/cmU9qc36aMgUAhWcSaCngIp0/6u7ZdIR3oUjLpAUthq1gaPdb+jriOX
eDgyxz9O1aKxbeoa/YXgOJgaK0rXxxpVb2xjsuNqIPs1GO85EGZi4UoqrZes+FR9
+TPg+uxJY8b1k2KipD9YrPYZAoRqg3pyt48Q5QDhITfVrxdqdnOvejmxlwxrIcis
BaTFgnjZnLBx2kEPeUxXkJv7r0IlBEshcQsxbB4UbVTMMidCBtw6QcgYrrm00VEC
rgbZB16UvI749CKvgDKc/d0W3wmyG6r/W8B2Hnx+bcZ2buRdZDkufBf/WZmdeaJt
Kt4Yh6+p3G0Hhrk3XNaeReVLaTM4uASlmHk/W3yTzOBPmhJ/7Qa90UsmfUO7Fqqi
WEdnaalJP8qSR8TYDaKbLBsVFlNTy42xahMUns6/zJWh3k3XxN0I7ftkT+2BPLsn
89TIqJJ/dOeLtao0WaV5GgHsw/BuU02n0cqC0x5iWYv1rsLl8qlDFwavlrtAQIsR
ndRvN3ounanyBqEghZvh9yNSkMYWwOWlasrjTmNhKmsAvA1fO8FwT9XRof5Xdv/L
FQhliDJ64fgSetLvuFGRV/KmQ2dewf0vZR1e6VGMBUXZq8c9N7sEIxs4AJvnpIYz
oFXWPBIo1dSxpoTBSHVLh8XVYPKNRGfOeA3m8+LGgNmjCs1vXd/T6iTQJXLOoh+u
r3g+3jSVH5byzWq2izMlMn9Bltq8v/SPHb0TjJcXv8T0TkwdL50GQ5OFHrc3KQXr
0w+2aYIWU2ZkrMvlxJIuFsTH4IERlDIMrzC0GiBaNYYwvUBgHYiGq2qSrMTwZooZ
YPzJXyoKv3oR42aUuwPb9Cbdn+nm+YG23i4WxgkLb6Vi7jpGRcbHb7Z5pW/vFPv8
y4eTj4ktrC/dB8PYL5n8TY+t7dblNMMaMZx6KFd8xwtVmr6FmSCSEbRu3nDr4KqI
GeJoUEoNOHQiZYZXm9qcOGVryfGD4L/fAKH0ia55NidwDWNJOAgsDRUIcfjIzYsl
1k7cPVcdijJXdLMMwh27PKXw/sX4OFucXPav36lNTn/4t11VRXxPfjiW+IxNacxS
njKW1TE1C+OMVGJS/sQ1vKrtiMzEPHPxn1978b9gAP4RywIA7nD33vo+n+LaGov9
o7W7sodvMd/GVXr34HOo3tpWn/VV37c/PCozfZrsWO6sWubDwz9JoGx9lxCidVmr
xdCj7Etbhle/9uEeYI0a4Wz8VWoTaIkpoifBD0WUg+eXsElj8Hza1M/2BFi4zAHA
6seGLSvph0k3PMoAe2AhPZxoLcw62h0nbL0vZ5KO6pB7d50Kfbe2AcdqajSegqiW
YiCniNADlfM80sUdl2XLexsHiaUheIdQ6x1H7Sim8FCQGA2BXr4JRyzCG7UfVUnx
hQu7uGXy6sp8S28IkNpNyhb57P9ZZECgNKtYFTFJ1dnkayQGd3UZHB/6mD9riw8q
BffMyWTKyhBWUb1uta+CxDnH6qiE43QpTCwef3eBsfFSxU0f9BgRYQI2ynUD3PVN
7R7ymNIQsp7B+4ABPgO8VLx16WLJl3cpLZ4D9gm/VqmWKolze7UFm5jSHQzWIGiF
XUh7YqoCIGAtlcOopTyQQd66j5gvyaD1us+uOGvU3uy+/LCqXNkGI7+ymFBCG04S
iRPRvbHUh8AiwTbyZdbevuXsqJhA9DU32ErGdWTjZP2jTXPJdCTaIgUX7hYZGwEW
Ej4MnFrpqFIcd+HmZqQ5K+fQO+X140B4UQMzJoVLiJ0Y/jGU9QmUhRXZS4N10eBo
zHWj622ielAnSSOOCz6MyQyRd6dyshApf0JlZs4CwO0Sx1NkpoKpAGHp10LoCWP0
PW9EY0u+ajXmmLFNw1+5kYXUbCQ4/DKE57UBP9n7Zh8NlNRf/QHFAx/fZKQKooIM
8Ya7mRuHCKg7I6qrVe8mc/I75MdsdXH3ecbu+plAmWKEKejAhJ4iyR1t9Po60Bqb
4tE7Helzl8jDidX+uNG1V2CvUBJHvsCRrnui83UdZccCO7C4KnSMXU70rTu+Hf7J
ud6qDrtIbtWJ8mGqYMJaoUDYhXVSbFDLq2suPpfW161o0t9lbTL4rqzDZQyCNe+z
AbPsRfApHA5uR8xipUzGr9AwPfldOp4VtjGcXRWwy8ZS8dLZib1ZeNDvx6F1cRdg
KcOV27CFfbr6azajlSc5J127eKzPSTID5ZhlAOaZJSUCVUTEo1KW7XQYsIWx+eN2
zMw8gtI3GGms0R6wmkKcnnkZF1E79XG9mbiwiCsnwYBS2lKp3wYZwhHV4JYHDOho
5CLAbjPPIX3HAqZhdO0ZJMfimobCip6XNtylrnQhqIg=
`pragma protect end_protected
