// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:25 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kGj7ChELPRTwhEJRRZLRo5nfscsa/I0wMTsx1kaZwk/QrH0NADmob/qcfGm2NHoi
1kYlRffR/BamClsy+zD7ysCUJt76NyVL0aszlVflMYfDt5SErPKtxWu2Bqp4w61a
68ChHfVGm+vyZTfbMHssrT03OGhWnZLvQS5kpa+3w14=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
3XVkSTnX4kXxlyQcfC5VkWsYU0lf5YNCUnBCBUmQZPgIuk8pgA9bixLy03O6GynH
GXAVVEqY5G1DBd6S0I/8Ui1Ffn28VlzEokMU63F93yMtdNazOFQ88iWh31LhegkV
dMYOgSKoVCXM7fTJQMkqnPF1tjMU5faiiKa4OyMxuldSsKKuWnMHsSodNgummhZS
R6Iye+O9qW2h6gvAogq2DRJAiMuYYOxA5O5owxh+lrEnFe3R2JJYVwVOzHC1KezW
vQIBNUUkdYylC6yRbhLAn6Oc1Qqw5No5dGO7lSJg0bD6e+Ak7SNN9ve9kNoEUJwU
BlmmGyY4kjVWc0rhRH6gEPVzJuHFW08lW0ad74wiLydltzxrKUzu0PvKyj7M7nIh
3/Ys4uqwo5l41qJHWwb3uJ3itVgfSn++vriFquqF+phbNjXRnFiWbIsX2sUZEDIa
SVhu45129l+T0VQckay9er/3eM0zmKSDd2E9O5mOTnC7qtMBWN5Urr83s8YdHvfX
NzWe3BD6xS5JelESC7vHEHZIDBT1tf+1NOyuQGMbLYQKbpG3gaFve+TypjrME73z
Kb4pGdcYG20hKuuC05En0jY+HKoG8um/VBaHSRQSt2Qhw0q7Txx7xtwpqJdYaIqk
4m0HROFMYYnSHNkELa+FZ7NL/iq+9xP3Kzh5GQxngtzp7I+jEJyU07ieRll9LKiy
2kFnSWNDLVrWyliIbCbrSUP4aReFNParn/NePAdBMkeM0+klSJ6bN8V39cN5iRrz
6hRu/ZRkPA6HheS+vTqc9JJiAUEfvAeR4SjeUS3c4PZXMpI77ksXQZmVplH8ZBaR
KfvIw3C85KurFT+YG20GkwmUeuGFqtkWunspXRhPdOKoIqsS4NKMZIN36JTeK2Aw
Rr4vMLBo7kdzRiWdU+trvTwslt6Az9EJCqOP/jAOhcJ3UEy+M37JOGeZySzRoQYS
7TpSSOHOc2t9V5t0qMnSdYruHvRwe6Jz8DjYCMGSrrYjNbdqDHnGV4QWr3CglF9a
b8yTugRpPNFJnl0qMyxNZiM7KhN2vMfObUoyYzsfxq27O4vPDWEo/9e2EPolL+MO
TS/F1/ygi14gHXQXDnE943l25XL3MuaU13tLeVypDIb1vf4gZJhQu8bGEw+IXhFw
zE19+CQqIPxjQutqCIY8+VFYOtlyNrFUGcRqhD+IZm9EOE/ai0onFg9IePY4pzjQ
UQBIegRvS4mIBKc2NV5fyEgg1DgAiEEoCYoSsNNEiuDynXVrANIbpU2MeC+91wzg
sW5fjyve5XZSbXg1tUn43Wsg6uameJf3eZSRXURuKKukoBwV6Ww0zGYwvxT1KiBE
h6/ki7RMT4IC3ig9thGNONTVmRIfKuSzy0Ad3sa0RDYZupoO1Rfqs0IczZtg7Ri8
Oz2XXZOWaq4Lg/deeG3c2uCWDHLT1wqItafCg2ZHFPjkMWVdpVtFqbkamnL1UB9v
OkSsBcqKZ5Gklg+p/6xKHepztAjDYIrgoVhkQcmAT9lonLN6DWICzN3LSEht3cFH
udRvU/5lWIFHorlS1krR+pegpQILFgL3as5rHGTha3LU7l2ou4RP+hOkk/jvbu1S
pqZx0/XeiUhZtODgWlL8MOZQ/ouYksjTJ7C3hOVl/4KjuidDJztVtAfo21UukDCI
VagKyA70kF0CaBnT1/DClqHetlwMRyjadxwfMFCHxNFDmqKwDbmsXlSm8ODq6wNm
vJcbie6AgPsBQ3a0d3hc4d/hq6RVZLd9EOaXCeaCFqu4h2bSzhcsANDaU/t0iF48
7j4ejzw9Xou2SoPk1fl5ZTKWHbnc0d33UxZzJXVWC7XuqEaRK8glJthp7LjznAST
qO5dsmbP2LBv33ZEYFxajmG6ylO3FNX9mpVvUTXCLGNyXntd8a5nmCISvVulEzFW
03azYyojxTAdjdgbv16Wmq1v1Y6ZgdgqXa+LuG9RQDJt7WnSnfaKaWEGDUHuIaTl
Y9BiQEmJCb+5vKm+p3QN35xDMYmE7FRMgml3k9wAHp6PnGMDFBo/1CwWZAf96uTS
MzSqVF1Nqm8cvjiq46/OCdNRLhOfqtY/FFSJ8F9/4ZAIIsTFgakTUDPQ1KmEKRke
lx808UsMkIkqRVXfxUvCDL3NbzdVy4f+3FWLrxRdMfA+9saKHD46csjbW9OyVy9p
LeJ2I9nOfqbSuKIQRJwYpQNUIf1Z106DgcK6+mMefq1BXkXTbSKPwYvmtFbS6WA9
wUP8XKKAdzXOujYy4JKOIUL0/FNsIxKF81OvcNNJIjMdaDHJbhQMh8bzpw14qpjG
diGr1fWoGpetCqvQevqdS5QbxumsmkoFsKDEyhzpHcFXAIwO9vLseNA+hFOjJR/e
YHvVyJcqc0E8D/mw3ql6BdR7v72feIUqoumGZHouUrzjNyeNOIzWYZzAIAda6hFQ
p4RVpXEYyi4hZewb/PWZEHLrgu6cBCr9sj1WxO1h1V8aZeDuT3IQwtL1CMGLFkWN
xGxt9jO8yIkEjWKN9AjE7FvGtYMOLUi4Gp0Djo5ueZvwItdgkxUuzcbq/aw08a+u
Z+3O2iS49RX46Gtui4h69DOSmpL4mn9zb/fQaqP3g7Xo/Q6Vmz4ui/D/yKaQWyMJ
s8cIK3m1shahvaUaYGJiaFGdc65Fzx4aSnAp5Iw+MldjmF4W9fBgKI7kbofMBcb1
+nwnzsexZ9Ypwh2AbqNhUcvWCSH0o0y83OzqB+mBUNCvz1Rs6khvkY0c4sUjPWa2
qzP0h0oGxR3RTSezX+kXimYXSkpcD080Eob0STIhmk7t85+ygGb6RZljgl+5zTKC
Ha5ysGXcmT6/gDrhSJi6c8OtF1xMwJrHcXKtz5FHYu57d1flaxuWRADM9SWI3Nov
ssltzxszcqEE7yFE8jcTUQEhnYXxEQstRE9qMhdSeRWh96s52gWDqamaKdAGq3HD
/v1izs1bTG+EQ8YNMe1ScQ8O4VbJxWghNCX7jtb980X1gjHSOl/te3ZJO3fdbhKL
aoxZCZM9cOLUD5YckWhFIThjxuvnIpRQAXsND+1ICPV8IRx+mb7pTEcdvZ8+BPrG
LR4iNQbhed2L9qq0OU8xfQN3zeyRegutdrqU22H0BlM/rCCZWPGwESnD+1+OZ7Iz
r2O2F/7/jhPv/pJ+JMM1Bs1ANZdVuBcyvvb6UtEPm1thNX4sx/8JB0QkjSoxxszK
Q0Pw8nRpBxVJMNPbbIExO7HqoGAx/sVwx5Ib+/U73EeKXN3DvJ0E6aAVcAinQ4m1
gSBXmmpIpBRqtoB6Uegv1ASUV+4chV5t8m/UHUC+r87wJrKsN6bHqOd/8Ygvk/3B
DQPpVznUFTnaB6XxNgmP9/vq0lpi+mFmR4K0nHr8URZvso37uH0lSPAyVJbq4IMz
VgcDdzVrgPID8TzGW81CR+sjUIo0dsSdfN/VbJD3mvmTQlcBxKofC4X7YP7+zSHX
F2pySE+eNlQhtx/cihDcbPmUmUESKTp3DeTkLAtjIapsQdmDg5DF+uuTFCF+ptTL
UzLiVcMtB97B99NNIaYp0iI6eiJ7jhEthvxNqbJXkro8slV36W6bYib/6DBrMWf5
dBTwz04p2DF8lkTdxxMMn7c0ps5HGJDLYrchBW7ZgjH7Mwk1Hl6gRp60+qEztaxv
jEArD5LwB7SpNFGirLsAjAOJJoPzTXU2YLMyNSr6ybAFpLsvXWM50UHxKFKiYpw0
HRCu4M91/jvTgrFoAJf+EZaEJ71Bc0WLTFDL5DjTY39OE5BSZBFNq72UGWGni8lO
28vZZgfHzS7fgHtV1EZ1fczFc0PHuBMsOfNs+vQAkvYOwddjgIQ+TwZDL0HQsR0o
/yIL/o7EmU0q0omXfbvh2GPQLxOy0Eke0j6Z3BSc9nzqoccqIlUQmK5e014EfI3s
HfRuSRbDkEhNCfh04pDsvpgfzEbmd7P97VbLxvnS9GYAG2aoD7oER1m0lhFqUyiR
IjZUklKxJPnWaROxgz1Z5xEDN59VIWaZ8AYHiHvwpV2ICtVyKniZ/Jnmh1/i0iz9
9UDnq7QJiG1WVw7VLeG8YBdlUpzSwH8SqUkTtOy+IK0IaDRvxCK6bTsWhPD6ppmd
E/ghyXQyuKjBgT1CPUEub5dzsNhgl6xy5ANVReu8ILHyqtNcjJn47QbPy/0QVp52
OyHHJeJcRhPDJW2XP6KnFV/XBKpTzO0DxqBN4okNCwZIzwp0CvDhoWRbiIUoFLvT
TnEQGLFRyyaUOcIrbGxJRvcnlALZ51ZahGYt1QsDB4auSouM3jmD6Giq6BDJgfCB
6H0UWM3Y/duq2nZMY4LihuawcCESH+N/f+eQ8yWV8JNpW7OYBVcjsB3FLXMW/HmQ
xzar/xPtvuixmoz7dJ1ZKULoX267ctDcvXokWrij1DUlq85Cy9ZhWOXmJxX6BF6q
TpmPellhoaRcEJzfsMWOv8RBy4Ma5H8YBc8IskZOUGSsHbc8+gW4CP2KQSq913uO
EcHUb/pIJI3CAhBIez7ho/GRoZXEun6b5n3xGbueR11wR3/xBCk6daiL2rT8ictN
bDbaiST8mRLaQf+IL8CaILfbkxmbBxRGDqI4rwLuWPKC2MilVWoMSNK8KFelMoKj
r4wTG+0B7lF2+NiY9VC2T7MKAZ6/MOyFr4dpR+WSJ2OA5FvUjFrTLXKbQF5nL29X
XCmMZQeX/reSSTjSY0XN/NcjQFhnWob8N39Zbpc0ESVFWegQiDGOlZxrArBz+Mgu
l8oasJ7BOMGAxpWP7tNZx2AUXw/ooNWX021CAgm+KYUaWwSDEWmdcqdzjVm46tLK
2J4vJXhMYKp+wr7+BjRQl0VDiknOHHhN6TOGTkyJJp2ZEyR7hnmw1nzkNPGle0yz
OtU+VDQWtjR3y/HqRdJkGEzMTgGlnggR6NWkmslPLHk5neinMd8M9M3srQkuZ+XB
f/TvreM/cTIRuxxEwZPk+437xOb4EMfqFPUqDnKzfH8Uq7sQMiqwa3QORbSWqQNV
Y17KISmQ/WMl+6mROKLZbLxpH/gfLkAekpgZdCZ9QT3ERj6rX13cWSpAWcr+rKgN
8Irf17Tq72gmmXXfBo2GZSdM0AAHtJbt83u3M5KagsbF+zKI9BJBuFNiF2kP6agJ
5iF7XukqdR11ijLFEO05j59CAn4FuFMWHDL86hvk71Frb87RnbNuGYgiPK0keDLD
0NtswjusKvpbWEi7ExNbxN3Gd5rFzjPm8bA8gQeYi89eCmpWd51SLDz6bAlOA45H
MqkHzg5Ov+S8PkD2kCJDQNmRIm6lC27GHtWsPlsSXddQ9Zu+Mi4V1xmz/vSJFsfQ
evDiu6AC4q7jCnRFO6wj+4C+ea5zNQSYG527G/ReD1QttEjMCNc1jUukfTfidbKa
72zFG2zkcx7OCwDP55l7bG8gYbPOun3kn54D8b/1iBTc33w6pYn07z+lf6jUwVh+
5bZNILBQUHrItvvetNUaVzYmXfY9WWkb+ihp51jNSd9An5vMPzhbF3RdgpVZzUgz
8a/cLqZVIAZHXdUYbkMoa/scqD2gYPUuzMWTviuIl9uS8C8j5yCuYQf/UAds92QN
ZhpmHSfK0hu+xj8ZwhKptXecAUC98RU7qiQpghR5iGXWbj6U+E2oYho0qDskwPi7
94GvIcxpBsPDVaF5pwEtvtjKXb/+/pIj6Ui6WIVT9dkx8meNSUsocfUxqbtVIQov
cLEg8DEOORtYCt0ojDdtKYZ/BZdpC+TN56rMYC/yjstVxxw6AuY4je20QfAX4JTA
/+z9fbFylTtA2aidv9KQtclkVQMF/eac8uPRRDgIihsPA6bc+oIjAHG3Pwph51SL
fLiTL5ivH5llEI8/UH19OTpsGvLTAcCFoPMXgwfCPgDeR4sSLAlbnmHqTsF90oWP
xE0bE9k5c9lGpEjLhfDwYd2N5cLlcIXLbp01bUaZmNLWp//2mLxjTMAwv03rAOwl
TL2B43AMdoF63pAmaHPouWRnJyhkr7jCjFVhmGZXz0xSp5tsZFMOMHNLcOrWdLvm
PPrVSato/nXCwHLb9n/bxLWivMwpR2cWHC8ou+bWI4pnP4/hfidrx6ymmVHNYxcP
t9W4hUvQcZ6mMtFYMsjutgpja7HsA8nPTfSphs0itVUPTzXbQ94mVitQJRV58aVk
rnAPjyEsPFJCqmVa9bY2yIt6F8V53rHHdx8H1O29n19zJDsyMFmw7Hoa6AHerHNF
sKdqOi8HQeNeXg3Lp2DMnq0dYZ8o74d5pxCTj3gkvzhdfleyiCWJPIOFMbwiKAXs
CkUN5bdfF7Nx0dNaIpI48icCeYTI0pvtqptovNDn2rhNLFEegouF9r1zkZx5Z9bf
3QN3N3nlATuZUwl6aTxMclROod7QXIKFzl19oxbyv5kKWMBMhaohx4UiNy+a+4la
aDvzkjxldgWOtkIV+nC1txL1165ZaWjD6Zq9G+sMljm4gpZ16Rv2taCNYWj3E34y
MkqebhX4m/7m0FiqJob9k3uZgLcw1UQrRK/dDw3Gk+pEdQugXXW+fIqdsbm31FrX
XgXlnkfjt62SfAtGZq0fDzIonh0tJly7LYvVCvbZCFW+G9v8iCjOQPthSMG7Gy0Y
hZjnEAMZv+WU7CqjBe7uMn8J9XpuB9xRjBe43fncwmDr19uTG3tJPUfuBggzclNv
8+eFiiOR1rqCWTf51oSTnuEEYF8k1K8oeU59IlKtbh5TM8vb+Peea5t5pKrMt+yd
5ymWZeW8hS2ToCtoiagpYaUqmwnzr7lxNcm0Ln+zXz/zyA3pQgUTHcq2fkoYiwfg
S+iR6LaDmV0fPs+HTbs59VPWJ63OxeCmOEHXO3Xnz7B+oko5dbMqQv9b8tYhiCio
+mdWuhxt2ZE8VkYnAnAVO2DoYIMfWEUprOoaxrko36HVVy1XO0R9CGAXsqyct++w
SM+3JXbdjnlLD4C/R+VECSzScwVH9sNJF92r0ntGXBGIXif/ul9Kh26v15dZAsda
OGJvKKr9y5tZjNEXoPfYyBqyu0mj63Z9fBBpUm+Jmx0dcxQ5AYuGMOz09x4iVeUP
CokeKCSvhBUd89hdNDiTit0v/kkqw6K3HY6HME1r6WDKAHNfCNd0sdk1xoBL9FRe
p8FspZpDocPXmyd9dkeK0asbwViCrwtnN84JZ+XNCpXiy1hhvcgu24fKcaBHYy0r
HywrAmmHpTw7WYu6x0m8Y8/joG/Ul+GJLmWsBhGZQepbhbnP1SHO+yOvdhKEMvx6
x6ojh3c6CsDtGui1VDSKtt4hGHosEVFrHKSi/c73vHJaVorrwdGbn1iP4y/tGA+w
8KPo31cgeDtAhWdAQZgrlhEUz9MqfgBT/OIHOL4NgBRbZpfEVtkKhLBizn9lIeuY
iQTwVvKeE4d9+XNrZvXukwZelbq+/+OLrq7B6UoBVb9wdq9LAnS5OjRrC02R7kpO
81jH0sE8RIwCnzKNk9AIrzDgWwVyypdT15PTPrczfNYLR3nWYusRAtnylE5ElP40
M4lfRG4gA8wRNDdGTDzsPRhy16c7d+4i/f3DjrvPekcbtxlWVXq9i1Uq9GPDOn8x
zQnGDFQalIa8zm1d9rNEQAeKxas3XMgfOAwAXFQlGdGxGXSZ3JamrKNhoUPBXZbI
r1qNh+QIwz4t9Y1iWqv7nodhosUrXlrc699OANVnwqubjGhudQCZEO1QPDW44WFj
vNo55C9sO8IWJQbsSbqR4ivb1qy1cprfNT8qY9r2wZo=
`pragma protect end_protected
