// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jFLFUSdOTcAd3shsEhykUwuL480gQ2DGui3/Ow5PHWL6NCULjO0TLb6SwAghtSIY
WqGQt57G9E37t4A+HD1svOaR2bQtR+gGv+bLRHhxDRfaS0Q2bBXXBRbLGSRWEiWp
oOcMsKCxKjSJJX5TAEQ4jt9tRCZsNdh9Fxo11RP21sc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7728)
QwUX31+pMPXsZvKjZgR7ew07Bep7KghUH+bnQFkM02ZB6MNC7/WI0quEX6GeSrEP
oaAAF86sMqrC3Yu3l40tsrNJrIhEiwj1DJIb96+r3AL5Jkl3G5Qtlu1xNZJ6Xzlw
G1efu2a/CFi4AZO0SllrCe9XiBuBca/DGQrFOQ+mDNyR/c5OKRHxsSQwinLXFExV
kIbgBKSP1eLQF6nrfhSi7wYikZ0grq/zLnvjTtealhdmHvsXR8CwSBhpT6MSi1Ry
4IK8AoFX0DuhSv65IKHcvr8LrZ0LzrZ6AjmiKfWqFm3BO36tJ2FlKjCz5CupAmvM
P2GMOPYUrkUvMjzMvTcuV7W1JILoOZlY0U/VtTbo/tIhbCAjmetdACcoCFasLE0b
VgK9Wvh5/Nt40sVj/gIw66Kg8vM6NnUJhiLPhzAZxUMS4oBdE7c1oCG5WmRdv0FW
tEERQAIHvk8XfCd3wSBN1uVx4OuA8G0MF0Tth2AU23yXOPfMZJaxWD0esNf08DGu
DDyNZwDDCFvcK4NNC1hmW1ZPEZjxSIkGfpvDf3zfzT18SdhTx4WPfRjQyOz3lGRM
l2/+RE5UKcb334ZRBCZOs4ozdQEgdKyzz9QgopghTWUak+1HlANdry5D1rbbKxed
s4XHxFDlG/wOOQY6/8QWzEQcsMMGCtPCzVC+9IsaS5WEOV3hQI879hToehNvdV2T
WASQr15/xfVB0fAe1mZrZfkmrHN4fciV0at4bg+fm3p+SKlEehkzCbdl8VX5qD3i
0khm3Fekuv1AY4A6hwY55y1jF+zi0tDIlI2kFG0YAiDq9T+ZcpZhNxxPmoWQbSzd
8H8SgvKkzsSM3F/kNz3fKnKWfSk3Go34eXMbp9bfwwGW9CSxcbgZQ694+GPYFuUn
xaZ1BHC/W1HeTQOmoh1gJF2aN/p0vWytQWTw1m5QifvVBiKMkGhKCGGvBzRk8UbL
SNbfwfLaF+GwaNQpdQAAlD1AJWm7TBSC8sVqCPupYsJayLv+fpjOCIZDS9+fsS5R
WigUicmMPzd8dYbyuYznAKkltk1pBeyZEqZYETvyN3S7mlXY/hGaM3HcLS0NoLFA
SKGDkrqlafRsTkO/Bs3R0bwegUhGHO0GQr7foTVBG2jdCqaHIRkYBLXZfaqFvFut
PbiTS5TaxgfQFudfqL0nWlzmgmsJqMkvz42XZufyJdRzmXJ4rjN3CzbHWS2T7y/G
n3+2RUYctCmSO//x7/wNyRMRV8JPdxsUShLPS2DBflEOKZyCL1mFLc+wVUkunuTJ
IG1wIbzZ0OiqHsOo4Oeq2ZOr8YbOmhnFbKGbLaRV3osIeavo75QNLU/7sHXnqLYQ
p7qNO6cvQ2v1eLTvB2MqTfP6XsYAOC4SM8M0MVz9DXuvO5vuhHTMQz1WJR4KRQv1
uJl/qx67nVtzVb4VJZkWijl2aJ7QhzMTkpVsw9a4LNVxZx654a9O2ohWmN3zYe5z
ZU4R31bc8TWVuz6MAj8HqrHkJcLxsMMdSMaODczu0iftMItndHF2ytHD/wtyyoPW
UOYksuhXp3G3Aoa1QjJcTXgIDFC11/Uhf3l4kIjWfaz1ESKHu87ph6LNqXXb8qG9
VM+1kZfb1JSJojJFpVCw1jjNqV0+Te8fkOhDPJzhQaMPTz5jj1vGo/1BomdKg1AA
BLYXePICuPK/BNNEnbDYipbCIhV23yTAzBwR5DrwUVO6HO9yQ8NqADrBIta4ivbl
oj8yKaJ4XLOuPsWdSoDDg4zqIyvIZS+GpNDAyycHHTFkSBx+hAxSQrId1n2tQXu4
UsxuK4TvK/eX7w9EtyIWPFZG+z+YrtBsBGRLIh+AmaxJN/0aFOjN0iUB3ftqwRmn
VBP6i7d1uis+lPn6KYbzaKt7ZGsFa8hzB2k43Rm+WYOSp05jPZpQo4I2Udx7sEjZ
52HDngqo37GUo5ceFOVRwLBk53O24Gn9RydNuszKhWBpv5vo1nUH375t+hBM3gNt
jnaYX+RKjW/w/LLNdcHrYdufAFyBkHYMOEkJpWziYlxPG7tNX+VvJAan2P3oFJ/T
VEHviz/sTR2+AbQ/eALmNEjJfyaBgzHZG4fP+jY3nT1jXbtLhLF41TJ1jcq/ZE3e
zPqqSrVbtJbOLLSzwx2mWUspg/WMsfVm0mGc6wUfIxXeefd579op4GUlCOpsfcwj
8HhUrJeUy5wDZE9QmcKE7mWt5KfOwg25ivzW0jOg8/JGDLrfylAwU0tq9vWT3IRz
bGT3Djes5j+AdShIlhqBj+7c4MCL8/P5nAT1T4CedwvWJSzuVHe+dA6tJwRfDwWD
dYcCaxMPuHpZ3dhaaH4Mw9pB73qdXcRrcCpz2kifIgwEqwy6kNRDV1bo8mUiAfDb
GFNh6pQxMBc5AANWnlTeKaWKf1bJkVA/tJu4mjN8ul8cWENTCWM8nxXX+TkBR4mc
bDoXealdOGQr8oIoCMJCyHqG6fe2p+8y/wynd384r1i1uT2ducwt+449JIfvJrB/
PkbQS/oBMfkvGBI2yhZ8px7yVO+vAb+mgAH+9yj1tvb89zeIDZgxZKISsUD1ZFUX
NScTE1fv2Xq7NckasMhFMiVWxErkiEeTmax2tkTV16jVQM1ds/ZKIBdfucFuRtmG
0m4hEP/W1s5GHq9QKcTXGFErz9+1blHR0oU+v5vrSXvWH7xTl/0JKtJeZu9HPiVN
wp9fzRroZEpkf19YThFn+Zoaj4KqY6l+ZNw5Ow7V5kbsti4emgGpKWkV37tPMC0J
czNd0WfgCSzyVr3BeEIjAVx/VLdhIPQW+b7lJ663zmPOikIq38ix/pd2W+Lagi+t
KO5+27a+ceuWyBhGq/rmy27bkjZPha49XLsvuxEf0DGhMZDD5SeSvSKMTvtvll0I
SNPW2fLIfQwCMJcts45dX09bLedIlPqULPszPeGU/L8FeppqqYP0ECNmIWQC+Md4
Z9UvQD8r7UwI8ATcBTqDiZA2SdIvAK5arsw3cp97RjzEyY25Rp1JzrcIx2LMPmlI
6v3kOiuscyeEvjfVBbQii8OjZxC+aD7A2aWAo2RP30rcPV8un6gtp5ry4MVhx0yI
Dp61VHJY3Z4nckA1mI+dTLgukdKGWCua15gQOTCmle6Lk+ApLEAwjeraSGJ62y9Y
RMtmzj/oe/X8aXu0+s3K7KhyRPCPSogPGu4U0IkiIrr0Ylj+gedlmSV/Oh47odRR
vGyNB+BCug6oOtnCA1i7Q5DieSTtpA0XuB9jiBxRJG8jD+r7YblmSCgBMpZS++vv
CDqTzjOhSBgzcVyGZj4/tURoBMChDnKGT1OuIti4ifYxHuV6RB9NkbDVILxLuF/H
7Wru2hMyeEp/n7VCxNqcBOFjgDdb/RKQaqOsJ0REPvOrsoEqxLYFYGfeZQ5l8cmW
2S4NzTASwoO1cI3GnHPszUX9xCQ9py/enzu1Vb83P61JL81PcFsMJVZBVZgg1xtg
uKEPCZSRYFACUycI3218JO4hUsdP6A0XgQNUana8tYNqLZSKqDXSai8UscvBXJzQ
1XxeSQitbHlPDblUr0gAFForLwwXqJ3cadOKDoqIy/lwDyx2y+SX86k+NfsbKUwo
hdjAJaE72o4B7QFh3bDtw/NC+TJRX4EAWiEyxX08OYWxTCDShTsR/p8HNkcUJ7i5
3CBPDsVgq1XhHmVXx//tdWTVp0lfA0r+ND7H+KWILmPpBntVrN28+Rpy+EgeD2IV
vJc+t8n8PRWquXD/NA9RbWBdyOnbVsghidU1TXqreuBBWzLqoiFVpdLHKPaThy+u
gxJYhHq7MBAbFpfFHfnUUTEnnVv5DvkPBDA2xnD7+80K4DbR+cePIVDQA4TqQFr2
VUm7Yx6P8y3LEUfzG9cMH/sZEttirsVL3r0FH4doJhacpBBlgXjTObHM2OSiehgC
S4Yz04Yfl2RfQGf6r/Th7hIb9gbBnpauUi8784mIiGrjkFT16kmZNh3TpBmNc1TV
DfQn07pQKIWBgA/J2nHcE+KbD92RRwVzOXHxIDrSbk6lM938RIgHf7tQnjLYWkoi
CF4DfcxlVQg+GhOz8pqdz3MOt+sgFedHO3FmRUR0ArEjNBzuWp1qhzHMSG2crD/T
g9efht2EPYjx97RvYwe6hSPC5UNoyDayQdeVWTpD4DRGbDAMk0iAw3qgSCmkZ/WO
Us8LSJhq1MjaK2fCupchKNmgkv5mFhvvONR5YDMV2qcgQmbtzXrqvm9y0FDnlLSy
D7ZXUTWVirC09RErNwAoUsxVpFrHk9U3lN/F7hoNVO89/EitYf9Ie2q1/JUPKwUa
OdkqZXUYXL8XLRuogzl68+LqKRdjQsrlwkyOBvTRGGccR62e2+j+izGQSVONL/wK
Wl6sWIj/r1IfxRj8irswl7yj0xAIO2bJPsyNbT2wTxkmWQctRh9cxZdV6iTz8qud
45tkxGl1GQAgaOJekNZqv42kBZJKBB92DSKhb9YBQH9GgKhaMUEbRKo2uNemLjlB
xB+fPyFow/ZMX5IUtfLKV/xu8EZM815J+iSBqUQ9TV7wEeTPzrdGPgPPZszYAM56
8A5rmoNzHcKDpGu5BYyJWFQzn/Y4cT4bWfiQ6WTlsWMnT/btgjMugm1waQ+YFB7/
j/HjFwtYKeQVMv+FKwkxn/XlfAr8IHDiZowZF0mnUQvETp8ss623AoX6ZCIfQWKJ
jzldbBou6pfrmMH3DtbeWfjxO5aRLe8cx68K78K1GTZgMis3KvvNGEtnEfv/u+f9
JkuWiAEc0p9Rr/tDWfQjGyAI19wtaeoSsHDT0xhm8DbhtcRbDSMfv1vlBgxJwP+o
kKPsq65M8ELiATt+Cx8UWpexQPGM1BZjEy4+Y00m9lQ3Ji5FLS1FANWkj3lonSTT
lP9wFb74tQvM2SGj7vDnkRruwqgz5POzMoNINMGVpWdIvgfRufL7vlGx8e/RVajK
99amRAU/vpGrE+vxZpsH005MMSU2dJIqAGfyt/bLVzHFbpYLscb2eKGX2llzTJrj
zdFkk/bLXhQCVKwCCTLs03q7IurfTRpH/qSPJUfno3u97sLPUXEkzRCYTQWktXGW
oq2GAUFqyIXn1i/PhLS+fAUIwEMI/+cZpEBFP+dSlY9Cv6vDgTmMKTvj5xqbOX9f
Qndog6LxZIq/CPrF9buva7tZ+I3g0fhSexYPBItKiPLiwYRryTKH8+f66rDecZL2
IXZLeZl9XCB/ALYWLpTBpRUNi3t8KKEFcFIlI4Ca5szUVF10yUjB/B+jFOoM/c/4
yDJJThpfNcl64jG4KBW2qwvSM1DE6WB4qigkHowkbqimYYZGLXGiGa46crwKspvY
em+8l7IODyhIzFg6KRcMgUL9rPDAc+GcTDn/DT+bcl+47UYGHkiFp27gTpCSAaT2
vGhPp1QVbub0ZOxhFwZHZq6aQ1PEfkwTESL2aXDAGT9DE4zmI5FZuKXq20QYsihP
MHl0VgBrNZIRfC//sb71ethLwRaJOoV4GfT2cOFmoyIcHH5cQyJe1sos3FKIedvR
48OMzA68vF0aJaXTUA+Hu0+o92Q9c7G2mILp3YeQpvjFpXS4Kn7ro9QPnRvqvGjr
s8iWq+ukWTc9BHdWO0JYPV/xBDzy1bINI21DMuPod/yaUjMHvgOrA8R4m5R59oca
fkbhBHRqYaEwqzG4WliA+IBRUrzNGQYrpwT9dMaGeJJsVmyEOStZEGbambiCBIPA
dgr1860YAupjQEe8yMGuPTEgVXOZN37HO1oeXfBQuxnENmbaaGmov+51Q89Et+rR
YJciI9LKBMBkAjZOvcqjM6uqR8hXjySuOMYFuszIBWAV09pssP0u/n/hozsAySGu
dALY/98YwVjKY/5hPOfrhZhkw46cl5SupmjQNAPyHxpFZ1DY3e99RUIYypNeP1ie
J31HkIXmBSI2neQDolICteY9nj7vCABPP/VO8I9pv5YqmJnNHKJLD2AioNGDQ9l4
j79cVpWPee2b1Cvq2zCMl8S26PTQApZuSA2Rj2S74l2oqcLd5JsFB4d+4nz4LNQm
oEGWz6jQQsKC1A7pcZx1aVCdnHwo0Ls1z+amyLyWEHqoYRkdZjB3ZROvZTksQO32
Ya9Fp4Z8EVdiNU3+I3t2aCyz6C11+deLnBrNSQBXkv3NJUYUtfZHwyJFFyrD0mWU
xKZpghLUu6dy7zpucyLX6YjBPToLGWq5nvJUfIHkxlGpoV4fLoPZuhTK4aGHOS94
qb13alOXW+kD60ZrfT5L5lvYUCPUpxYW77na/4EIBVWp+KCKx07D000Ki63rj53I
pdNYQAKOHqCD1Yi+n/t2+2BVBOGJ4g/8zxJ47jR3DHQoZIkvbk50T7quTO+qm/Hf
+HZT8Bj3H3BHmP3ImLjENWd/im8CEmeVH1gOVLOCpz2wy/HSh9+T/DDIebiM7bdY
/0yYF/hgF2oALJvbck+hTODouHPAlKtfRgTuyHW+zbZ4F0ZbB1pCI9/1Tt0fd/9m
IOMGOC3d/EE1kPpqZTp8gj6JFpJ8ZC7dhYygkSay+Jw60fMFIxzAdyjnHz4Q3DJC
oSQY8tStPHwbTWO+Vr6g2CUOrx7SDB3H3KTDFUD0j/javoTCRNWg/Zz+4gu+liyw
ghkBq30ee0YzGPq5mvXVZAXg1E1FjN2VkxylpvVKSFfKixNAaIxwMNl24gFJz3Xi
ltZ5n5Sd9/o8rLbVMfK5mnMY/xfyB65tsTYd2JwB7xNFIjxfV2ku5tczwOSVTAx7
dlJ+MYgGydjvrVpFb8GCovTmnLJFJFOtV/LTcP22PP3RoNpRahpVJ1IT+cxwVhhU
AGj4XyHd7c55hEe2OQu706RyYX4qlgaQGjy3doWHE+9tCaQ84C0hKhDxlcvMtGCW
lffUV+GM+JawlrTd+1xlDoBUY0WOQAUmU9yaHgkMu6qwmtIXKXytsxYDZiTYvsVc
GBXIjXWYruiB15Qkg6HV0jWWx2Ky/dWA9lv/vjcPTzl8cwmlgTred8bjFa8Gs5ks
RHQdRFQ2d5jm4gN6AKwccMlzVcIzbkfOmsompI3PzQ4O7QJ0zfdsJuiRUwTfOPqA
27saACP83YImzV/EXTVBRwr7qVLXzTtZP0s5Nnzbn7zFnkuAEsQNk83v0SQzjHhT
dchVJ7T68yPMhg7N0y2/6N3paKI+rWic89186gRxmcUUTOvOsSWoPALHWT6RyrjA
Zz1fVhlVov0nu6f6zYhL/8z9gzNTMvak9LnuCWQlaizl6I3MgjiuaRvpVpUBXHy3
7RMDEXuvVq/GH2ev8Y1MSxr68nWHPZHLEoG1Ksxym1arLSVcMG4TfV1HIjWsZlTd
8145J828l0SYepW7Vt7Rqvgo5jNEKrT5/HWOTLVBu6x5nOn1r66CNvCjInSCz7uC
glLkFfU2BsAE/6AtxYvWj8nJSvuUke/PhRAcA3hdhpk9uefQShWoUQ/1tpEEUa71
CizgeepxYVct3IN2666T+Q6i1AVg+UvKn7jD6wiJlG/0q5XLMt34tZ1ScVasekL2
KmXUuYYntqsl3MLjphWnma8mrhot6q1sImdVeACq/vwEP1cSqHZSeqbqWrRHxPOd
uNVWqt2z+b+p6lZeHP8Y5TNHnE+FXvfs+CC7vvmViZD43T56P0fK6HeQw4i/WYrg
Z02ZCyUuUpVJMitzmiALM6npRIMWwvCErGkMEOB8NGXC0QPO61F2AhFBCah/25Wk
ZXxIPfjefnulw/cKhreg3CB/h8EsxqwFWQPYEg6M9zDXMIkhgv5KfvGFSNihJxXv
eU5ZMJHBXGA5BzUCsfMDXDG9PxsZykLqB+5FFsuo05ZkAJrJocBHQrjg87ePN0Fu
E5y8gVYZiLd8ZLD3hzeNW+sI9VrOcYgPkqq29JM3H3zxueWoGuOAPgj+hQ9CyeF9
bafXhDkPyJOGk5zHaElhfCG6RDA5roDPGbRLez8k6Oqhph7miBxcFrEvM38fpJ0j
Cpu62sZsaigu6lUV9kMfneQtrNXTrKPH1Al6CgwFM+7HmLoAp/rHXKEhvF6KNoiZ
SygV2Lksaz449ofpyJEwphDQGpBQHuF53VBY+jG9gD3v8COOTKmYedG0vhirziLe
gL++VJx3AzX8KM6Rum6apYdXqmSegDWucT05Zs5FRswb61Pec8I3jPM5RhuQU5E5
j7tXtQ6veKqOShygqO8mS+nDI4TPQB1cee/6q5VFSQGoScHYk94cDDXxn7OlpT5f
lgO/yMc73t472goOVJixkRv0iOCpOdw9agXk9OZ00V1VX2BibwvNZXUCtqhEswgX
t4Gdkx/Ud0rhjLYaKU4NSuHv4QQNLQ05f3ZcdMF47qYgxiS2FMT1Aq0dcx+XC0qD
GxvWmy3Na/ZhYwX5I5TwPjVsaSFwyDY8Xyp1O9PKcoYHsmDpkCRgVPxVE4qWYlb5
TlmGYhcxqq4L29BGfOi+ifE/PV1Io30DgkTXCJF1vEzJ3zUixM+z3/9bgDrJVo60
Pn3iV2onmNidOwzvk2ivGCnNBjFoClWNCHlm6+hyO2sBxaOSsIIHTg03UoiiBwJb
B9Xh53rhJWKzQrINKsLqpz772F+dI0/QdNE+bSLyWt6wuzQ/r+VhRjms2RhMGR7v
tJfFpuO6ehF4oTZwQi5WccaN7ytS+5sbAB3Li5WdQqZGyEl93WrDet075vH997KI
CiW4vmKXtubxdFiy3yBthDPTSOB0sI3cj+iQjpgW0Wx74Nu5n2nQsi8GS+xibsLa
M1VAc83bGpW+asgFd2BZPT+5jAWELatAZ+8SbuNQHAXn+v4gVDorj3VLGSOtd7ev
6iFbQnoboyuWsxzO4Ox7oVpOSHQsZVgLC4V8F0qIrGuASOB8kHVUA5rMB8suCAkE
pooSV8SUZRvfef51N+rAm8DKCF0HCiSFehXKYREXjS2VaUFGUOuFGGX5r7VXR0cS
4wQ2QBCuNCnALDbG4+Ssv5mqsg8HvVLw6jjQMnTSt0p/BvxrByKZEuc0t81H77Qm
yIWbk9y5WlvDV94rImNH6c2Q979FXB7z7aSy9dLKGruqfJWFiy5bgjDADClZZvmI
Q3LAsX7yWudoobdfJdUtdkZ/65ZqYeaaAbgVuhE43CGXSkLAvG0bsbx9qtNyziTd
G+r+sQZVXeApF7tfkFUD78goCJLrLIJpFRxoMEAkxrlwrbfT0qq2Nokq/uyG6Sep
VXNMKkNygs8ihg1rsZYph+fo54QrFunkLmo2BgqCOHksWkBW+0CVegXPAHKRx63k
WOknxBF2kwATGMHa4YZl3yURimFFDlVtz3n0DFTzbSo26eIkst1cHxbuNX1On4Pw
VjsjBPUSAd7wmvHgt7qf9Ijmmhgb9QipS8b7Aqpg8i0khC8BMR7vsD82y0ot8idx
4HHHsJ0WxxcqPI/OV+7yfrYfPdGwyCIu/8pa3alTf9XWm2gK0/ltqY5/G1Ru0kak
Gm+OjKleIe0wNpuBzMtjXqObAPG+blF82PN7pPEdTcyopwXAjbzfiUCLXtGf8v1n
JykPTtLF1lkrYVsVgd6uQ9uUXSq+AafiUleZlOcZ5vefb5PE++ZOvBLYhC6DT63l
x/KoE55dm9txWLjnEYI2/olxpLAIR+DxQoru2XzuPzJqNDomX2pX+qxhcvu9+SPq
dmu2RblUo9+RY9ODvuoM/qC+bO2JpznnA9NooTjOS0smCSyChV0YX8HZZ9hBCf45
Se0rMEFwX4nSYSKmuoVj8yZvxKjiXhY4fEDh/MMnJAoagqKwxZRizvzOBFOhNUQv
qGTC8vckIPv4Zdc2Hy7zJ+Ly5Ksi0cqep1rOQ7S1UYciLqZRVNMWupsyKIfS+f+1
+UMn0NE0De3iJVW8r8sAIQPE9TJCqNEcy+/revarWhecjeRyFo/xNCmsa4r2mfxF
i6T+NV4Rp73KB+udnEsgP53R2tUQJL3KyWKeIdYKiJ0Ufnt9qPhzkiObuK0zpeTL
jXYjkvJM9tPOv/1EfIs04vCki9212aC1X+vlS5T10TGKpCG4n4I+B1iGGfrIcqxL
XRUEh3UcoY7rHH0hljd97nxdFcONPI0sOgIXXT3TOyRmmYrTQdDsoCF1GMlI4ETF
s+4R6mUemGVd9U1Glx3RnKv9nFn+IiroJrtmsnFQcrtMrdfQqf8fmqTaMiyzfiiJ
Jp8Eql7Hz35nMv9AlR64KHrzDSwyoFvfoDj/Yzw/25TvzD+EvDfNCBy/qTK8w7dY
Ubq2jMnsxZOgxY7yN2v/H8ESyCqzx7zXvy8F/zGtSh0oiHrXMxY//lOtmBtxPhZs
1kcVHZudjrpmbFlYHQk1JkSwtY/uh/ZU93MePzoA45dWvdmjKfjCAijqdIXVt8kf
`pragma protect end_protected
