// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KNllBRit1V1xWm5tI8LlhPhsBdndnwK9966teJ+XENBsqITHH9+mLYDzjS622TLf
C8mgFeTVz9ZzK13uygRGA57VWJja338Rq8QcukIuI6s42KDhhqMfxWiHJW0z4T8B
X9lHPCVhCNqY5AWco9CM19Ko5EBdAl+7nVulbz0ROsY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 123920)
F4yfeQu5Ropo+lfIuObbVVdiEsEF51G1GosMZ0t8ZDmPb008d1oXXt1aS1WYI6lp
Tp9Ky1HI2LlK8ivf58j1UZ4e/AC5xr3SbboqNQSJMbT9nlnwnIK0cmrz/aiN3ikJ
CVFMSFJd6SEx2CYr98lXFL8j3i1dyMQreEbvKQXz7K1a+4C8h6BKt/2+SHBByqag
1cbUP7LjNCch0SZ/QsqNGBWe5pWCYCMuvn8q6O5++K91Qqg04KBIbiA5Xwfayr/5
sl6G0zP1Ufp1JwE4des1jqOSScnupCoUJpS41IAWKxkQaYLxx6veO39G31vVrt8M
9jTjjcz0iHnzAK+6hyTNPHt5M5QwSXRh/ViU29VDCDVOrzuaQtQpeEbvXSxue7cs
eBdBzeNVR1iJJawHqIET3e1f8zOGSN/uMPnvJBWOEBOyeA0W9eaxwlUfzIr2wgJV
IK7qKpmuT3CKPGalzbzr4MxXn+t8FJLgRH5T1CwKK4ahxOTOKoQ/NdA753u2GzDn
qQxXPuE5HUN7WWGMrG2BfKuOEYa7mSvCqwnNWcmYPV1yKdUhs49bZu+vWwCCjePr
jdZiv7fXPzfZY9/UqAJ27/JW8eDOO/nihB7+jE6p972FImpxDvge0Nw1jlW5SvBv
rmCIgDdtvBQR45KeevYqrMGWXXjGco/43rCzdgoCydpPJRk5hz/8VZpJ/eWm0Sgs
C1oYStQaCIuGC/GNeB/R8MRHMc2fIz/nKmNCBa62ZKBHz/VDpORe8z2Vko4cl8Qs
+b2TUvsJc//RbeeIcaKL9H6EIO1khQgGSLTqH/nX1ocxJRS/ZO5HKeTVdr32KnXm
/8uzW5Tt7mVa+LgcTDFe38pKO8qlQSIOyQa3ldy+tyZCiZhABtKFjWEzz/6oCWch
9guzpKUziVZfWT66hZW179YQLAm8zTdyh3gihzFpK6CCLXsOHB/3qZa4JJFLOgwL
4NUOmv4B47vN/TknX6seQbklJan3nZGl2Gr/GgQP9Bug3ilxc0l11X85cabbFxuA
OxAi60l5+s0KvK2OPo6YAcbuksGD5Stg1wqO+oZJgH0EYPW6DPOa4Me2UFKONn4z
M0xqIQStNMds8l9cl/oaIIg/gmNv1c9pTreKjtwsxE7suaOXFbP4VRto2Ahm6S/4
aMLtvE81h3SXkrHBV1rcNVpKUdCSfbauJHGpzh8XbjKM6FsMm4YAjPk+st6JD7kO
r3TyBGdtEUiWMBhAo5gVEEtbzYbi0Ib9GGGLGDBdCxGdzqyaAieHQRlKqTd+XPWh
9SIMBEdN4s7WoRFzAqLVXBb7Bqdz3FipEJw1y9yc81Blk9sg/IYPKkv7sEud5voM
4sgNUQj7rmqJbjnONdSNCVvEsbMpXnjfRkKaIBLTmb72GxGOx+9ZPRwEYBQk+2Bm
ZEwcgYrao5MNyCsMxfr0GjbQek3a1CUi/0kkNDuqjWt3Yf/PdYgNwo3Mih6zxD9R
bj9zmRWZFvR+EzWWV8b7ACqu7EPkXk/EM6xtMhRqO9tgLGO9STmPlmwgQmaitBS5
mrAqp5pw2KSNzW+UdU4M+y9yW4QKmNWDndiRZMAmH2TsVj3iuG+TMTNtGfq9B+7D
Fvdr3xc+I6dwwsAmts7Oyf0EZmzdyCPYKna6F4qzZffOweqNrJ8N6RvPg3KFeOBw
0bGw2jKQsaKMQqYRCjEG+h1CmZpANeNzhVDwU+Ecer3Oq/wBsTp9vEiWInYxjAwS
pbz0nnlYiJ6Bw44Kpmt9HQxsLUtReQi3PIfUARoeDiR97psFG6y/0eo3DZbdBX/w
Vogypwiae4ldQFy9nhGSajYWyXznj9+KmAvUf1VHmdXWFUklebq65gjC7ijWTihW
DHsnOqgQL7T6NSztaiBBD6xkw9meL/3gB48F2yIuykhOL7GdOIc+0GUqYCkj04ht
F5x7V6sjVE3H6JVXqeTnONzRRzviSUoOaSth0m/kXKvHWLNzEdhWRohGXNbEPRCX
zDOfro01isjM/73Vojh00Hcde7ktC3qRV06tmRIC/6Cdg+lZIWTtl91t3TNKr2yG
ffXd9dK36GxKjivXHsUFLuiNsCjftJquzp1fwRGPljPJkrIz9j3ppuIhe5Nb5Z47
FbuBF2PNQdop6wY4hRUCHNjOtNtDreavXFRiimUkR8ZoAK797/Zk1ol2cuSFmyeX
+61ohGnkVODgCVKYQefD0m7WPo/dG6PvRdiJkDI9FwUCwpTVHQiXnL3XPA1UXkil
/QsOa/pqwvvd36ysdT3kGEVe/5W5LDl7YfLCZEJnXlMtFTHxXXxXhWZvV9EsJlnP
awU3/J3dayQ0fBi7H1k/tA/Ry//4FYaIMW+8y2VBJg1JYT7IWvwa8NVVhzDiwMgk
ChwtjqFT9q9EyIn3gbeNgzkUxWNJJNAFAWpPaKxHdshpPm+e4kNTgh+WBMZViCsN
E7MRHQKcbdkHPxPhyKQc1rp8TUzaaru0eMLG1ecWSEkdgbxPc+O+kK1ukiITQzb0
nWjIcE7uKrXIvPjn4fBwebJufah0017SpLPXtyVQaCpPEJp0p6oJTsmybIEvoNSA
be5QrDmH4Z0VOJNfF42wPA+u5hFhQm4wqUeaZo9kqjQ6xBoLTzbz3kY0fCi1eDC4
lLG6LsE+eU6BoGjFPaN711q31W7Z/kQ0D5kcmLZxrcnnNWr0iO1QivaHnaSs45R1
/ydSo0ojQgIRcAsRgJzA+2xNoisrG+kJpHyzXxod8qY17b/LNcDod1B+W+w+ZjKD
vE//e7t57lPuyVDtft2V/x+5sKcLyfwEHLIwdpHxZtgLlm8rKaBreyizsgaxkZi2
Nsk6yGjRv3AXL9pOgs5ZaK32JfOU4oDQiSjYeiqdVusZslqaQn9t7HRWQF1vIByB
DhZzwuWJVhYc2qZUvxAXWItvvakL44enTMHNcc7JzlfOavDN++ubmz1+QxhaXbS7
08KYSt57GuzsJ7B0ph7wSuDEDBHAmXTqz5C9q2Dg0RsiqGzDd/Pb3bp8iHMOUWri
TvXA6pp2bWzUqo3K6JELgTsAu/3x41OQVNHJaHCD2mIDOEi2NkpxASzEw/KsdAo9
DEf/w4X/djg31O1D7VdSEou2cewyfGwzGVhGT3C0snQaQ6D+q4t2s6iMoC8lx/Ox
Qq8DcP2LBX/uVS7MKRjKgGPBLRhm7ZRmg4GG5eqDXchaaiWKRKZnDYjWqZRL1soR
jqCPKhB81Tf9MQda1r+hvIjfxugZTyzymnjQO3QOKXme6M5TtCrAOAW6MKdiF0zR
a//lzlPkYRv4nYSvoOfPiAPWSqqmz/CkgmMo/uO4cScQkAykyNXF7CYnlSXqCWIi
Or76qxfFG45zctXoYh26UcoBZhmcbC34W2YOVjXu5AC65KrtENXnivyEYcB69BaR
VW3zff2OjIieiNfwkuh2tWv3x031lgpdkIT/r4s3Mi64bag1P8i1hhdLSlQ1R7GH
m1B10pqMxUMuSVNoswmosZ5knQ93gAOPg3rXP9/gXI0sMJ5u8lv8nu3OzRI1yRVW
qJglAkJUApRqL4WGdqrRFD9vJrHNJiPiZQj8uq7RdwUT/mmQndoxXYSG4w/TK1U3
JlfinpgBr2mHAzZ4dgWrkaXT0LS/ic6DuIAwganZxZwjpyAFRICaUV9sY/nXfQgn
SUtSAOoHsqpK3rfdVzCd4Kwrk2d9bgmMyvJRLs+PsOrqgzq+d5uS7hbmu9DFnHQl
54S4wJkLukZrSi83hoBkMz/WXEJneEbSRx67/sHvAKBVcUwSrUqmacKpyI+ic/os
2jlKg6tTarOTF8y0nBar+ukEnP0oafffoSVztokB1UeX1TqY6eF0PaTZTHeQsCdD
qaAJ3QWWKnS+YQEe/qSEyy/TJimYOOtOc/E1u50GrNUZ7uXI9leBNtcF0GrMZjwY
Ocvgs1ZDOcMsnFwuI5z0AuUTw3UsDmgSApPxtvEPuyAf6G85j01qY85Cuou2+WqF
DhmvIs8YAVzDIA6PDqU8Z/USaOqf/fKi+6q8BzMFyYHVMgMDqDafQ0W0QiapeePh
akHGqcBCRH/S1xZl9spfBr+E+q8gpQnXgMeZrwp+xKkqMPa6MX40ykHQs5deYWhF
uSQpw84COyjrmpiQ+NPTgniKrWytg57QohHR6vnh4DiAMUr9UsMrUsYGIFZOZBKF
gToaw4JyYGMuY4i+S9F/chh9+WC2vZg8KSaNBHM/CVr67ctv1SR5Ix2x47zOg8L2
LZAvbkGnrxx9GpGotPASpvy3AZLrzFKiA94z+m9dmyXJOW8KMnvb2qKFrPRl5Jn3
0otekpPh1gncvnjicOfpRhjVbho+zsfWDhQpNMUsKglrlnJ5dutMlUMi+fgVidQ5
4KiIuV7urgym9e6zvDNBApS9K5S0n5xjZg9RPksFEeJwQciqEGg6UEKbptxHYx7O
wFuTpapR3IIW/yZofZq8OuZOLe8sztOxL0zR6eKv77f13ggHv5kvQtIXHoZ5AqRB
GkQAe93FJHAenR2w/B4c2udNKoPJucGx5qWW30A7gznxmKmDtwEQawzR6y6pyrgC
a4yBGWb7FtlryhMe78ZXzZAw7S+ugwbuTQoXb0WgosAVGRToH0YO5xRdWhBLMnav
2eW5h7K/Txrw6sGLLr5vVgy88SqWKSo02YCuFWIuHQpVK/R2YWoGrtizb/UTscrs
8+7Otn5P/HeUucWBCM+L9vVnNl4lmNrgv6BrwE9jXjv287RtTvu2TCGPSntCXoFf
kylEF5ebSwEJjrgVukmOKIajocE9UQ/cWs9wtrMQTevYhKAnXlielmMqf84jIK5o
mL3ulSlM3quiTBueGqhl1/4zim3V3lFOXSZU4EZPz+LkLG8lJj5iKK3TR/USaENz
4CUu48Z1p1ftowEj2/TVTDV0wX+7YeLiQ6DcsCNWqqo5CU6g5VrIxV0KlIOmSu66
EK7Ss0Q0/IMGg+N8Ph1P6S0UG3fwTuIPOGIrzai9Ajak2l0CIz5NkFBODKL9GPRP
OX8BfVjWoXsv7/Hxa1c+vs62P8R159VmQv7uX94jAhT7tnxNzX50AlGWHEq+6UBa
HJ5Zkw70U7OM0/zT9xu9D8ot9fYvsDXbczQ5fBtw+t6BAJZFP2hAoKEooOc0OjaS
hI/dAk009zz3XXYtuIZI43EzXzfQZ/W+9uqMOdiKCNoeLXkmPTZFRcSwPvXUwmMy
UUEs8X+KnqVwbcDm1FVURurGbNf6kUsx6rfnmRluz9KSexJVVPn3HbKACLrkoJW2
toiSGdAIRI8mFjr4EqN3cvvN9Wksc2NHDH51kWmg2RA5sFKMgc/2BXnHyl8TFw95
OdUROpWP+RHQcPELuiRcitxzH0ken6dt8edQgrIK3y8zbtoY68PjN0loVOSqJyUG
1SS0Qar7GSsucLaFo7MQ0tjJlnrOixDjohfJGusUpIDe5k2zUpPoae0nlWYILc6K
UDNNB7SzbSnVdAkOvPfQVtjy4m/nZigconFr45JiO21vJk+KZ6f0rgyqP90FXlZZ
ciqJc3hvNe3R4j8UTEM7V8ue1lpv17k6eQV8z9maxzQuNAm08+CawsqNDxC2JD98
qQb31gmo5GS+iHO4tkuKJ7b1CkW/9JlpIMmWuG0gS2C/UyoQ7LcQ12J4TM/LWH+h
5Ea/qaQ0JzurAd2QVusmDHHJjottpxyIZq//HWwVoQ4Vqijfobga2KIPKGBPvU9d
KpHxpPh2bkdnuxZBIJLa2/squS1l2k6Ah1p84wkXObsCE6QRxv5t0fige79dQlRL
k3tcErEenX5Bhql2VDvne0yxjc9I7Z1QuTtcs3hl+5unMgUen8d3voiGNnWaFCsu
1SFG3E0QTYfMYgskX+vDnBJNVLYrZ+p94lryI/oip5sbRh9BWS5c9p21HwhgUjsn
k5+accOtmMfIs9vivgHB5TwL1Zj0utQZRoPMQHE+GuKL6XPc3gg7hhFbq2GJ0f5T
aZPVHEPJxocU78RHRtI/YMDuiAW711TSQzHXrYwnhrbMyZyoZKeiO54VKn3ScJmg
aq3JsEovjsa5SvBjk5m/i3vrhof//MwCdhGiZnhhx1+STZ7nh/efaTpkYYYElQa2
4XXscehqhzN9/wh0iy9GXPsqv/fY6mNph/hsV5nRQW2juZUxMel6FkC9XcJwEa1Z
BNMVpJ1SK+0VHRyhQ7fx7s1wi8ZndEWW58oVVVeHoSfPgAfuS6vfvxY9/lu6Ehj4
87ML7sx0UL1Exkc0aMgHlAt8UorNtvS3Tohh9Zdnw6IBS/LGsXgRGPj/fOw7uI+u
e/Uvl0p4MHvXgDdEMh//2rFCFDrD1iB5gK6GuyXtAclqVGWLoi/FFZuygSbZUIqZ
DxRIZzFyKJQc4eNJ+SsmMOE12lV72BKEzY8fXD5fov1Lmzb9J0y0RHKPHi9uPXFJ
MUDrUT/1jPJK6CBZKUqL9zpaKnQOgj0POsv4vQpYKd4Ipy6XgAQV4NgPYheB1xb7
rtnQUoAXrl7x3XzggKySm3PhalCIlDHWF9jXVXOtU1FBvhfluQcrxOOX6iD02lId
W6IpvJ3g+KirW7IjjHfN5fV4gVFee4gtrVVsjPoRSuqSkAecuZEPu35k6OQpNdFk
dVhpYMlFL6TKcsr9NJ9YbW6EAwPTWOIRCnWLLglsb1r+aVrQk9I1k+CnRhzsigh8
jC2in3DkKQPbpgUcgKs82nm/fYu3F9tCz3FMfiUaCOuaD8sCktNOs5IFCaKYQB+D
Jt/6ZX0HLk409hul3WcgX3uqHkfO7HZwJqWeXC8lxaG+uCrAuFzVIZ7LWOzCBfry
sWJa/EThow1aGU5VRLP654nDIsiaWU1ArwIVtDrZp+dUHFY3JyD7KOoFe34K6vq+
M0cGg5kC+goljrZWOWeum0lKl/WdwihPJj9u//VvGYzzlul6yc4v9JApH5MVU298
tOjlbZMAycwb2yJPeAnJrUR8Vh9dqH/KG241uj875R3fvHrjbaiFjIeXaCbG8s2/
Jg5NhmmNOH+MAFoQNXDzao3thOwZ3XG17T/BVscyts4zWj/Q+fokJP0+ecWjNmkH
7dndqtVkIxo8wbfcTxFBZ13PXP4/TxmbPlZu5h3uDrngInH83Xydjc8FT+n28Nxv
TMt640f3W5DbRBJCsYZxurxF2EuGRRLm7DghqIYtB8aIRFmXt/1rMRlLXKx06Ssr
ZEBmj4Tkk1tV+FGiwizLwJmvkU9GDfCoqdpqHj8W0Vmd5PcA9uSlXJaXGqjPWunq
UChP0mLoFVK0ZvTdhX/WE+1XLH4Rsy5lTHAfehyP0RaB5Z0EyUMHv8sfpuLxOQzO
LX4WN9VsTRfBtPnzRKkxtrLY7Nwuv85tClfAC/7YjLzS/ZFhKYvX7m4jm5MURzd/
L/UlYWYxEYhtAQ/i9MGaAyJpAXf/PAVofLmuHp1anr1j8Y3eEa8tNNJjZ7D0ZAaD
+9d6WlnGevGS+k+mTBHmoS46MHOmGpTxtDesjE0cwA7jt8/K2JjI++TnUXfS2rUK
hYHhjQIYTPFXOu3WlbIrhPXUGC5Jx1CbCtBhHZM5yAFYPf44PwCjK3iDkcgZTQaZ
mSmbgFBo/ut/UEQyaoA5HK/1Ep9HS6Y6R4xoS1yNIIcxDdum2pZAofd/fba0CpXk
kWCmp/cU7onhPds3pfvhHzs7KB+xMKikzUrY3kcRMT6VIQt1yJj1Z9eIkzzJBDWf
zLU1RhBpA8AWXzjROI1lOUVrcmBX4CIFG0sLsxHMHQXjZ8/98UTG9W7PwWQ7Ortr
R0NTu1SH6QjE9DKEOanKfYmtkdlWUiE28b3HgV/I+VyZXYQ1KLC9vMbmaarxn5C7
hxJRZyOnek3YRIhlTdtapZn51OTOIEMSoYQOOxeLKQNxf1k2BIB2OPF24EUikpDf
0kq9u4WIJGVtW4sSB8unvnPq7egt/G/E3WtZcEQVlYuWgesjvzOXEJMs4CirA9N5
aOdWG9AZoZf0rMMXdv9/DGQ1YaWSd4PVjV+994fhlIRe2IFdWMqgULIVZJ110l9Z
nDyxDERbMDgcwAFtvRVn5bmKgaJu499vG8I3gsYP210kdQxVBxFtfTU00Y2ErGIy
CG/T7udzLTuxIxm9mW82/9eQ1G00vQZknG6NBMec7Qbs8o9ZNJWSQlLcm4STRCQm
JWwSorEsI80oVBOWIbJqjAWwpHlwf67E1IkP380Pvw/xb9hbkJlS6FjjxUZ3ztoJ
THskioAmoUpF89ZwME3Vb323B2v+bnvrSk3rXlXMdwldcPUJD1w3F7Zv1hNFvmD7
J+z94vRdwzCuMdzwd75YqnwM2FYlZbMM91cMiIlrGJn8o+bas79PgaVaFh3QLfaO
eEZfgXIJnckhLuoGiVRk/RY0x6XwNLEuZnAg7fkhZUoBb0Ux5OHcLPFhYw35yqWc
fn+pPEBJ7WrxSm+R4IXGA7YqsQhzPhVjuIfaFIZoEi3/Hy/o8XQYVcryy4oeyNCp
X6WZdiB86I7bJtwDb6xwOL+I/CgSVIDUKWK+2U5u8P1WX3qxpkv0XqRJYtVc1R1Z
N9cIUIC3CUXE42dKWMDrRyLJtKB7/7Fnac/ohrQS6Cs5sAPHDN1UXKfqsOeI8Gyy
9m017sJz25BAgrz61EFBbqWNO8j9osA2WrXtA4ZH9XhYEQ9WQ9hpRWMF4kYiQK/g
4Th6ojo/R3MUu42AKPA1AtIzzWuES35q+k580a1/bOkhfFvTYHEcs2VqY8VySi0G
Kgel/+lnL2SYT2i38CkwovOfYvCcGjDds4iFDF77uJLGnnRuG/QuNieeQS5i9Trt
OY/Y2cPGNkM9Rhk15dyTwvBXh21NZMn8U/d8yFsxRxGURNTnLPMd9KcAEtJuYxDx
EiZWVX1CBeYS6t7chSCW6vf5cIVUM/Iq7gyum0okqBHLYxo4OQFbRV1Sv0xhSD8A
CqJmvIJVEAkwq16aPCtXYuoTgOFvC76qcQnMe4j8oWPZnYBxnZFKMpNm4bUgRLjV
x/jCkPswIZ9oPpNgtI6gQxUBFc57rO8DCPageYcqVZgOJod0/dsii9aSRVMRKBBH
3+7ndMcNn0BKgsQrnZr9N9aoELgKfdCzwwov0bvg1jaT19mf1mSKroruemf3cPHZ
0kU6T9k+OeaJ4h/pX3qA1SV/ch82NxH9+L7j6E+x78PFtFFG1eGtGP1SnbOi/5CQ
9D0NJo8zFlGwklW8NHVsdm1BCIdrRKMcd+StQtH+AeMYp9RfDbfn9DftHrEOMiPp
i57qRld81/zfhCzxdwJ6qs8H9lKdiVeMHtuFyWGCYa88DPdbwMUSySIpajlKBvme
NwGnqcHS+LdHte2d6xdi7TmL8eMWPir3220MuhLOlFdcBi9TgwwfXjeHhMMr4qAw
lbMXZSVP0mMnUzVrBWW3lcxQm6gQRXR1700RfM0OZ4NCfPK+3WWfMD3fQvrI/E8I
MVaS9F3Mwz5mz7xc92je467yf57Vjpi3cnTNEZDfcTjqGXgfaDIH07KgAg8M/aZf
ZOecTqrpBhddW54JV+xk8rfjMZCw18KxT8tohm1kZA+2F2DB29boRFO4jcSDfdQm
yYuVat9mXN6biq9QNVQBtMIIPc3IrzNcj6QpMaAWSCL2VgZ60aYZnkAIX5iwARM1
yMM1uZ/taPZDvSWPCbIF8ooo3p589sRVxS+itCp6JxXLOBSsCo5zgV1Hpp4XWdpy
7aeXqFTe80fUnyJbzxEkgeNIEnIXq/mEfYpzc+A9WkayU2pYq7DWEa2PZ4czlcWA
fSic21/XFrtQhySh+nixJX8duhbFwLqS9sF4Exnlz+0BZtB0nQhw8yVL9alX65f3
AXIaSlNDB8UZVfI/Vw+N1E6LF2xL5fviEP7iHltOvCPzFY2u8wGLTEviITSucgIb
QLjFdXt1hwzlgrFugYAjeWHOTxpWA7dy6IR7Ygpr+T7dlgCpGvtfoIKeWPRKQaXS
U3auOcdj/JzhY8thpHxXNSExPOaUbpGZaqfHQMJj2iPLIonsawJWOv4RYB3D9dKS
urEzB2p60oBBJHdtqYE9q4Z7ff4VTcW+h7hgj8SmB+eJYZTNq0mHAe5ZMBS1G+0r
ygC7qvvk/7Mvm6grvYFhXMlxqiUADqBJ8pOUgB1aTVdrtSsN8MrF7dH0eh1RuFHP
QpUdELS0vtz+0YHEStXWKgHvAzS1p0wpUh2GQF2/8l+9RRnryyjFdYwYAQZNcoDU
KUW+0rDPPjzSfqvdPTNFoa2+7AuIHC44LNgvSo9y4ESb7KutFTTD3w84WVTviD75
9rLpMxO70+w35NHbperEyR/BmdlqBnukE+xz1OzYKAlbZDMfG+YAGMY4aqyJo4GF
pQHA3fqwsrNJuw088OWWbCCkQsNNLR6bFGsQMIVyT/Y/XXIEAotUdvfJTBYNEXHh
H1OfUUthy8W5hOdnIYwNwHuj1zcAyNkITEmoua9wHFCA6GsLlskVQsGdCaoy4DgG
hLv7WuCCbTkQb7eQ3vypHqC2pnMAB/AjoHx2a6I983ivTc+GvaUNwZzpLbQ4mkWD
tA9bYC5s09kPZlcahG9weD8l6HBnoM6rgAmRuzgU7FeSNBgUlKV+y/HkiUVQqEGU
pTDjpGLYMoc5hwjejM9d/Z0ooFJFBZrf2VuHrTlyCIrwiIKbwORuKtapFyLZiI/3
Xay31ITJu0S0+QdxP28rH4AH1/OrcBOrmJ0yADnxUxNbTVICwgmglo8K3ytJuWbd
7s5IiRmTXKQISlqoXttTb2MLeWD3UGXzH+UsLZQCMdBypRYq2bO75q99Xi3yDZR4
p2UE7w5mRitZJp0Cs6YjRUJgD7VS9Ki4mWeR29nMnj2Q8nFbmwsjJ4g3oSHNGZo3
G8etd5zEu/R+v9GJiKtNVGt7aTSsU/CKo0IzDrXjPG+kwmjYvG8/jZYC8WniYGLm
8tXDGt2Q2Y7yWjiUH+IS7t1q/s75lm0EnbT2EEOjmA4wqGKVNpFW1rgtoTWGMasb
2oXCp0UvZL8CbLgU7wRoKiv3lkD3jsyiod/9QQw4lI2izdRN9Pj5qCFAe//md75d
8itDxci0l1t2isDz8kPDvQDKR4OLH++J6WvERN/cgwTkX7sFvt+CJRz2N5ewBi2c
7m+XIQiYx55RF0BeAVZjYiq5BVfJQsm63+ZiHb3AI/Qwgcvob8mRJOz5axTAEWvo
n8QfVhSgpLo+ZVbIgYvJePupNucL/dVWuCQEYKn47Z9wQCNyfVfKEYQFTyMCHEmu
utyenMkWqDnmGvDRwkLPNUwGVw4ECG1MmIiMZR+BjjALQG54+FXskOSF6UXiJNPv
djLACb+ipzPP7cm7qrppOlAMbirLDUQMCW/2BpFKXubMQ5SjAl4jdNwyMqMVu29f
RyePaMwpu6jazwBN/LHI/DrFxsK/T16IKVs80WMz4nrKk/t8h46ITV7x3+wHu+pa
K1lplqxv2tdqTZ6H8mWNFxrBr9gLPUSeDC8kp47PAGonV1DzgwulFlrTcKqY8xpY
DYOYC9NWHErruEZ14CjjH5M3wPuTAXJ6XWE95KNonhabeyZrSADAxX/aRcQq/9Ew
OTxTsiwP+LVCcu2cFc5vkMx+dCEMuKqQBdQOhyfQOwyzyUr2Qc3X/u1lVzzPkuTh
8Lu/QWS4F4XKngZZlfzGYeWaQUBhxCPfLGCKG9bmEXDY/b5n/fFhXhcgAfJgeNdp
Tv0AXDsWqb8yimgsOEm1HzxVRWTDSlsYx4unPq1S/uE/10fbKSXxnr454ZAYn7Jg
StPm91VoW/9h8Dzq9RHZBiXZ71v5uGyoSFhiqv6RPlRQ9VrcmlTuUQSIx/iMXBOZ
8V3jE97qPWKGJ2BmGmVOkNx+NTlNUdku/O3A3IcF4zppKR/5Oiv1vnJK305K8WPK
TNzPiAYD+KLKMBhsMKBfwEhDMiEPSrNpBm47aa93uN1JVBHCzRotI4G8MpXyzgXb
ZamVNV10NNqrLVB6HWT0OienjPGLEkxDYyzCD8JoTupVtnsEj+U8EJwkjL9hq1S/
ftvFDYZRrVOsXgqf9esNUBJzywYiihNIxiPr6qLGINFEqMCJOdn9T8JG0PSTpi+I
t1okp2i10oY1tD+8Km2UvuHcc0zX+tqyBJJlAWMy01jXII4Q6VwFXYOGuHHD5CeF
ASY8VeTHPinzS5hBRQ8GNimUn+9lbT7zfne9nNW0k+Vl/ULRheEeCNBuIsvhBvQJ
3t/rGnvsnPsShvG70TG0WzClxk5L2lW5qV2oS8I+6Ttp+ir/RzTco7VHBBjK73/G
zqqwlHadPDZ3zVzL8EhH5yti11KiflSNtc+YpZUQL/eh03wbE8xmMhGwymFMR3hk
ovKez9DzT8ofi64635AhjufniJ4ZcKBx3ScRNKSu2L/EWBJJGUFunwb/H43tuPyG
d4bTwgOgIB6cRrzVNmX5xqWgePsMSEoFY0b1pGVVhnD0lYdPofrX3C3xEJvaT/ks
Go2iFn8beZ2ZBgPxQNH7mY/lAWXevZGZ6mG/j2uSWbd9fUciPHqmeyCBmGpgsr9J
zUrFPPpORnBvKjJmz+7ytoMWReLgWlfvoivJrH4QSpuE3/WnyeQXlFB/OsT4Htj5
HYP0knGvv9VhMJAQiOuzQWslsWr8OrXfiGbhaH2glJb5VI9sd5MmVyOXl7IkN4Hu
6QSRgE9YZVhdEtbahvnORwYHfyiAyYhTLVS9lN2XiBbk1Soq1Z1bNFHfwuNsonee
IROz/6tIyTf0KAtnmD/dgZPU4hGhDYxfYO1AjsmoM5IiX0lRg2XqvB2rJW6viAH9
TTxGhcMHd3ebFwfpGPVQMA1zGABrnOnQPXEOmpLmGYrTj97rDOtkWwfjyqL3u+0h
Lsr+fJY4uR05VrycoWJn4eoANXJlVUUFhKKx3cEDLFapYMXuzdd0q7/VL0PNqD1k
EEbxmlQKfo93j2QSB9//Jllq/rZdldxENci//7/7oYNmvOBMiLUsLpBmIX8PznRp
XgIF5yyEQOqSBELgFb3t0sYPLCT4iMrhbavA41wEDOZe6Sa7ft+2VitctTrQ9e//
zOCOLZczPoFQkwDMH/alp4dWz/C3xsy3SxefQ97MqrWtamGc1i3Za27Y37DdDHse
vlcyzVKNR4RxV7qLnmEhxAraIgpeDPn26UMBHVXAdbGYh7iUwI9L3Bh7DpW/zjfV
Mtl74/InZ0Q0R7RFcpJGHYcY3yIvamGiZJ04zv3NoluPJNX6X9j5KtB55Uo3l96a
hY5EKJ68CB28kUsQ/mGIVz9e9NuL17HkbWuuPN6DtgFimdOhwyBcXot4kMmPZlIb
NbBVBFfVpRSODD2eesXtt0rg/S0g5kDhbygOGiezrrOQw1g9XlapLu4gjf9XVk/S
x1Q5bAU7854jsZahGoSUYuaO4+sHEgz1krU4mcsU2K1FAHF2yhrrImspnlVtcMsO
wiZ/lqlHqKGsRfSyOq0s2ODUK1MLlePSmby+Lfhawy5F4z9lTDylZk60GPD+mw8c
Effc9TyWiP2dmlbS2lexAxoblc3ff0byruBnfrYUr+JC5yp3SZImnG6SbbAPKpWB
76ToEuraekFMotYDGI9gSWT+RF6NM/1xx61dY8dWj+jJ35R5WKv/snEHEqCQhaIX
P+UQzdjTsBxrYw6cTaZDgNDRtxDKSj4Oi/p4kax4K38ft9UDf247GBQDTXraXCzv
KTygjjoEUSeFM0W1ipq4dMmCyYp8T67ytYADcGVsVCj5QRHYSOD2bFPrjMRzNy1G
smKE4PH2i7GnuJUSZgMUUS7Fuw70K3gYFgKx/WTj+GsvVOQ6PkIuW7vnwd90btbH
EtyLu3CS1yZV8ebHH8xxbjsBarmLCbghRkvPfzw/Pl/dqtDrmI/6cOYNQ6KN0mFj
y3lLnFEshLY3JyUXit8OlNcxutqqO8u7imBxvWwyIHs5Q3u0rh5eAA4QN0I2DJXh
C6c8WwIMLz3NqWFv6638zrDCqlch/iRyyVO3rdzB7N46b4/tNQyONGBHKnOCML0B
y9gMn94O4nawRFepzn4h5LA/YstME0pkraJh4xYjw/Mvd7gKqZgRdFWVJz4iejm7
lnhLZfZbyk5f5j5VFG7y6WbfwnQ8UkagBKBWkoNgTAO7iQcKEnnq6BOF5+fDEBex
+eNY5JpEA2bE7G3UCR+1RT+XTnR+EgCH3aP2sFQdmmdmSCg3uheTwQrf8ReVTjrF
JsGOe6rxNKtAu0e2QHhP2Jq22INRAYJTB9S/ncxBkLK+eIIAZ2vO3doITbMFKNoW
HnI8YgHaT6kSjT51+F6b3e2Ia1v2K/W0qsmqNKJcS+RKJUpuVl9Pm7A1fJDFIBT6
I7KPMG2qKsR01QZhjVMkBniIlZ9saHGY1QXNAHxZS/Bvkp6yx1HeCxQrY3oPONID
jcaMZQ5rrqHkm8mts4deGfvPv3c5OKnQ563Y2HQbH21gxPG0vJG14O/Wjaz/lUh3
KTLNxsdk1XajjCmQeqavgE66uAzAsDW7bFrM0W5lg5UR0YDxVsjM+lmScpdblaNj
sd4gL5lzXzE9J/rsAmIiiWb+vMJne8VxWETClS7KdvGqT1HLB0Be2tG9/apcfMGL
hWIF1XsYxV9TdU28vulOvGQzzKTjvM/kBAy2xy0px1JHTQoj6ScwTlc7V+KZ41bM
6zLhtsSCigVLFzpAiMqyS8yh1nWocJ7S8hO8oAdRZX82iMcuPOFeGwLLpT52FDO5
PzXx//jY6/eI91br7okUcFAnhHqeCrHOlqJqgkrxn5FOQAG3ECHIKl6Y+88dLrhO
Rla1eUMHSVJV43bgIT2h83Co8DPTnV9DZw1T5VJQnt0LXtQLlzBHa+GgGfkBTqcl
eYTNKjaTsNP4/j5RQ/I0W4P4gd6Sj3wOrj/crnlyvDXORpqgB+geokfsmr9EH5gA
dxmrIgTt2lq1CrfNdr+1qM8afmb7i/dwVnFP6LTdrK4yw2z15GOxG/+GSaGWk5er
lGJvb0zMZ+Gy5nZKwsGueG43JY4i73ddmTXu5JqOm0N11gSrhNHXyERj942oaM60
DDDXVkL1BYyfE4+QytRRxu7V1ntW/H14mF7k2gHonP32KA/fshC3UXOAnayLmucv
X/wFoWAesgB+q4+5OlXC21AsJNApRaVl2i4ZjZ9X6NsipP2KG99GRDXy7gczIvev
AVSdUOHnuGWsb4/OGQqqYgHg1ssi5PfhatbLFTwwEpDVDx61fCcX0Y/My+J0xbXn
iM3Rljm+hZ7aLYv8XEYydA9EQBkURK58dwtqb+HNs4G2atyWLBWMDXU3saqmt5rv
ISm4LS3zyiOpjgnObKiwF2lBM23D2vNntsYpP5LL3e7Z0TyemjMd9oCl5rZp08d9
J6KrTnvJj7veogaiNKJzv+UYGx630I1/nwFCyJOOtUFWue7hpRdW6BwHKlRBwJYc
ayf4LRh2sGSMXdHVo0cBvibcnR8JBers6yYErpI6ond6t0GUkzqsYXAmEltNkQWu
b9Q0QYD8odUazBEnF750kB1uE0CRFhOCLC41fYbFixPnN0bdQiS0V84gXr69U1nz
h2y5ZflCwHU6yEby4i5BH6eb6XWxKwIKqPwsuUJxTp+8XJko/NTKuqQpyIo/3XXt
SxdlWsr0GIPO4WJljkSCWsPDV2fR3Kd5+7Kw1eAMjbDpS3I+xCYpdFzRG3NkuOyY
lgiBzvQmvQo7+EAjNzxzw/4KmS9TeoUXZK+H3Aqu2FgUacf0jNWnWfMQ4S0Y4nbd
5iYrQoHGchnIxtZLaLErnhYar8ukUjAnMkCm28ujInEOsOy2XHVzSEk8IRzSKXt2
G7PerF+nR5jIyfgwbRuhdKUEDJNDoRjVPqWK/UJsxB3nI1tMcg66X+7HuV4Vq9cX
N9JxL0oVp4ZXpNay7UL/XwxfdIBJ63j/M1BoWFtboHwoyKkrLol1wuNq7sfvr9jV
7/uIRX3RP69gkrozXlM2EBZLPlrMaR9ok6WzKmrwYBstHTgo7Gym9SlRd2tVoMp7
1s9k8xZy6oQ/3JMA3TxV/CY1SyYYRyDSbBh48DW72RcpJ+XNg4etkPoWCRyOdU5P
4iuQTyAYoLKjqzJ2WJsvOkwp6UhyyomC/K1CAXjMeKxFRuLv24oYi8Ddl4PCZKZu
jYVA3U/hJvX/xHbhDv1ToU9gQ1Tg1vXiaWTyxqjedskxASNm89yAMXD34XoLejrJ
zEp5lCQH2iD77mNuumLkM6HjA5rBKcAsc6sHON9IXdqR+dp44WYqwYZsVL6Bdm9L
LLNle11HqD8tKKgxMlVgh599vrxKADdf+rAmQl87+etMAuUIU0sDgUVIn/OtO4NN
/02OLMKUAZ33/iXkxfxlyEMYEtJslEN8V5mQ7fkBFZVb4AzzJ8TiJKCTLP+LV1Nw
rMFhAbts8fxLF+zGxgMIZ+owFsLpOEocWODymVZidz5orEo4MSK5jUN64ITR9Hjv
fU+RJWnuObOF1EhmhaBF8/L9kXqRoeG9xztTpAWyvWGSTznLqW7JHkPGKShjwsur
008eHtt4QVr6k5YS4BfacEadWQfWa+gUHYimCEyPvkzPD6MrZe/pgR3PQB/mCzOO
urPXvypvZ2qvPbhdyTqa59tzK/knkNOuiF+PVBEGmvzUYcvwargc9+rBMnjJeNHE
DY4CuvNXZ6yT/2UMfDsegMh9yhMd8B9SobEE7MoWlVtt/KQbncnz/fuJGtj3flKg
3LzdtoFPyH67uiOhOEj8nWLfGgxMEXk9MjRNyupgXISVhRa/8Jxed0EMcdaq4vsr
KgZVa09vPMncXnWl4+AQ0H1X8SH2ArtustkfDv643wLCAI+7AV+OCJhse8woYBkq
C/YHl93FYRadiCW6IjuYxuvv3N1dwu+0Dl7WsiDyXIEdy3xCK/qdThLO4e73b3MT
Ybjs16urZtRmrm14KI4Yd2jhjjnh6JcJuWsa6dbco9DJFvvu7W4yAYEX/HH2SXfp
alLSt2tiTuEx1ZQdRccyKYV2OgmRqjj3GdqtLDxjC7+7cNU9weXbQACICNyqrjjH
R6oIOHa08/G6p6ppfUdrXcAiwvJBy6IQfqIBOgpl3z0p/GI+05K3DVJl1rVSdfsa
D8Wf8EeUbK0MhUUam+VsPa+xpEZ8aUfZzsOBOI1U6moiYqenxcJEZmAIW7Cr0jEN
1zl3w1JfJp2aO/RNtbkEFCSC+V808/wPP6RdnKvTwN4wnrq3PPc0mcx4BlZ9DR6y
aNKABymaHQNOIr87dXHXLUXodePFhAIP4o6l3mmHNkMC8CRj5Rv2RngWYTGv044i
3qCZU517rpceawNZTbT+YgXj4XtMHCwYeNm0K6RcTw4Q3NSKKhqUM9a0Zs/ORuUh
rfKRJD6//5bHH7vAAc1WfceHnuZWOBShU0GnlbouOaBL5B4krca8H4oKFZdsuiSd
ro7J9KcwKB90b8vtoEIgY2UmJQvh+k1jT4ZZPgItpf3YjfXui6LZQadGg9i8pSnE
qa9XehMdTQ9AqM0Aly79vNWg3jRnP6kYho9HoLEuSfsgxrhxV/oalLE4N0Wqwp5I
CLC0U9GFFwik8SBvrxy574kLE9maPKa0zwy8TSletKs/9I/oPAMGpMdsGAsWN2Wy
RiXthKfMd8IyPpVGUwz3+CHM/CE1idwSQjVzYgH+byYYe11qk0Uve3Xy0gYujHOX
xfZL1pGov9MyuXCnomRkWbyXT/7FS7vjNz3uWv9rfu6bdGxV7IUn6RPvIiMI/Qhx
l1fB1upWPIQuNPGMmIOn47pkLgMR2/bkVgQE1QG/tP4YByS1Xn8Pdf5jEqcWV0No
GrLX4YCzjV5f5sFkb0zfwmcBZ9fIuT2d7L/SY3aqHr/bO00Af3oY5IHgRhTqVMPc
7SjC91aYN1REbQ5Ypo7jwMi7Vnf0u/Dy0XHSUSh0CvWbzBVIq+ThmGlu4YVcuvjJ
ZHAdTPC28zLvyx4Y5NxEIthhqcV7t7Eik4DBLnNpFUIcBeVkRYVuYdNKdpa3ntmL
zCWjL4+SixTduR1siIdWgLv4hHHFr0/3wnTEDoJsymUXnr2c+5iyDdT6wpBB4JYF
JeMxLXThGqRNC2J+uvfWYR+X+o5VvcOVhXd2Bn6Gftmtgoa9SSIgxXyPS5gp9loy
jYmPRAAfOExftaWlkVDrOv64TgGmombJuVe6q05HlqyJEBWxOe2Y89XLYlT3qYGv
g50Qm9uuvPOrRRMqBSReWaI8LC8OAQa9D0OZaa6e/KeIOKsscBmmbe+MOkKIOD1K
+ru+R7dhSM+OijqOuLl+8wNMAdiKMla7GrXCFiUWFEdPDF+uGVQK5364ncbAG4aY
2PiOx9Nl4EjuV/LkSceUDxMGNWSnRB2kBzVZPhnHPCtfAkMvZpPuBSdrkMdWFnwG
yYmN4Gj4uxrCA8GcYjrMAOd4IyQBbWmwrekZRRPMBip6c1+99NJhLMMHTzp+6q3F
8z38hNUIFrI2fqwDdsKO/5f9MPJAPR3Yl221Bn2wsfaKCBx0r54dJxx0eOjUYqu8
xvkMB3EdF6qxzhWJZF+2suQjrHbBiDWyKh7uPy0VK0jtdeJStKHJ/g0kzCp/ZDhJ
8iSn711nZTzngzyYgyl+S39kxc9ZzJH1/kwow8U6syTo2n+a5BU7YT3HyBqzVJ1z
WhhyZnVD5K13um+3Zv7RTYhh+HLP/081wvdyJvkj9CUGBmolCcDn4wcQsAJqlbb9
jFUwJCF0E7dQQ7DJoC1GpRcdfH7n4pzdmBQ7fKhFX2+JpJWOzlVR7UeXHAxLNu2T
NuzuwwUo+NGNj1mUxw9QGqLaexnPxf49fivW3fQlD+3cl6Rz5TDeBRKcLfgF4l9N
FF1hEUxwNYDwx+CvLZLveUDoKSvFOmPGopogLp3YYMeokuR9nghr+AwWaldqZYIA
fjsZkUzW7QH0D8x9WAcsWnTWEB8rJhVMzSp9k0V6Stth9DcGDlHxO17iohgW0BOY
AUzeZnkduvGPwlh2wYrG+HHUPuCA+bytERBnKY4AB8VpGwYlVSQVGSBnfp5Cn4Gg
P1fB+wFcvf/RQHTmvdyci+k5oxeCtVzzrKDle84JPTRoB08q9tbLGBjbpgz3qM0A
KkkOFoWuMZBVvgSkOrDADNH9dyZfwyO7BqnLo0TveMcDfGFZH84iG8j7oXMfXZNZ
bYBZL06pcQGI0DUnPaaPb8Bzzw0ctWHwSH5TE/Tvzm0lYLsm7NRjarK/b69HUSFy
DelpoNgtF/dqQkC3OKIS0lyA3JBB5IO1PtGgJ3yOjAfNBsqaNbBnLjzhQHPxXUbl
1ExARkK4kyPoiqFGEatulN3W67zinoZh5jExLk5sMWb8h9EGBEHIQCGsjokdF+Gc
vgTXCUbjC2yvRbYxvPwtDNcym9Nzv/jvwqXqbOmzeu7dRFrcGk7/Sl2HgpiUZ9u8
L7n/qwKKhyFZTaegyIvoQkRehgx4B+HYb5x9qJIhiMEukzbGXWjqR1psbtQzffHh
KcAojfDnH38hllIbYSDJ2B+SECKjY8DI6bLhluN4kcl7rz4Ercb3cOIngN7h2U3L
o8rpGkqx0kW4QFjC1ZdWlnaQvdvOI2TzxMcVVK6Hs+qgPbd2S5WdZebv35Pq/iED
vJcAEVYyQ24TDq0K11ywLzMIe9aAN8tWooEGlmKKyv828Yg9ZoKNAL0RpJHUEe8u
2+YhDgd2jJuUBpSyNGjA4OAzUxOyP/pLKldLnxl3hQ+WBdZAY+Hr+3ubmxSCO0YG
S05HLGkSwoo5O99eUdDBpubol3SgK+y85VRcdHSdjT8MKJdeed7vWhaDij0LWnlq
hr2OknbuWbwB31zzR54RSuPpgIi8tZxVh3KXu83IbGG1XmR93mafG2EO1ZF9PRK+
+L2GO9zfAaMOOIYyP9t4ZQ3ij9xKEc2K+ffV9nu3307q9wlK5p9NbLseMUOs9IDd
T8SHGa8PcM97YrshECe+kK1WIZvcQgVexaeUoiMrvg1kn/UprIKfC5/YWANM40dO
NIniFvd8Ql8UI/W2xcsD0hKkJuPJXWglLGA7TU0z6ODp8+mfbbOnSN7ez/QZDPkk
NXAri+ZkpMlfSDXNDmTVIZKNUYjNK7MKdHEBmbfbcZ2/nd8gyvmfuOtuXtlPONW1
Wv1GrXLsrlpJQGynaggq/tcXie5JyOrD6VJy7QbHUkYlzBgHQeTKZlfPmTWXgxt5
OBO5dhoBM7Y6bake6d3AynIR8//4byc8h6TNC3BLHb86fXROWyGCYuHVWIUlxmOn
8hK91tZ1eXbGg06e5S1Jfkt4nUyG/fkPxOocp+/hyzDIuHuW4rvUlTx2JsLxyY9i
EChOWK+z3IxS9M7Pa4YAWCRymTUiPNHlNM+FuAJWZrxlkX4sJ1Xu9w8CBzfmY0bt
2nLAWpVOxw0qtkFxbO5+WOS/co/gie50KCs3zw5pTw3QjZqNQnooFK8uGQgFcldn
jWzOjibUqlXo+JDd5S7kYHZOiDZxLMrTFp8sopgKFmo6A+uO5ZAjIsqMbpboqR5p
RUnibfMfy1HbKHI6KKHwGRtlqWZWQBGgLH/PedBPU5uU8585BONyGzG0qjv8LI9J
xAlo0jUx5C9qW3RVBSKNdLxlXrpaKRrXbY0uvmoiSRe2BpmwgsW90KqllnDJAiin
Cx+CWCAoci6d9IE4MSN4agVrqww0J6oNtZaMIfzI04utUXB4RyfMeSfqZc5UbtVG
4QQSgtJXP9eVertxmGWmVXUSmjJNXfdXRFB25QyUPEWgiAgUV21V+AQkbAO4vJZl
mfh/slyb5aKufyHXN+e7rGWF3XKX9zP5+mblcq645D7Fh/MhRWd2H4PGJ7BOEGSb
NQXMb1rnM4ha4zQ0Cd5hlIFk10Fc4UkIdrKa0/4Wgcg8r/xycJI8L77PBbwpCxcT
pEKYm9LI1lbH1NnAKXO2bQ8FvPFR33RvjTs4R5sszgs9XL5V31Kf5d27qYGK2Urq
zhiNbKrZ/d/rDnGAx9GKdL0qXlkBcSD1g5EWv94n3+RalDLGnc2xu8hCfNkYj++7
Qcn9QxDNeL2Uqc3RX0gpnCRT8lL1ntDVFjOCRwgtoJRD2ScPtNNq+DY/aJJPxgDo
DD2/qeKo4+RD6e9x9jaDLxNHh2BLS1bCNXgaxK2ZvaakjowuuoYwx73vJCwvM2mQ
0KET/Ha20ShC1Cd+ZrXMfhXOEOzPEFadzfcpC5K7JBfGQ+7cgHUSMWiYDHm7ZIdD
a0CsffO5fRIOniVD/keevY1Q93xQIrLJew4sfiF6P5sc3vqP6qyPNB0KquZwy8Kd
talnbMf8RrCXQ6BBcbZq2/Diujwc/48MtV2owWRHNabH3SBb3qlXGcNXLkPUhrIz
egeOUG1SAFYXvRHj8v8+b16kYTFWoFKWctDJIeYW1E8LSbaBIa5yMDyfB+RYWdV9
x68C5dXS5xsAwpMTm5VWJoV4D4ux6MeNMKxD8wlYZfZQbJP8mRcOZQ7Ck9qWvjKI
lWpQMrMR+/qvTI7CCsqSGPE7putppGE0jv78RISfl0IIe9u7eGUd5z3soTeohFNr
JemBzqIoOfqcKNchZYjHFdlKXYQ/SsnDuKI8l2JjdgZr9M+u8cl4jbG7AikAmm3/
XHPjzuRXbBoBk+D3CBLAavCbvZpeBQH6ZPWueAuSvCxWIrBSmX3xFT8Flg21kSEm
4IP6UwYaaFS2Jxbewd8AwFjkMdBxRNGvtnlrANm/ZylmYaOXmb3ycAk1/fgKJgK2
Qaq2zCkDomu/TiW2WT3Vtm1cOOk6mifhuiBesPdvvZdnzarVp8EvSa6POlGQs0in
AeLyW/DJQaBssVwDElPcFSl7VYChYoU4SG07SvJFgMDZc8A7wRiTEHuu2+0PXM+F
NeSuoQT28j7UYhNADIRuVXY+2wtDWMlG7T+IDVOF2+JO9UdquNclImX6fL6kAiW4
Lgun+5dKe2+AdHTHlCO7yNsGOi/Q/rCURtwlcMWfXDdbsibR2Bykg8uE9FT2pgPn
+KzYe3UNCrI3pao8pvuCPfBu+oLENbH3FXgp2P+DZk0/0ld7pkr/lbfZpMbFQ+zn
eUJ22zgvA7tBn1WFecgNR5kjnhIWwTjv9Zjp2ZfZZP3DUa42jyHhH7nWYr3Z6yLn
G2stsgM4q3akq9bYvUvTzI/LtHdOU/6KP3SWDTdhEH+UYrJ8uSL95RRqr9HZSr7D
/sSJhRlMC20/dFpyHlBGFk/c2lWBexEe+LLwtCo7GpEP0jobwdzdhANoXnJE4Yal
cSG/LoINB2UIOCyq4+ftUkdErMQthqRcXwjQbPsgdlUL0Ugw6rhS+ziKCOJJXHSo
c52Mgx1ozJxTUN6+fNyqH1WLsV6kICj9XGRQQnOSUlzuXgSLS15B4sjJVIgiN2Le
/iHzxMtY0QBYMQbVkJe/qJO2+6I4WF6cg8jqk9xvaY8oWBEryU2pnrX1INjWcX/9
Cf03IvJNU9CSYmJS81vaJhvngcm28+ySKi2RKagbQQhU8BLSx8Nrs6C+pCR0uroB
LglAyzdCicDk2LAk9/swh/bTEb2qxaDNVj5vXwXI5P+TVoJLOD2/VwTGj8tfJoIE
/ZKIljk0ja7CGHX6kcbbx/eFyX8jyfJjmjKc4l5Ut8+cZHJ5volzwiIt36qUofhq
CedczsBnaZlDixBL4q1j0v5bCkJ9NZljxN4KGQC47plpdtKAsYWN93iFTgOgYNTG
+gRpBr7/Y3YRZnRMYeMkTubPwiQJbhkIotinaVXTgwOiJVGLr+8eHeBDfzejZDSA
vGQ0fqBIvLnjS0RIBxztf5sWfVSTMJOVnusQrHfRKU511gshr4e9GoJpbIywbaXp
xZe/8vbWwpAIF+v7FCKudNE+H/iUslnb8GX/tZ/fha7XnFW/W+YfBCUT0n3yroyo
18kTBR7KJ4XLUlv9HE4MWNMQsj2phIRReqPG7PJbKguOOLl0Yhbv4RkqlNzj2o8/
Jd4p5IKez2KMWHxoovSssevvp6l5SbZW6RxbQzhY1q04m2jf3usuxMiD+BG4ZeQi
XNDO8ME+djcpmUEskldf4BdaZoBaDQHAUBeVxDttp7oUHvTRZ5mcV0HXq7IFMl9I
surAn5lnC4Nq8/77uoz453CcG1WojURvltCGf84nVPluuA0132bvuRgGDsvnWMbB
XOAZta42BFGVyaXK3Zm0AG07l3lMxyktj08CelrXCdFBldYsxrH5m73mH2lOTEs+
lYOcax1e829PkNkIWKQiFxTWJSJFYrGBQJTmlOToWlyra00k2p3p6dt0eebKirOZ
5p6zHXZkxXi0U5rfXb4KaHT1pv3VpOgJEebgdgJnpSUtpv5bhgOlD/Qc1GzOjnpr
wkfNUAKftj44jkwm8mmvw0rsEI0XlfJw/Yt8aVTYT2DEdHu7qwvLoftcP5Y0UT9p
D5jOOFXCyMmiWQM6YBErHZXE9M2aU8DQ4OmAddIJxL2BYT+Q8x0gYNFjjoOlb8me
1m9WsnuWWD9c/2jrZVvhKws0eBtgWMJ5ADx5F+WSXfHTRa1xUih3dtyppN0AKv7+
0SlEuajkfzpAZ5tqHBqM7bmvoQCRpEwgFnI1dPC4IQS7fn10h9rG6KLs2QD8AZ/0
zVPjZMJ8O4+QVM6Jf+H+rR5pDurFLIOR2sRCZ56f8SyiOX+wlDu1TWINfJBh3qQ4
2OhJ+sEy5j5n7k35VrUrqzDHoC4GAPVpy3kcJxkEphd1/sFIsfKpJ+3MjTLp4TJw
3cbaM2atAjnOio+8sRiHGaoQFObJMbALfrs9YhLrEvnFVAR2Fqv4oV5R4RyWy4nS
jXTAAHNx34HIcqzxWkuRSrzKQtkPuAwoDLCI6w/paX/CCcTGc9GCM2G5rfYcJbwh
RBkGCrkDUsr7pFuv8h0zFlcorPtdjD/T37+sVWkjrOvQddkhaAKamgVmWHOYGwV4
T+SulnVE6LuQyJqqGhm/LIpX42VxlnHvHRVgna1P9jSif4G+ppeUMlZR5pMM41O5
2RlXrkLT9F8LW+M1cwO0nC7jSzZZZ4kBt22q9DTV/GBcA2FrFjsZO7SGjxdRKZff
r+B/V3D3E7fEDXPqJeo8JdsqVPG6BXNM9ZqUqrrgN1fY+XshDsB/46NAO4p/mwVI
rjPniOA5BoCee90bzc/t4p/Hm+WZnegu4eTuFqq8OTcAzuUXwZQMcaTjEVWTF9ZJ
e0XdxjKgK+e3Eat62CHRwyEQXb4NKcIXpTdmmlrIBeswV8NINNErGyLbwym59MSl
Hrh2geE5vsEP4ie1E8pEAUG0kj0O4+Um0SeBAxKBuh8Utk52GzZ+gbhnpQOuf/OQ
jKyjBdcggi/2jC3Scx6dmUCx9mdb7ZYCBbefU0fJHyqHDt7SZsnKzW5IYQjCHdIJ
BJ+PltPDGeUzRxEJ7mmtYnsUV4PY9o1fgIEKtaDMf0hazfz+9mRJ/SjfAX8RME89
d793QXointabyIZ9NVe6JVyyMwlJmx3WA/R4VI9L4DxULaXOtpmsvEP4D66afNay
w8CN13IQSGwWut0kQBOZ5wJ62a1r3wdQ+LjhhgWO1XnFBBUgY7+U6FyPekv+TrHw
iaVBOvhLv0ZoxPOiOJCedwJIyK05i/s791+scBZoTEqCYfxVZjv3WE7t7pcQ6teb
/SVCe1URG1/TYgWkn2E73fPm8Z17AT1uAZCxsaoU2lNMGxkQXwoblhwiQY+L9G9O
o3BXUVIhGWrPsRT2CGscPKdWHJCSNPOQxrfdY7WbG4HKaTM3MYTBI5p+2/YlIWNH
tAMiVHuGhbhZKQIMcLjnDFNMqrOjnOpO7AeXSrTk/Fv6ehdN0NRRLanNXxnV6z8q
ZnIvrLaHfulgVVzxvWm4k81IlDEkXjhaPgEtuGjtwup0Un8CgGUwXB34/j8PlvHU
BkjpeuGjwzdPqTy7wQteprdGR4taiaI+BDB9a8d9F91eDlnhEosMNfnPG66UoUaY
ZeQ3f5nz4pYuX2TQGqSRQ/JkJUzfwdN17xjyMKCGnwUyDkw/UxUBJ7XHsUEqOPEO
fCa3+FVjMzrwezaDB7R/wRlyOjLIdHLZr3ItYh2Dk2GvbW8XygGh32B3aYRNFRTa
sKp6GKSMPJhZ+bj54DWQV3vomPGMyw41gVR6sTlkekGDHb7jVWVLCNPQ+H4MbD9/
7Xg1T8kdPvk/1EncAu1dgPPO49RofE6zPq7CzsSHvbE2kDILrLdeqNjUVVtZuiGS
XhL3ZKF7ZebN4TBijjd20ox2dVWXzJOkiQqcClqp8wIva8ZVE7PBIKE3yNMaWYBL
f5iT77fVIaoXSBIROtwwP2itF6Wkpd405KxOPvg3r1bhFQgFdBNW5hZK8kaVe1sX
Wh6byy23dq2sLbaLV4mfG4s3Kql1m0/vFHGWqSDX+HDwweOFUBGRW2Vk57gfM1Hg
sEAmdg7dgtcmpp8oLaO0JuBmKwthd9/RxejNGpHMbwKjQmEL0V1RsQZribCO+WKg
8qOf5RfZEUm1n2slax1DZF3YLyXHG9965hOu8FW9sNyet7lC7JHccuS3Si3kl/0J
9E41AwNWLZaJbfgx9+Bie/pm63gY4W/nSMGzx31D5+aJo3LNpMZJ+4jAhZ3ETQk+
fEjmeVG1N3gTpgt3sIuJ6knpFptJ5XMophn4cTtFb/QLKApsImPoC/Zu0/Q/6qbs
eogDM1kZM0pSI8bOLHVDXxVLp3gXu1By4p7fwKUYFx1WY66Vt6B58OwadGziiAE1
Xv77uqQVqziIYTWkqVjyTfqbqMPz1L2BNPWjM2kKNtOPjhLI2FMsrnNR+JHacl34
b3fIEqZ7qlHjQd0kIKKuhrTafC62AuNgIa/mHeENg8ggq+FU98hO/bBccsPhrGXD
Ns142pAkhAwA3dAu0VNZyvVBj290ATf2byCVXltLIjGPFrMC8az1QyzCg9rf9ula
G0UAFhgj9AUnsvHO/NhmxU5aPaDmcYfGPzFFhjUe4F3KgMnz8NM/C5vXVF3pppOp
E2Y45/roZpO4ziLrQsq26Nevs5rK341HOnu5M8ZpKiD0Ryerlr2mz801mZWV+J60
kkOs2LY5XcyAzFakjmhWseFXkmKEOcqnE51p/rY1q7DxNYnJ6CqWftgpR/h/QrMb
jE2nOhjeb5gAj+haHRvT1EQ2CRkprXA2geZ8/PpGoNS0g2QAy6iK/ffiOrixyAQJ
Zy/tUfog5UznHXJow2Fe4j6jvbjyr3oTHlbelPCwZbF+WAGHARpB29gyCzw8vAzY
TafIV/3uRG6WqyzcGwSiRr1+pHIVbDie74ydyBw8Czjhyy8/HFn3vJ4sJf6g5fI8
fzxd+RAxCgWEWZB3wBmQcBJUZlmBs17ZDEsydRkl5KjxyB3unjfO89xyvywaXUsn
dPZ+V00xZ6ZNun1+e764NgrsLGcHNbbNYdTUB683WZRSvetoiwLjUO+Nh6EDgSJL
G9y0lnR+leC9s7vtiwBNzZ9YOgNSYhN7LBpZg8yb96UMXRcR0d54BitPhhU+6mh3
S233TU/4/jzpbED5Xjdab2rAUvJVySs96rVvlymd2/Vet/c1X3yifTyZvoAaG7hC
ab7c+QLdT4kOALoA08lYKvX+ws4xCu02yXWI/IdH850LfJS/x/VFF/1+MkYiBfgT
5M31wBCAqwQU2Z0QTrAveHWhLXabRcouPXceYdX5IMaJXUJfoAKkbp7xuCqko5OG
fn6nuXkvxmW43gl12KalopUcvOpM4ZDeVa+NPHa4uMPzsgHadN5Q5LabmMFYghcY
9gnpyifActF51H//PJY8b9Q6U5oPkkDzXpzzJ+/XlnTkeKr8KM3Iy7/HEK/5quNY
fSDzoMvQ9qQ4Eoz11k9u54VZDISk6khkQtRF4zDuD62B9Ve8bYBWtiNF/G+NR8tV
Li03ru2i5pkKHYLH5l/3GBhSpjamjNxwwC9SohgPyzJz2fyLgGEj0B8J7s4Z8vPs
kA9yZo44uvz1ER9ED4cOcAargQOWD28IBWM1Yuo2gHee9uamktrdlUEVzXHRWpsx
XkcmDccqqrD0GF3ncT673fgWxMwpo95h7G7N6ZpBJxnSrlRXz3oH8ElA4QHVfIwo
opF/wfTUGvjmCrHXQpuVgaN5mnT3zQuu8eYATdqNwJX214DDPh9OTfCp981SEu2N
F5yIM4J3BrQxP+ySDITSQ88CxyrgxdVpFwZ3phjUKdTVy+edh+lJ2pVyRkYXuKJc
X9iU+ylxvcYUjGbSl+4hdRXJIILp2d+dDxW+np3asSSGV2qQOFAvTb00f8AeAGPM
mWBDE1uY300WmYsMgN+wo3MGwzHkcg+fUIoyc9nD9LCSIK37vN5EMxuzdH0Uvf/4
H/e8cugl3/6vOBT/sNRtllN74BqpGuLojI6FAccJ9Y9onqWHDl4FIeIK0DKqmXNs
g4+OVPYT2ft1Pmo47NUq69PvlgrL7vFqq817UlN3afsvmkQQ1J/rfbjxMI+nrSvx
IuJ1t3f4OS21KmZdANBoX2H18pEEXga0D1nCwg11A3C9zWpdx/2HSsd1LPGV/F1U
XT/TuhqJbo1tXks/UeYbougRWBLe+IQ74GQkQA0KN/Gim2Nf88SUYJQWCQ/pdBKk
zfhAuneJNtPBuCtoaQb0Grbz74PMl9EJIHgCAWzy8CM0WzbCqrfwtW5HWUo7OKR1
b4O1KcUEyh/GoK2TTX5yneFfb34DNCSyeoGQUm0J6gFJ7bm+m7EAsDAbrwcvArHo
yQpOSELAphNV58Carbp5ry8vXRE+A1D7db7qHLFq2NatTo4e69s6Kwi/XxybtTho
TcIQOC14LQU19h1ARysM6R5Z2Cee4OWJwHDZy2+RwZibquHA3cTz2gXLXP1sFgjK
c4BHzQsN5ibVUW/Juv1WLH+3MiurmQ7JAqWyclbbgJYh2obEHdvg7oj9SzHasZJN
kfyIDRZt+lN9P7MXlivF5M65rwieozMuW+gfmq4eUyBGgZOORoVdmea/W65W4lBn
pdutQ+RAr3Lxza9ROWVgLktfX92IlqYopet3295zLe+ke/KqdhxPTucdbyeKjdYd
y2YxBr44X+vbbiLmVEDZdzSi2vd5C48pmIeWcPtCwYlm6nxsOjHb4CEUu+zADq7n
6iL4pMEU7xPynF6uezwImR3+AbcuW1F2fICCNzMjWEtPMYFUo+IA4pGrOgrBP672
Xfv7D1Q/sFdAXYeumwDa5p/K43Hg656cdWBL1fvUu2SVP78jgJggeTlrjAE1AUnf
aWP8AzogVapsEKR90a5XNdp0rmpOZHyqbI1xMEuO0Vh2A1WzhTvefgZ8T8TbZZOe
jH0K+ha/7eOeQcf43/+yVm1lLMzQlz2TJjMLVXThs3KdV6WNRFjh0+UCTzSpqY4Z
QBHE8QrhYkqKOpads4hsRUlbk6oje86x35RQelN2jYuqD7QAOVSCQqlwCyYKZSeV
oBmgdJsq6c14KlC6ebvoEfJl5L3mUqpoz/WhXe1TsjhQp4IcC/4ww8G3RaZPPWor
epane90qwsHMRfKOJcVgxflWgMjXKVdjD2Znq7l9W8vYd3i4F1ypgwharMmwfWoi
WRxZeqLHe9z8iAeF6kcBK6aNWHBtp/GXb0dG3nhPOvGZJxChF2Ak4NhNPooP2eZG
APpaTVzGZQ2zN0S0QIXvG2YOOkjWjekdSBMRUkyw7/9q1z+fMbeXQTeGhyrRaYvo
s7vrIHtmSNDrERFdyATSP3h4skYKqRs2hJJQQnpGZ/DC6Fag2ridf/CW76N7MaJy
KoZedzK2EV1g2AgD5DEAcdFhl/N/W14zawMDDe8lRaEuNwaR2fXRDITXJ1sUQco2
xbavcMFvQadbpT5lpWYLAJIVy75OUlXJAFSU5/jH530bqW58uKcYhR6wT6+hIAc6
Bv05UOJyt2Ov/njmHqql9PrphjCwRddT6/nYrND902S5wqBSfQQ9Vb/piwzec5sU
JbCO5PFpnYufUztcQxDNna6T+GQIBkQVB3FvHHC3PdFhecRJHWEI3bbj8P+q6LTi
n/9Lj1Aq/9cnQWPHlX4DVObHFMHQgwoRttJXGIsvVLq//DsMFvNqYZV9rkcxTTpi
VlNwXhTBaf0YTzkmrmL59RZeldk01SXSeY4cYRb5WOy8qyW6QfUJqMfNCzr41RPp
o8qe7X8mRJiDPoWSaoeWkEljQPID2TTRgAHoxQl01S3eA3VnMGRNxBUKzakIONU+
/+CXQ+rD3XV/380X0ZIfYGrnwLfN8B1OoBWSEz+yki/93Yt7+U9Krw9T3koQ2YKZ
TnXytPSoblXqgpWDB/1K4GsXk2BWzJ5fPEBlIWbEeXOwlsMyTcK1op9zRg2dSqVy
yL7YxFmxmdzHVgsD0aj62ueDl5FtqSxk5UgZj6jO9VibYFdFID15KCT+EfwIaDTv
fIxfCx22lXV8BzRL/UrJR1G8vkggeKv3R9aCvFcUD77UZuG8x7pAbZjfR+WUBHXj
fFVzUjenOtW130vSXXivWZ9sbFtofL6YJghSffEQXESz/U7dhN+2XS/MCeD2s52X
1YAWNxjqrKSd3Uy8/E9IH0moH/70X/5LjoIvCtlL9rTi7eKmUbluyYeuYhQxAQMG
79mCdzdxzgqvNe5ROtwzEl7bmGSsaJzNgzEr+tXAXXhq0dUgalNsYB5PKkeCJ0F+
k7p7CAojWWiWBCgV2bVBpOM3bikGFVWZt7MVr7PSbPhobP+bmJ/LpsD21coERMyI
XxhVgNdvcAD2G/7jKW7rRlV7LdxWdntQIfK/jfV43+v7jgcIIXsxhRycSuRkvZT/
PUGlnP5135mwHtplNkuV3nWjacHdbTJSWw+IPG2EjCyh6ZMJZRXwy08l7jpvPzA4
4arxScCuZkA3e7BGiBTdIEg81hd4vkvieR9rIDl9s3fnOb+m8Zumw9+FPBNG5lDw
J0x4N4AyjsJ8LfHpzB9b9Lm0eZEdLHL8wliup//frnE6Mn6ms9jlpnBRPh87tDeR
1Ddz6IRl9DC2GMeYW/0STtAX8MOx3McqvOK1qZWayK1pRwFVNCchXSyeb1Oi2xvO
9VVYUdDJurc+t7ELmNp5r/f1Hb8vkI8RZz3WZbDXf/Mse8WFTPwzSWFQHdZTby91
KE1GKS5APUVxNnCFrJGm60ygR64Pra+77MYiTotXPHlsqMaXoUhmW9j5Pp583w3y
3kOYuQQ4pP9d70ZLEXT66eBkWI3nFDs88QPeRfTWnWubp1NwQfXMXf2RPufPnKPj
BsgGkg9IqNVAMmY2UgYmoywwme1+chs1wtQRHcn7c08zudpHz/zvoQ12p2HW6smq
Gngn6z4rVJ0ukd765/Q0Z0HRTQkoYb0oFF6HAZ70CYRLjXheUKiXs51hIh4UUnPU
hvpfP78bX2m5RK93Dfag2aItWt1eenat9IAaCCbD7VhijbUFAZisInHX/B9rYSCo
EoiVIOg9RdWNgOsmZjs5Ka2Uu2Gow+MTvM7EzLZ34upnoMkoQn8oaW26DHV2cCie
3hJjOOOCAp4I8/e5COpXvCvWh7rHbcRiK/JQH0zkhK+o7kZVg3ujGGhRrzRkDeQ8
O4iqdRQpZLkX/jgVk+kGj3HQhilu2IVuu0LvGC8Vyuv6fj13ZzO42GgXbs78J64e
fEAO7tH2Md4omldnTN82F0kfZHYG5DpLBn641ZlJrObuOUuPsx4PD1YX3pR8I6WM
gzbKQrWQbbm00ZqPNTxXuz75UaXyMCGKgI8h7XsO1pBUcMgar0Syid8mHIjJY5I2
HPvvqcvKpkEqruVfu3ABe2sz2Uv/tjV211a97q2f0yhmOqlxf6eQiHcV0EjwMnIX
yIlQsqmGVKvwRoLkMhztRlCE2ITh5FORFYg1tHVJgA8Ok5UhgzmamTR/9axsycT1
btcLHoTwSQxYiVKwvF13OmbTUfpdWfx7M+9zn3NU5QTGkW2fnifIt6+DWRSe6bJp
mS5iAHJJrPGS5hLY+JmeWC3L4Cd77T2iTD/tFTHb+U/QyeHaeDiF/vi6Y7DNkNfU
rc4u15ZMR0/VLtBu4wsVY5OnCYRxu4Mxr1Ne9qu2oV9l0woTvrIL8Jyzz0h+2tNq
lIkY96XBwFFX+iHFeYTpt0fUmvSj8hp8G1bsHT8Brj7Mc8OuiRkKV3ADpy27Ho90
IW92AtuIrekn07CDCnVzivXT++KzFMmAgZNV92mCzmvVgW13EplXxgOhreQbA5Wu
sTLxH9MzmDbpvERnetfT3/fHgKdA+3ZorZ+yZS2gAXHLc7Q1CYQCQMsCTFQrY/jM
903/5Zvi8v8L21f3mBL88KFYRqOUGKMiTMiobyTsj2m7cuFGMCNx1WDju0sQkKlv
XpH/Uly6eyrfeVu+6jCylbFaVJS0QfJYzpzRJm3pDs6lijsZby1e0lAqf2RlaLiQ
4248lkVwb+QyziSekwprOnDjssjTWPDnQs1yVRYAPjbPJkWjvkPGT59KZR56WjFL
PD/m7LQ2bJpvJvFeLM8Fmxi65h43dM1XI5tTRwFXSxeI+sd7g/Rep5tss0c5YZRS
TjzA2TSO3oBBBcyXhJcbf0ke9I0ObA8SafqCXGMBi1Yww5Nqa/cbc0HTr5PlLSxX
prz3kxpB0AzufEUNCIydjcghdngRI7cYiGKxz9vdOj2q8HIWb+L9+QwlYBlb2A2X
WAzEBB+EJtF8ow7gOxlwpxz7xAyUMOsV62xflz5AnnYrmDqD6LRRoseikgbUmT/2
U3VmB3tU8Fc8bLskKCVn5gZi1xL83jRxIwY4gDaCaCbeqVJu7su2geq65iYMo+8x
1FtibsWlZ1Zs5WCujZNVjfaAnENJG3xAxpEvXcecQsMwbkHpxGumJf9TVNkcKPvR
VI2r/AnjmAC/73bKzwzT5SuGLjqjPyoMTv4zn/btEAvnlOCIEs37gJajuVnOdmi9
xjrvsSYwDjobkyc9qJEEyvoC/qmD+QQkvXWAsL29hl0AfUJxt3qxei+lwCpUlj2q
NnPbmVWuvzch3FoEe/gI8AO5GeCa/yNlYjB/1uPynbOt/K2ALY74yvKuTkIQUcmX
6egW3DvYWM/5ezwCIgbMJRQJhBO5lsfb/XL8obL4WKQBguyieHt2IswVOQTSEHPs
+CY7ZSw5857ljYvyFNY4IbDyMhEyWj2XTzKf9p+SD+y88L1KHUM+wzO8k7im9QjM
EkPqHnAVLPXhGa7FRliNvwDggFNw7eLEuwrn9YcyQbuH2MyqOCuwRCMJcNA7bt+q
NTbLWLtVchliKILDvqOdQm6n+Pov7ERnxcwkJUnDpiDdKXWWkTYHaNUW3y8OdyP4
MlwliFrDO0CNhbTIplkS689FAoBQGXMB6lerfTjftjoLNwhYOP0lNFUwoFUjB4bk
dNjiibbxMcCliW9JUmXA2v80lRlluw2YGPXBf/xJMrd/QHkIWJbR/5p9L7C+n7tB
wcOw2Ywr5+eXA/RI+pLzRtUI+U7oNOyjaxvlljqcrJRYfP0pDhAI7/fUU6jrqsuc
0PKbLGl41nqoKj+3oOlyCt9+ukVpz31ideEkFzPlYXCzJDIn4yf2OyoRIX4SWa+t
NgYOz2X9jVAs3A8TzhrHhWhLh/7f6eeDSgBKZX246eRkVPH8Bd0HHeQORQ+uh88W
6p0CY/KAnaB1aXak5x1syc8jj93VzOJkjmLHiGfmFIPqBzxn1IpQXcE7lbLs+xK2
Ilm9U6UP2EkSsLK5YkKcMVqTvZMKjUUJJ97FYYLGyuJazTMqD+xE1hhvMzP+BSVR
6k4ZSXneCupTuLZGyk0xpeklFNzVtOkQm1VlThX30rQSoKrjH0gDZbbVihJWltFR
DMMr+zuP8panSQUcqi9qK9qDwizxXkFVuo3vHDjD1YXL5s7hUHjaS+IWgZnFxJrZ
4oal08Z/8+OfdKlt2MpqV+3ET9E3o959gJ4iHIWa3glCBDo9mXqrcemJ62YvrIkd
ryu7kjWqYpKzbJ9hpWnWsUYFk20VUoTB1V8uiOene+dDdiItw2+nvamCG3udhSWj
/7Ps7EBxLKh4se4a8L1vsvnTa30Blu/H3ixBjyYAU1y0mOoKmFZ36ogpp2CIEI8V
fpWB2q6JTa5VHSSXhzKP/lShjkDV2dcZsp7vVbid7xg7YXFHdvziDbF/uJY/bfoW
FJj++mAajQV+5EkzrIUrjoVFXvaeqNjOVKMZXnrZEZKn0Y32AsOENFx4GChsVWvV
EqOI5YejIeKvtRQO+Aum9DoROi/Px3L1jkq0h37XB2vBoQwi0V9CNzQLYj2hKOm/
CxmYPNQYPAo8Uh5pKCuoYQSKxGBVK/VB/CNhjUESpbeSLDvNwLM1zxJNWEuv6jCI
G/Kc6TzwKCNKTRV30pddzPj4ZOqU6GAta7jWkpVOBS9a9hK4Xz4rswnrhPHJbzNi
ekmJs9gZje/1JjbzaJ4zG0ioJwI8iLYV7QtB6FBYug73m51DNAUWaGsF/iZe1bot
rSdx67Dz3oOXYNnhbfpnpsqwCZtNHXWkex+JXVeCNCC8fCcN+DSx2v17mK29GyYW
MpD6YV51nO6WANGwpIX3RdSaw+qmVMfwR++C5dGUa0uuTW0BJAxzwhRbrHBoAwJ3
vmLFU8i9/lI20KmGeKaNa168laiBuLDG54WBPMwOeCBfpZgnmdQnDBtEbUsHvpYB
B47tB9Vz21QqHAkUEvLoehJqyyCc+CkT51fPSr/K0YPiZ89fkEv6160P9o4bWoIa
HuoCK3roM/upHrqR/rsDd6OlEE0CdTJkce2bJ0WGBO9E5uDNnRoTLBCQPCYWh87F
OBdVLaTIyymlWMvGeTq6y4C36/5Lj5vyYR81UBJZj9WNqoy3n82LzkCEBYolVWGc
kzW8oOgV7r8sTCB9ZbYlABVKLs8QyUTYW7Mi3FqyMoXCWpMiC74pJHZXUYKDf/J4
SOqTTIRKiFDqHSlwTxE+tEDYABUD9bJycyAKkkPCGFsa3oruXZ7AJyFIv2A9sQMf
ukLwYCynjPKUDMVksVqnugAa06dqTAo96WniIRaNG6ctWc04P1D0fp9BVvlukQt3
36BJrHYgvLVGmbIytOlaf+k2TvaS6uHoShO1CAdbkPhz2Z8IGv6bpTYl3mPZGc49
IH17egRODvH1z9409VgspIwpErLt0q5MwvAwuFTWF8Ihseh4zQpZTjm5hkeXYauZ
lhZyCcQVMTt2x4Uwx38jwwLjwvAwWYq3OQqxpBN4xpL0wHL9D29uR3Qzxfbi+5Mr
DRkUcgoImAJvggoRzXKuPLQK9qNaPiYEmT5AWpn2K2FhFuySgD+FXh738TfJEv6p
38ycmPu/4Gkm+Pj1P79mivmsL72KjHScwtlFt5dBfEoCNmHEYt+5EPzl8pQN10fu
suqSMb8cHSQM4zW91aYhSXR+prLB13/XJ8XRy6Lizz+xSkd/rKoy0IVEYetPgpst
XANjqX6sEt2iyIgddvgFV/THvknmbgi0MWw8Yz1+zdyuCUQGj8zwtrq1kG1EBYWI
NBypHadTWkli+ngMBxaoIa/zZTtxv3hYIeeNRH5YjALBxxvlxXB+NEQ262AfwkTE
0lp/FpImKb/wwYK35f88sLKR0i/+dveNMmobIqkFbVoU34a6C8jmwDeDhfX6sFiv
NWFnO67Aayk65Qz/eIKrWWyRrLSvYslmpqPFOmFSNWghSjyTrZ4A7q+HQQt1nM5t
4Xe4LFBmsRGaBFlfLh5yLZE9k6crs5/rIwuF2C6UbSdFNSXHV8CFm5psWWQt9ANI
VCvMl4r2gfbd51Nn0+41SHA8CzJrTH68WhGTbJK4l+z7bNwqKzyeVuR/kBGdI3fV
lI9YZFBTfMawBzknLk6xpGlx4muYwG9Y/N8msEqN4DR9DO+x0SHhwA1g8LXxgmrm
unl1yPOm2AXNF37NIYCrZePHOf5Cb7/hPb4MGKv5JT/ENwhbdNHCfEduZSiMf436
CMtFTp5rWvsCE+V4+APqUlaj/5CVseCQ/jsRE7mK+bvfQeewiD6dBNwj2qiNdqAi
SGfaE/bF+6Qa5LmdLSIpqdNJ7ReBJKUhmjuWJ9T0fPfxm1GLZWX72LhORczlzJOO
lKz+5/EOhhAWMZVTnUwGvkLtkuId3KryI0O4BL71BbjF3hR+0SQGVMpqn+PCZ46Z
NiU5BkaH+yUAjc+nX4c1EAuHmmO8ygIv75fTtNtsETs+p5GvDtt4N34CCLChsynX
bV6+LkGC/l9Nise0qGt9l8KbtplLlbGNROA0xnuQlJLVf6md/FVkPWZmEzMDlzH9
6KK5iApBiSGet9jFTCfO/9F+j6zTzQhkHUaEAY2l+kIG0EI9oqUGc7+864h4nFJn
szwYLtvbZDKudlrJiCxUfmJL0eB2vgVQE/UEqj236vYLVZsX3eeuXSlh3LDTcgRZ
mNoPn5FlNE++UlhSqRu/ZGkeGakZ7+NHrTuzXG7vngNw0dnANy2TecUHoETfHWDS
bPJglWncoofWzkWMvaQKpK0dthxKRCP+1bjIIuDRLW968CLfSayCrukJWmbxhC2z
/gD2XxKRkZlPbgQKrUaJdQfwCq11lvK2bOjGhFNKUvSRh0yLcrMVerIjnJimZBPt
04OCrWjNVxk8RyJF9XuXB5M56Niy/vFxrWASzRKelgMzyj0WF0hA8pwJ45A7IX7k
lf21MqPq75RAVVfOc83v/AhNdgnEN1KXd5DXqLxMKZFmdOeAqlhDZyGbsqayzwEf
hWcrfj+M4j9OnTsztyZ6FGfmwcfAH7jHIkD0dZpoBn1aO/Yh1lOwPjGy1zCx+U3T
0eJBvVlG/d4vAbEi3mIuq4yxaW5S2sIhMeyNmVrSL9dp62A7CPrctlaTywCoiDWc
xanUGFMdiHRiwDAe6TYtktqCqgMDtp2HPmNEragPBC221rVJ17cPLZGZ42wxOwr0
XhYCnuSKruipNNnKV1iOt0esrBI+kGxi56P2da2FJeBCrlia0CZeZTnusTJ/HdhA
mvShIvSlw0MGZm7S0jubCQzuX6AZn+ipNy0UOpRbazIvx26C8CmV8IIkxCbN/2xB
LONakUp2C2frLs77Z9CW2RwE8PNWx12vLEcwKX6k7vq37Q6Kkz3Td2SEzvD89GkL
VgU5V1ibIIapulv3NV5v2LRFjxgdfDlCXuv4zABOL7hXduEzQX2Tht4DwTmr3FW7
wkfSZgQA5ufILyOtoCs6zWqM+4rOY9JhKx0odbtaqLpY+E0WnI0n6C5eO4ny0/n/
9a7cht8JzdjpBmNVZ+3O94bAksOK+O6sroCrdz5HAEi40kSjQmrlrlxyc0U1nK0W
nhMZ6gdBHTLmgm/Z+dLqrR37H0tOfEGC71KKFNon/aNqVM+b+LU6sXxFQ818nA5r
am1CwSyoxY4I3OVTa252yvVT8q481PHwo95vmDnI/sNx0oL7OXFC0xaMK/AFGdR3
ATvBfRNhPmgQHmVCjNgXYkW1c1hUCNT+rdZk8j2ul5gKMJuo6/JHoJ2DbJDlEZn5
WflkKmHKy4OSnwrxd4Wdo27/W2deOgcaWAiDwh6/kfbzgNwM16A8eKXyQCDoviBO
c8lLVdeouvD1jHCFFR9SrpOsox6M5p63HMRZcCayqEWtcUp2VUpOgZY8h5alHbnf
6t8dOgClkoiyl58x8tTr8DFqN5ixJ83rks2kvqLN+R/plcRdo5Ia4Slawehlhy7G
pXFrS3G0YQcFjAmwTslF8IjDO4/YM2v7kYZnMXTCUw6H11pTK0YYPmjkPBNMnGOh
kGLxvRg9Mx6icZHUDt0rqxjQ3zApkUdauwpdm+KGcyiu6IyOhjx01S0TflkXGP4C
DB0h/I6pQWK8HVIFodE3yr99VYLcNE33WPJqwknH0+UFXuPtBwrCZ6aJhL0qShAR
EBSf9zoRGXQFvUadDn4n0yajRu+ttvqsQQOQRGGPY2cIcjp0I0PuDrtXFSP4PEVU
/i/EQwOOgBqxMrbvRGO0ecXP3kAkmngDKrng2inL7Wm1qjh+oftFxmtiviu4NDqs
YdrnyAlxHQQkuJri9r9RHBTN6ep4HRgJfYKHKRD/C1KyxKvf+0aw8Z49Hc4IGFje
0gA1hp2DOQTHIFl6CReCb5HSsnWxb/VipjJUns6n5l+RZgwgOV2swiIGser6xkpI
7CdgeZEEyNJ9llkAMgZxqgq031Q/RISOvkCiUlwC4kUSy9xZxEa08fEvNpXdflyl
OoBcycisyFYMOpf7HBY2imsgG+A8hgaPhUR+TkDNNGDeEUUt44RbC2Y7CHTz7UjA
NeRbmZJ2mFeh/4FgZN75DOKH4C9kyJW1kVvSws4vvLpSPYMMf3D+4+urQUklvquN
HAU9drL6o4rzal87nEuNuw0Yj38MVKQ0YmxqKCyWT9MEarqrcAvOI9STBdKhusVQ
kBAiWw1pFw6ddERhSauW6H7jIC5kH9vhVJleUoO+1JjqlWpUgBSZq8gcBTe2C9Pb
T4ZDYgm8fPKuyDCU2RoEUCIkaWUK1qF7yMWieCM7KireaQhGAn8stsz3Bs/QqdV7
S73wUxXl2eRP1mhavDGVIfVc3RKJ4PjJMgplxBNkE5v0VEg4xUK0hei/DLuD1tST
ONASFgE0WUSJf8ayVIjmS067VO8CmJIiye1ylfzjpnaW9i1LOzLNKx4PZfEPw4MF
5nCiEICw3eAqPfyff6xNtJQrj73QpzYZGG9ok3frnhfemDATmqQlUIbCjZr9DmN+
+Amt0O6+7yCstrxLqwBi9WirUksvJvHlIFay32ORFmNNIzhSaMudqrYxlYv5lLx6
uOTbLXU0HoMKcn/PQINyuNOeAn2uZpmTAN2bE1amq3aicmcSlBesJ3MBqJ1AQJ16
aZNwCWPr8lpM5WcOAex7wFpXZlUnc3LjeqqJI0DhBm7IBC4l3QXNeikTR7/THqgS
b0ppP8fcQl0bIdsqv+RK4BiRsfojJBDkXdmWxqb6GWI6vx9byZtQsqqcOkAUU0KH
fIugk+pfRy+SWwWVl5AcUyqf6AR42WqEg7UNBDr6EkR4vTvXAOmbSvj2jTXkTXtX
/+GKrRyh4YQjfVn19TJMNHpRRDaA1+1LE7YLQSLUnBNNx+jkJ/yZRwoSvvV6WoBQ
qnzXl6TR/ME4W/S/aW8iG90B7ATTsP6xVjbLl8oNKYxxs2da7S2dpk+0Rp3qXXQu
phs2uNZtJrZWUBz9DzA/cvZtG4DuvhapbtPv/S1MVTD/ryAl/I7BJRiq0Tyb2wPo
qgEA8WC2sfxLZMpw04A/sBkJS1VcVWN+zIEqULsLWpjGlt38PhjjCoAkdpgRd0ef
p4j34b6Qsyaw/mMOEFEA0SgjLkpJCH5pO5gCLTo8D6eJ5b24t/V+LelDPEjAd6Bd
QtDr3/Kd8ImXNL1jNrnDknGUtU4nPuwH3OFSMEPFEhwrE5WFHDeRNdBulynZ+/yU
P9joDIJzn1SbUtgcaUoQ6/R7HQTdw37BN+BJlndoTxWpADJD/9XvRzdBaGIc1yQr
aFg42h0mHuvCjhFmTrUZvWcf9nxJSOu2SymNHF4OQFu1Xaam8p0o4h0y5D0NHLZJ
GNdjwM3tVhcY7ivIytqxHomb/war2dxNOfCz7fm/fWqT8/K0roiwdaSn3OyxbEJp
fDSshpP4jyK3evhf0S0qeIG4XHCkfMlCBhebxtDJjQDXqrtn5ykdX6d5+WxrXs7V
Q0q9OhV8JlAiLD45AFP85PZmXubFCQ8PEqxaEjIqiUQejq9X3PPYfx5jBunuMlIR
v/7a3A8WdvJzKOICeyxd3q4yUgu5WQui8Y/C9do8OxT8N7c8pIC/2VXVJmBvE17v
s+wHmCmT1kqS1PA/qub4S06+iX53TH10ndGuKJIM6zmq7Si1Y3VLYsQeZrOkBRmd
RR5+8iNX1vqWzU1M0DihiHF03H2Usy0jcLjBLcAUbNftmAE+sfAFDqiz9f8PMRsM
dpahRSiq9SdDcLShHsssUbL+YKdQHa++D5BA+Q1NTQGwQoGK+03hJtbMA1BJg8B8
dVWunZCj5wio0UUOREB564YhYUoFfayzsCXzgwyzsHxihJV8SZvYikyn46lRZ3Qr
fxDJkq03xJD5ZiU2R/d++kMWlE392haj1PDBqCjrWFFoN9ful0US+NAIwAwP1yQE
YvwlA2VoASlDTo8h+F/VYqV+U9hg84gfCisdmCURlIvoA/e6Fikc9nCOhpymWJe6
D9kRiGjEHmt66ltttMykGQuAGdtBBDaWgJU5R/oYVxl9EtCEWiuyhhw9Xd4D0M7O
B1ndbnoxKMys33PXRdWdOTZltx7m7rh1iZolHbk879eOVcMeX8O8hrZZeRvfDtQ6
iOmZjobXRlPcAFkgn2Q4Po4sJ5neycfCgc1iQwJvGoiWJSpoRr6CI1fT/Qjqy3t+
dhRXU8xngXNPxF09y+FCAWmsMum5c/0ITWNRsIVEoN36hvVpJU7R/5V96U853/t2
9sFEU8yTCBkAIWlEpj+wO+o6D62vQRNcLz1sJFk5sX/ssFpyXpfVrqGc0H1IFrr5
wWmVu01F5xMNM9Iw+ZX8K/jtKM0HidQa8oUWGNKo0BZecZcvhIDdXpfWletupIjh
rvfyUQhrC3b+6R7kX8Et0BDiBrm4QdU0FcHK/DVkAAaLkMOBo++UB79OHi8Kwb0q
nOyTM2V8/1os2SSJabW3PNzF5ZOKUCcOd8d3gYV2sxj45/uqYV/VgxEtxPIgM7fi
hAbjKctMs3E6tVPdp/dShrS+trUcYvDoO7nsTliPHXB3ed9X4uWx94webpU+Wzsv
1uG2Yk2ICUfoTh+QEhKTuFzkOuaqbA1M/hCeU16fcrqgFY2D4sitPeqBrMAIJojz
ohXDL9l7waY6IIxCjGgUX/uqHWUo5uAEjBgiT23cHwR1+jNhTpOT2+jT1ZQFcTvJ
MxIAoDsbm+ByUe6jFCztcflFR7ES3TT10ymCZgwtlpPTwSOjRROfKugHLEvQ6lZq
uirqOZASJOayxsf/jgQJ+d+9vjMNkCLUc1n/IxlidyI4GOhKoYQhhyRXcCv7Xxsz
C7mmE+fPvZ5DFZSq5qqu5//A4HF6xZLaXg7ejuXkkqtEKvQ3dvJj2R7ZHXhkcYTK
sVnIRRMXGvgmgQZpuRyA4VZua+sGnPOXxsD92gmNCEpVYi6VGWacHxMi/DIEVpa8
8TQXfLawc8zWlLHeXRVv5arJRzgV2+ETi6yY7ojstsGZBLxb3TuF4xrzx28GTT70
2n7+S8QFpqF9cdm5p9LM8ZkDBJrRcY58ckK3ogm5E2yz935l8IrOgLH4TNAgiPT2
SSgGCJi5lfPQmPXwyuO7itUjqUshpDrD9wYX9KwniUasFI3lvswvDamH290HESik
UsxrQKcjrdsSBkvpa3/4+FgUI7ip/pdbX/lCbhUhxPAWHqC31cUR+CNhlOnPwZWu
HNe6iEwNu3UzOQ6EIzpfJv6133AIiztL6/YxJ6Gn3PPWc7ppUVeXxL9XbDO6y6vB
ndvKm62rVYucfVVWFecE6XcjSK33twjgCUueoVzqOYo0oavVfYY+mxEoEHgygW6b
3slhnw7LBZA0T515cqv2EzX+/ZiepnTRsnC/GAhWYG5bJgv3VUhuCmYZlZ2LaK6H
XQ9/rgxhOj5yNfTtrUS0hX22fq70/SxcTonZ3bXDJMn3Erj6PyoeWmMtNIC8Lm9r
xyWGpNzA3U8KoG/o9BfSG7Zqs43tFPwDMXqN3rejIahy1HKlxicBRZGT1fZyxDyH
zG3dmZm3UGXC+D6MKPxfvx1O6pknHiyLVInKkPGQ1pj6RneeVYBqsf664GD9vu/B
43C/2oUyKQUsH/KqRe7yucmrrRnII4Zqu5cxTI8jES+X3ZMgztRyg+mVoPUVtTLl
HAK+3BQA4stnwK89xx3m96F2klFrVyrfEb8nwZ1t78rWiM/F7VvTox4H5eHr6b36
uBhHUgg/VqV6lxsF1aWcAezFBNXs5QpRfuPjoCCMPSv24KHMRvD9WC2WknHn6KpM
f4TgdHjvQYcudLED+kZN4wRz02BJ2oGhLn8tW1HFon2NY05TSDDbrkmAab03B4th
1JpuUcfRYgjPj04zrqBSIxALXLvXKusKHIP8bHThPKJ4vk5/NZUq0FwpLXY4CvhG
okeZrR9vXLykKCqp81U9BH70BTM/jPkr2uz7KM/FcWTDap1U+IGbHdL+EF9Y9MDI
84Ct9epPOHQKKlHn5Anp0sEkUlB/k32dtKizmyIGgsYd5tpz32WnIPPJGRgJEmKT
KNBLhsuu8hpHZCKvyZ6olt6W68D0Z365XEWettSjt+gy7GoKnCpuK6+cWYNJTyGt
BW1p4wxtogLHrfB1DmcZZvlk64tT51wcCRcl8DRifBDDM9DZM50cFyN77vJyJjwT
X82iibTE7vRQvb7aXZuDK15Mvzc/qsMxa22FuztL0xYQM4Q3h44yGd5cGGsK4HSA
+/XKGgmFahVxtuND6+U6CbjTnnpGxpP7fF7VZp9VPMjcDOWBBhtk+6fK3F29buKk
piN65Vvs+xwiqzqGUaZu1vafZ8Yh7bulyV178XiTb8Mr/9HakkUjSsHqaQtb3i36
Lu4GgRcemA3F4NsFUTme5sm5UqRk5RxywyNCVjxpxosSG7ZmUDQR2MajxoA+QSpV
b1ezr9LhgBH1k6YJ+k2RR+x6Uz6S1K/3L4zdErl2ZgpukCzgUHdyCVXGjhueoEc5
YvTJU2kZcb/kRLuRZ1Q8/4DKm0OdLp0Twp+PK/4f368ZJxT/ZUByl5lWsYRR4Yqg
NDDtWITTglwdr1Mnjc5vNQWl1QKqExzxWSGsqQ92dMVul8kGQGqaSqJOppeRU1ln
g9N177I/ZqJV5o2/P67afrHLukSsa76ODw4y+UBmwa5KmhiCiDhy0sknHxGDh5eY
Hky3LiZuyCpx9FIvmJxop78iLpHo2JTElvwTboSpJTol+vS1cR393G0GU4j8SWKE
M3169Ram2NHdvGJgCCGo08zwzvxFGzpGX+axIzVNEFkk9O/rVsZPgTUxz54bQhKN
5AW2IP9Zr10dTYhrNFAM5JoMWQa88PMjImtBbB+4uh2M3ZeVj0j40uvyjEgqWJIv
Yft79DbpFnnHO/iNVrHdZ7V1KKduU2T6+aB+TdqvS9oF2DO0ybizjZszo6zK847M
vwb3w5sg2GblOTpc0O5hjceIT0pZ+Auz1IvzQpY1Nq7sdLbarkThKZ7G5w5dDFwr
MtR+wVVRTxhrRTyYMyTuFqhAlg1EO3Kxes9REEIlQdgVUsSSvtxo1wQaDc9vvylE
LJAHopKf7Fq/qFh//c+Unjo3m4W+63TsoRTH8WWQr3WE0SCeq5TP+RPUs8t5SA+W
U64OyyYcMPJTM+Se9eET1d0+wMGrWk7c3EIIcanRzhJv8/K3mTV9E6+S95bT8v5F
NkBJDmi6aZqXTiLquIWmJSRZ5Tsy7ZcJ1PZSXJxK6fxzXBio3/oOf2wVKDiIeQF9
bR9+MnLSsKjMKrKNE5lVn5VUI7ZljVxCgilrpNZ+7wsqph5wlTLR9kpj3GHRQvkt
+CR12Z4dmq3iQjXG3PJ/E/fYKtqCrf2WJ3zqo4aYHWbgqSkuDMCpVgCmyiJIXgG6
dFLBAjKokuF4JltpXeUox2GLtulLNQH+I4O/uB2qjTmCmpNoWcm94ugu+aHhceRH
Qh4gKnApesGzIGs9r3Ttci5wL7UbJzHOQ3fIcvdTvGmQlV3XBTAfBZTLr5SREfeH
Gh9sVoAucHksYFXrAoJWF7TjEVGSxnQn6AvtZ3GXmvnZ6VA/wCvCYxkdlUa5O+ME
yCF4njFlPMKP86CgxAPNAnckN1+KDoIc5EkVAdd7u+6Y1pzi0MfRuJ2yjSlLNx9N
otyV/aYu+9KpDrXswPNoaHVMkz4tZdf9t8MRIep1VPjbzH5OYwJjlgeM2X7qsst1
S0uc3RHsnd83NxSEDkQ0M/pc5U19xuGeL7OugR5ttwd214HaVeVzWHL128g2qi5I
6XgWzgiabNCP6oCDW64YnQJx2VQCXU9Ajj00cfZa0m/7kynN3IxsUw3xQLdUJMPU
wflKHzkdNFYCQTpDPIkpMIH/+/gb7coN7oIiabZxN/w9TWKAAiplsXrR+J8YOnJM
U4yjcaCUABq8yfze0wWs4uGZnj1eqn/bo8KH13xau+wzPpb5zrHa60CGkI0FTxYz
L24vmn2aazUQXuS+SzzMlh8hdRyq0TNjGcIy8k43rlYo+DFHLp1MiV1wdDtBYj01
u3CNAdajZ5lUMz9sEH0npNaMhA4eUZsRq+Wvl3sGA3RhmUUzuC5Hw1ot+KDllcMJ
TKTozRnWqPGRUA+MuKb/xcucq+pyfhg5M+Yex8f2tPO/9U6s1UEbkcxJfdl9a2NS
dh+enQlfueFsdkQj8UNgfJiaCOdDyITVEZ2qb7EUZafz1lVlfXmBdx4mWTNcZdhp
1lAq/NgzsQiVgE/PGaU+FRz32ZknC74t1xSvBWPQLzTac4CD57rVwLh+rw/hZ1j4
zafAP+/9k05fflHkjvu9jyLlYnrROE862bwxqz0ZzQm2E4wPHAsJnPQRyWaTB5aV
CHsVk1ljBZGhYnhq2j3LT4K8+i9C/OIXBSeEl8mNSQ1mYdAP8CV7AcSiGNNRnvC0
rBh5yrD3weS8vgrrrBFH7BraAZXFqOSZvOylPLV7LWyHyW8hJJGeTykydwV2vpvP
4nEoYYWJaRP5US6n0sDMy9IjWyFw6+hkXxzHu2zZJky/hugyaCd5RXT33STFRfCd
8nraO0wC/XA6cOuzHonT2a/kVAGOj4c0y7ALe5F0HkqJoG+gAooDU3NfEXaTlkh3
BibPULCNsQRv7oZxm2Ckm/vBtKFB/LBdL8c3t2LlmNv8TP2Qlp2Vm1ZZXXtWut4a
TdnqINu0rZoQgsZEe3cpGl7rxptF4NbbPv/y/KZhtGSpy/vEPFVE9Vsf9opaRaTM
CfvkZ/msrOzevb6cQTugNdC3Sw8DqfkQbv1PPbHbYGTr/wd0JOOPiMVhoNKUm+XS
x/qvffmfr0an7A+0rRVoppcYHch3pZmz5JGon5+zX3oTazpc0UxJrPHZMckpf05h
dHU0q3PWgyR5VBodkh+WgaqVWlQlhoj374fcTdNKU5m6O4iAwfvEzizPAJM1pLBp
eB6ynnHQxpwYErod/cwLqq94LC4p3vE7k/qYrMIj1ZGPvFvlgtWhJfQKC3Vjjudc
4BLZ2mAviKBxKayT0pTFibMns/ogIVrQCleIS+xlX0HgrtP/rorzruMtZ19bYeWj
Z/YnPnZ2HcsUwibOHQ8kXmRG0/zesrnEuIgDvNnM6w7uPU9DFsfu5fQRQ8bn4Xj7
OTTqqcwMGez0GG6k6jxH8oLwpm5+M5Re9k0z2AymTb2jE4QvZWe5KLDFp5v+7t2V
d6fLnTtxmcKiHA4n9BPGGFMIocnEpX/AtNpKgZobwRuUHjF8KEkl3H/rYkgOndMz
6gDW7ON5TNnjIDXQK1G8te2kos+/Q9zs2bwAWT+7fKS40i8xAGSbN+u0EePUYBhs
ud2/e27Sk9reFcI2o/yAGDqNaQfBuOZSFzVLFWdnb7fIu3dRg3IKHH4YjDR8yRMD
OqdOAqZEpLZ+NQJnJcYxCTTKMc5Wq4KMQVCkNLqiZD8Eu2pd9Pxzii+IMvxFEIsL
OHGmxdxQ7Z1Uv5GwQgfWliHKfqJbqGbn020XxWZojGi84MeudvbmVrE/daxOYJET
pvJR5vWV30CcEj4cU+oxiPDPKnf5NfKpmEDwa6ib4Xfc/plaDUzwNzz9kjWSd0TB
5iqsCVPMR6mApYMUL87rv/zmmjCl+Oc4ycCYFxgwNrKz0wcnax+TvVYe3FndFK4i
DZ201EhhY0L/p9BPHjtXmHNPqW3KSmCRDIu5TK885dXVMCv0NbTKeFS+9ubnijW6
cqbU237a/MMfdBT0a3Pz5ZqN3AjLRS4me5hW+KRHAuXUP3emPscRSW+GEjXWEks1
5Rm1HymqtucaQgKUCMqXClroyCStxh7D7pi8bNaNTKHPYXD6VZxLy/qRlCuqRrF8
ZrFKTeui/fUjieU/54M2+T8atHwm9kM4gKBVMdKjU1moziMFeyPNiRqBhu4dc3oM
A8SzrNfQ6XFMSQfRsdKheE9aVNpAwxVy2iACzqVcKlUOuGbp4I9yjo4S9Q3LzKqO
jCReryo/AgVuBCD25HRhZUaVG2mZv11GhGIGF44ysngSD30zedCT2lnGBj4UOxzl
YpA8hZbh2yQ9cPukC/ls2O+L0kS4+UDGUP03J80MUGw+ziOxmmay95CcffAM9Ji8
NDi8bkbmxSudQQYcXn5sVbBP8eERLu5PvMU4UopiFDoBctpRvPS3xG8xpF/fpN4f
EKK2YyRyD0+/UOEtyiHslPTUc49GJGit3ysMZ77jIbNBI6gFNxVmqbxgqyzaqUnM
vhbApnJcvNgLydBj3W69eSa3xk0IiMPTBbxB+auwTye/FSIKv8iHQbYh9JpW7flF
e/QRsSooOrOm0x1r/ZXBfKf1syMWej6RtPeu0fkUQATU3mG20bz72UpNZ6qAtDf5
e3jt2A0Pf/Sm88XpvR+QUSGIy6xEVDEZfnMyTg4u7MRTVLTRz3CbQDAMCQBEDgTg
b9t4sYbA7uexYd8TjNGnbXATNN+j0XX/xQRACctEttZ7AKRFE7Vll8oW8XVaCX51
NVvXKd4CYVg+qHLWLA3yxPLFzyNiaQ19hGE3Ul8z18BBxUnA8njpN7fnFQgomKOx
o8Sa1xA4y24m9Qy0qW2yDJe7PfSiFsg3scCloVRBeptuIe1NdvpePQBKsGvc80tP
8WmD2AzHJzUWLLyK2bNrjIyOSUo6l58O5tQvai4YVNBY+dNQfyeeWrtBeTv6Ogrx
3LF5M8Ot5Ba0bjjiEDLlcire5svARgAFbQ357JhpQlVDQxHhYvdF7A1SQXB81vzd
F0UycXgedYnlfToyiF57hjxBM4akXQRPeKS1nbu2BTbX6mUriMTQdPQe9p2XJBPY
/id3NbJkW2HsQe5gcD04LS5h8/OsrnUrMNcKscEp9lo+ugZxGeJz/r+WWZ9GEjqY
qky7nAprhJh6IJxBBhmOwcDvi3wdRKzZa/jPd1m41LZqb9nQ69GXW2mwM1SqBWr/
K5JvNO9Xk0TuihMGQ+oWp0CHKWTNOMTpt2xnrp/YZ5hJ3Z6aIUwjutwTLh95hYQm
pE2fqPlPt3KV0iUDAUzNaYjGGItSaI8D++Mg8U37E7RxbcoHKfWL8IHo6hqPEHRI
HjQXgDaujWc6bNSv3r+WLZoDNlH+2Dxdq8a/ftw6bXUyiafKxWBIL3cQS0X6s7Rv
OVAcmPmx/CVyfBYQsCEDAQ9OeNPDGXQAqIEOdUhYDLeJ/fs1qBcxTFmezuv1v4Of
Ck3NvF+teEO8XBUDhNC+EMsLRMwaTlA7zvEXrMHXBDJAeCEVlEZSXdTssm0cciYo
ac1v1raBaITQyE6p7cChS+5nKCxW9lkybGMrq94zgchZmnWfHwlYqQXiA0d85bS0
ruFAuRHMd/LZxr1CdOskX6fmo/fjAQjiKFiFyWRoIFFeYIWWNioGs3vr9soeGAQ9
AiT7j8ykMoiDsc3R4tD0CkT9LMo39P8XT/y7ZxcOj4MxWydGmAJ16wVP/HWiOwD9
ZZvG9whsZd91UuhF0YeCIGktehGgnZitp04GyIpJ0A8M9xwGMtL55a6t/1664USZ
x7lqN+MlDAwv+E6GilZpS3+p3fWrWBEOS4UQsk+7vr/Li1fq2hH6Ze1QxTJPockM
N65BhbVrDXwUXZiBNidgejwYO0Zt9hoPgfIK6+rc/pfjUFMTQ1R61zQgKrxUAVmo
vH12x834lapq3b47EJw0l2th7gErFqL6+nO16EdGlBFqWfxJL2iNdfwp3elLfFcz
htlWMc7vb7nxuvCe8IoDS7TicyO/srD/PV+AjNIuhbI2NB2M+r0zB2sqJUNQbgC4
hUkNaFHyiQAKXdd0WiV3q1HV1xjMFFr0+Gf3/QO+w3bljrVT5J+v4N02+yHFReKu
vSCTR4yz/QErTC4uZn/KvZtjwUJXlvBUZRPJOoG19OMvb5vAienkoHsvldkb2NRU
rXvcww2aU6gmnjTJidQcPuIlC9mexw3krvcclEe/Q6ZkmFGvjBBWU2LNYes1Br95
C68V9TCel0yTX3wui9BFLnhC8wjmH5E7HUi4vGc+QddlwoloCrrdD+qEZYvnVGjj
Nwr7/QedNzmdJPi8Pdek/i0g9zAJJeCp6s4uN8+v1WKlffGUQ509krwkhCKT8wuS
0iZjugZuyxrS/pB7PIau2lnNKUdq8Fjyg5iUx0fOFx5+ge/twa7/pM3QDpGzgEVW
/DONpBGsfWdYP4M0nj0jW1iQ1sMmFrXJEKmFhihrAUCHhTzLoZpnpvhaOixXWylw
1V8MjE0vZIlbYgN7HT61dxxHRYg/dIDbyRjyBcAcQxzwIW1gVVw+oyFVHZp3NK7j
BSMz3Csc8X2AqHBvgrZXNwelp1q6QSCDyTIXRf4WrshMZflwJ0Rm/4xsTuKgz+Kc
X/U3ZXC10KULkNDnLNDMJyXFUofFyel+/WTSSFGzGkj9WxGuBtKqBvBo/302ztCf
9TRqc4rD0WJD70ya+Nc8eg7EFiNeeT8+9654FUBMoNTeuwNqKFnZiUHIWMWmI/hi
JW1MnS+zCi3LImkWOqK28pfeZuUBcg4XSezQqUPT/VDFOR71PQ56rNcVTag5ht4f
5KhxAVLuNzwKjfc+pWXlJjf9iUfw3uGZRJ4zOy2Qn+CUUPZzVVuWJNj75va5QuXR
SYV2EzGGpte2HlQbXSLK7t89FQd3uxz9B/wQfbAZSykNA/Y5r2rQLxkJQa2wxI3w
ZpdTHa0S02BD9A2vcYK+3JcOGQ9JC5AAXEMM7S9Dp3csS/bATGhYO4NZ4BIaakMR
kyfV6HPI/1rpHg0EiqbhASXSTcJM3l/xMyVGBUEpvWqACOupHDockQ/xD3+0Ph29
xqh8ZOFaHBgrXx0CZcoHR2Hk5hOokNmEHR+LZfgPQ1KDKPFtgaaJnLM1v9S3jYgQ
rkzJUhjjz4WmN4hu4854DkHHV2iM9p/m+DuZ/51bZUuNVGMe383zpyM86paZzaAO
R3K/Y+7KyV7KXgYTnOHGT+YKwP3t1tgiERvoP3IKeWT9JjqtHJwHWzJGSxu5TGmL
NNZO8C/PeL6tr/AEgnU7GlB3OnzbtAAP/vJ5TzVeN3pjHNTBI5cRfkJ9JUlXUl1h
EDSicX/EcxdM5nWTDmg8z7TrR/bgOhn30+zMRQmf0rYZTtCKJYYyRUMoxOs39eyH
1rWf+P1LCP9/AupJikPeprkHCmOubfaZNJPIA9veuqyuzJ5xnuuL64etn6Bzv4al
UHb3lS5B4HbtF3hGmoCegH0yrT1cVE6ogFZyWL7c/6VDJfyzow26AmGzQUJ13FlS
/HzGN9WQqJrQ3TMiyQnNdooBgDy52CoQrFbrF8R5fqSSjmmpttwJoHPL4TqBbOXd
j0eqqqBmJU1eg5zN7iwCaJLidEeKns+Fz+GddFn1xjgT9+SghlyJKJv6LxQNCt7a
coq5QmwLTjJv0hxavDG/C3h8Vq9olqFv2tRJN8tMoexfQp/Ry3h5KLW7Uj40aC7o
CkqYTaVxvgmmkmX1MUZH985e2p8n5jDJLpcHwVvmvm5maUIg7Ws5KNxAru7tbyuH
UjqEVhYUK++h+wDKITSpancsJkWJOvwwSyRl4f4Pz/zQBTSwHOwPcfgFtaMKSPBO
ZCntppi8egNW27T1+w42vczIApesyeATcUbprNuzFsrvcesNUwoXoVovpavKUcqC
EGZWyVXf0TgET+lwQQVuakomnB8VesvX/Q3/Q+2x99BtN6AHhDkBwsu9OVth8NyW
Orh3f444nkKDHg7/t5llQD6lFeX0aLmE5PZd1WVtcB9jalnuqxHF8DcXlCoomg8V
wM/hJg/DMknsEX57OmDj/KHUsm/PgQDSDN8LsW0NycAgZ168bcB93QinP8PLhSEr
2+wB9I9mDbU5JdxqINuvjkRK5cZCCmigef3mGqNhRxn7q0AkqtrDW+hHvSO0CiQ6
6dncAphKCSj0HBccztAUvqhviAiZvAkQpOEUt/BX8QKqtWq8IoH01gxEalEeRnLx
eFuxNgsw/z5AnXmOe3GrZ3jC3KgRZVu7Typ2gNwLhek7079Hxr1en4fn94jWZd/X
n3DmeiGBiulL7PeTjSGikLIb4KzGGadPopbi3wDk6qk93AamdpqmbM901Q7vPl/1
5RyzAQlCGzGZls1EIFzZODOk0Z/MzOMBcetAg3vyjneP67iMKveC8yE3G/xz649I
aDmR2KqhZAzwkHE2cXD3upLHv8uafJyV5h1tTKsYxg5KjxJBx6g999k2qkNOccw7
0HO7g1VsUmfV8uITh2bgvf8n70Au0l1/n0QOHCgXlDXkA/Sp2i0cpxSAJ0/p2y8m
ISqr1kYe2E1LDYCEGb8ttDX6UtdB+hsbcqSSIVFlN3nQpMDS1YQ/RjeLfcEQ1r0q
yxNmkatBPVU6OvZH0Jh04bOC9vWwd7iMoy9qx4ZCBm22KBtR0W46rMpaYGuAJ7ON
IWkAtJb65fGebt5DagEp+Y0lyVk6YJJeB0lZoCxX/hhXEEIU6yBdYQEoH/Dqk9Xm
R4cJnncaXatIRUsR57WGe9xLzyNlsAgwGheRqT+ubRU2Ehtmfc6j3WDBcZahJNBw
sF9wU2SkfsKDwDlSffci577iUvjdoyVtCJId+AdNpsE4K/Wxa54AznGWZ0hn/hdR
mmuLmCUXIujwMVwyQ6b6iUxA8ev9fIAswP1YJ050XLmJCmYeFfsZyOh35BNv9jx0
TZa6wU7oIzNBldjQL2BTb8wtdam0ELlnJUrfGr0PS7WldZVVbfj7CLsExP+bQp/B
A9JhwkPNJCr2T+9gclURMF6kImyo12WLIdMRnGztZEb5+xtdwTnN6ec7PfmkTE83
bFlrlKvSIJAjoDF0xlWIAdkluaeVerX1LRKm0xxubNVvIJRYoDCAqgHv2NYbSMkX
UyXbj5fPpBdoI0mvgVjSQ3dGeR+IFwwCwQh34yaCEm3X0Yt4B+8nEsnKS+4jdfMm
UK9Aot9uDXehML2d/LKUqNIhQRtdYSaxtHIu6Kd/yx/lAlhWo7HdqPpUvuJEnLPs
gtUQ3CPodNSpPvmRrB+lwYPa6JNHUU0RIOQk/FUs0jmJZf64BeHaP8lkLhmFt8QN
2Zz2KGi+R0VYRj+vxmcsVAGWUKl/zBjFLcC6MQZFGgFHcNdRDQWT8mAp8M/nECui
34UqFzy90ThlWgxcGzxG5/nQ+xB3Dg5x2ugfBfmJcxDhxyK/2vvVkcqkulRCsBkY
+AKXtQO8hZjxe9j2yRKJNX3wPbpjxPa9AzfmzKtl3ANZeAA/mGUteRVHT4uD8Qoj
30fencTKSWnmnWU/O6lwpw3gQ3TvJWgQo8c+rRK/jEJBgMkF4u2e+lLD1NMt4EKt
L64LgY39CTGJS0Kjfvr6/dyq+Bttt8ZLD1X9n0pfbIz1gAxzy4vOU4+EO4EMK3LV
zIIHdXeGo8n7DFdWlZgo79fsayEDzhDotpFfu3t4GoPEuQwCjBf9JWmMAmd5nSTs
glJOSGVg1CpM3Ploqb1EGVAdwg4HF59KnqyKDMbtboKS3t6QQOInSUHJCaaB6jI8
7mqzRy1eJClvNHrAeZn/JcLM+dyu1S4LSGLxk+Jd+TKaVlGEXyHikc7XjaHBmqO9
YNbEazpyue8KtlxBkZdnY8Fns+wOHqH/GkV/xP66R1lt2JQJYurWtR7DeYj+wwDJ
ugkg3PaWK/6lJBndiacMOvEmba8vlu3uQZ1IP5yCIX8D+HMtpIDdboiNGOwVwCWb
VNTN+sHXhV4jVSwe29reT6XyRNypYm40CbTPHDkyAbFOj8NbIeBWt8EdZOrlTrao
KO0SK5LAR69zv7BGmLYJgxC1JrC3jF9w2d8qWYzMfTyI2VW+LG1MH/rElNFWVpYQ
kbZd4CMo0GsMUuAGgVS3jE4iMtN/xZw6skqqxvxdujDARUK2JbjLVhqAzKXF6FCt
tNoyPv6X/cRLG13DGB9Y0vHBc6uH35Pvkhh7k45giAnXWpIIkahDQikZ9cwvSdcX
o2uYM7f+tD8oMTLgFxdO/Yk7S3MpHZfk3zmkV4RsB7uJ80abwWLxaNLmnvjaoQzz
MoiR8H5MGrmrbuuIY5NjxHuvkZdEPFaA2qVgWiWl+A0enanHDMTmHYI7qHNNA2uw
IMwMHpIfXpK+N2/4+CYiNMc78OkrVPCb13cXQbd952+RFRmFIoObJnLAR3OFYnrA
eTg6lxhMiXOnDotpcUr8PUncP92Hyah/e0PUpo6P5evJehlYJfH2t7Gtl8T8jLph
lj2nNID8Iyul0/KQ3dkoCTNf03yqLoFAFvLS/o8GXdkdYeEkoB/Tla6cONsYNwfl
gOvE1YUA/7w69LPkPe7VnSuYTOMsA+pjwhqSw4lP/4Fj2Pt1QeuHYcWHj0SARdqZ
Uwam/7t4v39jPwc0bjrDmueOWHVZIMWfjzYxgS3OZ4ssJc8XPDYXSMvxUzhqx4Ug
wPtUYQ29acNVqSa41lCM+0gIf07GpipisIFtxjtzRK1E0Od3DdVurp4cfYUhhMeo
vzJ+YP9JlEClTjOyFs/1OfY1a0PhVzs49bOc1a6zN0pQ1XEwCMdhBNXe0AIaG1yi
5ca3cS2+HJDzBcu64j0ETVmxCYYpjSgdBG0o205cSZ7P/qhwcPxTPUgGi2k+wdRF
BEXxtw0YjN/sokrCjqADVRcxpIBBK4pLaX4kcQe9v/6JHiyTzNMjgFU33+PFqtW+
XWgzDoF5pRJwM1KXn3lQbruXGUQGI4HYvaOt1yWHJVe7s3qROTvTY6tAVtx0l7Mm
D+HOqUR7p0IejQHFAaUoBj/+8/qxEU9JAMM1FBOaEZo16/Z8kQxueE1PL1hm81TE
cF0UqNa/keCpNDzVyvgs55DUynNAGkhmx/SQbegPNsL0nzGiAh+BLKm5tw7NAnpL
HFjrzTGaGwWpUEd/QJ88Nrgr87v1s51h07zFl2HQhoNpPiZj0O5PVU4gmNoa/HZR
+czovaCNvj1Zo7HMhU8VfUHweyDTLSkIlW3oUteRHRAO9KbQuA/1jcLBPVW62a5w
Cr6YYJSuYO07Y9Fpfz1t2HBES3RSaiHhAcRyAAcALWvXq/bm4fMnrErdA8dvxAZh
FiSZqcHk04a63oRxrI1zqm4dMQHajsxJB16+bhCtn6DSPV37kMylw//YPFhVMuaq
r3vpAcKlMkm3Xr1IjuYJ7FfbxLmr+ltkUGUqrwO05DYQDbSkzNv8Z9vW3WYYydP6
/mBqT+L+fZVVMXo2132Wvudxa/Mneyk9z9v2dxGsOUtESbiEEILmFLOQA9E3DrX+
QKJZEMlfgxbUlofxiNLAQizdp3JMFaA1grYi+p9+QGno9GIljxtITEox28/lOIn5
ga9sWDqsZNmOJVVNXMJ03wYLSi1Z5CjMaPX4MT6xjFYfntfC+gEwhbSmut4Zjquh
zqOcoDIVFZ9X70tLw1Zq7aWB31n+bHyhXt1FwlBra4obeHkiWlqWjmWAZO5hHSTM
KvaD2A8QUA/FGso2f5vX8ZmPeYgorKDH8n/uDNAXsOkgA8BReVZiAef2Qwyiqjc/
8HEHN189bBLhea0ZOtJ19v02qK1tFrBl1u+gzWc0eMptE8fTHku/d7zSGKfKPgeO
hCEQQoibMmzQEk12T0gB5wlbuKkIu5rRHSBYckXWqKC73lKaFx7YFIbMkYFX9pBa
zRvndLLXcTJ6yW3xnmnmMuVzpufqFLazYsZrkr7SeETd/B4d9LColT2AOPGRTFx4
43BROZqCboiIG4MliNjtX7nlWfwRotDncBR71HAEt7MtytsrloZCUYYIti9oogKp
CQ2JbeIutpexxIQ53ODCEZ+YRm7KZIhyP52l8dCx5Db2RxoDnBRVkSqgwEarWaSq
/uZCVWaBQD3O6ec/+9ka/bHrEe1NkJPmd1PpLXIoj3bskqrT4CMUaz3IEVVjk7cA
Ehk9pP1k2z7PB3JmqZZoP7o9BU/dgk2bWNekDk4maJzoZKZ5G6fDxOEOamBVKclp
S3KRUBCmYniUVAmTAL8CDpO7FnBEBvv1GB628rBQc/RCEJd9QR8o4EokVkRV+EVS
dGuma2F0w5OEOQ4k/Dn+U9kX60R73UXwfFYyxjImYRktuPxXC9a3hPbe0LQ0OXVj
CtODqAwdCTB8QzzKZ1HWlROruE5JJz60uL86HvC8GvsONGDa1FH4ykunNsFy5QHq
sthsikGaq4+pkjxCfSCUT+3q65OFpZu0939N5jVngn/Cwkj9yrT8ldDgpymvW6eQ
yBUiAt99eKDyqodj5ahfjJWOezJP7BOpk9vr0GwICr19KrOxamGHMJvz8I1GD/Lk
LNGPWDW+tRKZTLFlnNngFxNvfZ9pgvOLhkNTnjIHZU7CIBVI6Qpoh6/EB3oZCINX
i6KxKV+UdEAQgts9BaBtmfLozKg8QGeeGXdKN63Q7N+L+qThRPA++IWCAc9B96SA
LDJBh2Dhv3pdapD75S2Ltr/wnLWv2mVRYA/ybOwAuXNZeBAaHWobui6sJfLRhfmG
FUqIpN00QNsaz09hbfCcAT5r7o1QOBKntTq0hLWeY7gUBi/3/JTYdunfoho41Hx2
8/kD2QvHWJxIRwH+VwJ75kkStXeTdg7Js3j7XQFTKt4yl+uRZWMhfBFeMB41l/Zy
xMiKGl6FE+P5ZbluBR0x0bsIF0NS62INUZy0bs3RtXXfaAoA2QcfpeKRH4mlJLAS
GnA1Bk2vsjlaWwtl+4FP3tahy1QvDWdkFwp4E2e++mJhALjVyYjlocZkeR3o1nwc
f8q3J/oibLJPRrtSfwJNjpz5E8qVpWFSEdeS9MUTmAjvvTgsKBkHUHqhtY93wL44
4xoDNti0jeLoYTE5p+rUGXbY36xGltcBuIC1rjw8g+YZaeGj8u2jI4/LJqI5psE0
rFXSAw7PNgq1+xBPLQrh39tSNtfW+9fZR8Dnd2SG1uLRFaV5Ee7bo80pqb3kOjIk
DMCZtxeR9MK3HTjBOBBkmZ66cefac2qO/Aml/49ytvHpoZoTdfe09gL1s9Bsd8ls
z6RQ+vx5vlJoTTbvQpXSYlt/ZftvFhcSW02BeYlGJht8UJC3VZ8ZK4kUGLN6u9nl
64OOYYv2TePBXyHsqYSTKpDMBgcUDIxgWX1Of3P66PPwW9HeFeYbVcKY6gULx6YU
QRbnEjiuiWFutyrWINk3TpjOz/ux9EdMHJP25Cw0dWYTLq6e6OgSfSDUA4NUI42u
4F/ct+FtNI38gPpuDibcFNT2CRBk/S9MVg1ZkwuTtu8RHGCTHMPyEq/+/f/KRZP0
jZzatDMCS7wp7oBB/LFMRlvVD51pjtYF4uGHrB0LW2ouXatc3+epj/FoNkzXQo93
Nz2gZXjPbVoki3chiq9ZfTxTTtBBqFZUkhINvry/rTkcCdsWZTe6+qbjsZC28qWm
0OFozgdKt8vqhQ3Gq/2fTRio53k1I1UkhZNep0+weKB1Bhp2sfGq8WsbBCHaB1EY
Vbs7m/ivoV7Amr6/8apUVRE6kRkRfcfwa2GNUD/ykovAduBvBTyH6HCH6r8GOC2a
hB7fZaH/pnBcvB4N9YOsi7WASUQMiDZjrjm78q9K8tLNGY8BlOwMQg1H7I+jgdBV
sU/BX/48YDaXkBV6KqIM7y1OkTBChxvbp6LYftNgMMcKo5Z3FRNGT35W8c8jQYVc
L+C6sww1aX/oCvwP3AfjkmPRlh6UEsDOp8pHPxrMr841Pj8TVWCfEfkowy3B58Os
4wE9LCWQ4Eu1Us/X2kU86kH8Q6cEy22pJRSi4od7tsXwjxmb1nDWYo+1NyqnTPmQ
KjwMN0cYzl+K/S75O+zYAooL9q8pSTcKtNunuDudbsl3aSZJx9rD0qh0+ki02FU6
i7Mi3zJ5iHPgkZ2hBoDwyRahXPcXuAe3atp3OKNwFt4lkWPKoHcmUTTM4A5cg3xw
HQdcqtdodSfXdt8LZ4TkddAHgmC9HIA1FuO8mAzIn1HYG+ToB6F3EFcuda44SLOt
3t6XDEVyikyCMvk5m+AursPV8Y7D8QKTiBnaZ1J5oWUuhWKWK3QiB7zKCBOaaulC
33UgpqM6rOCkq2bbExpyGwuVjkAMvFrqKK5pG1+RW6kJx3lhu4zRWg+v/b1Spjgn
xrYZiHODcaC4iPzv5W4ScwctBdPNPvOV7QrN+5YaP5ciDmWmS3qsP7oMhZWB7N1N
U7t5SDgcyhx27oSNChaZrQnzZOOBrM/+hlOjkmx18l3XPwCvH9w+biP6pKCGuyy5
ZOKseHXgyRcNMZPpqMASa6FCh8uoWelVuduyXrqe9o1r0SZWx59l74HSRHlEgI0S
Fl4AC8Aj9qRk1UFtL4SPe1hz226D503ptHq4uP2REABNqxyAlRlMRsVRq14PPZMx
5yxBh3H5MlM4t2/nuAEUWyeU6I7/B3P1xelUq5GLfAUPn4iV23ZHYDA4lOphvNFu
7kvV2QHnn08Bexx2ExujquH1LI4RVidOFxRX7yw9nxoysL+TVA2wbSaQW0YWS6wF
GBvMr0yhsydg7mnUBt0KAYtuQhOHfKT5A2f+cgbImFYVDgnQS5O2aNS6/eWyq2UD
wv6N0lO1ez47wk/VKSKn3/s3ycvOiAyBtdflOf/7/VxTj+L8oblZOweC2MMnDN3+
ZNqQ2N4YOvskbrWNoZGNmM1ZaK+mQqcknhpN/bRP78tmazBQwAfEC0P1uAtkNtte
9bhRc4r1tj9+kveuSs3bI4vA1/eWs8cZFeYpMjUSfwIilHkWTJKBm6pFkG30SdYB
bS8Eva8ztDPR7aNKmoyYaAfrkv8K9lccTJQ+ItbS70ep/HeR3CS1z0Jkxm+tpZgx
0TaWrvvELS/RVJN7PHxNFpk0OGsn/ufbWeqGmNgG2ZOT4e19VW2pcCDM2fzuiUcc
5yA6sQOlBzdVvrkKyyLzzGeSFXe9Ql586Gvd8YX8HN5vROW2sHwmcl39qNYzXZ7x
nGWePj4A0D7+gtXnMJclVVCV40X4vpCRX00rC8UCamC/xp3yQ8W7FaMHFNYMUGxv
ZSpFjaKfI1XiGqWAKsgjNcEn67gVn5OeBWvytw+LLModDYUTeQ6Iyl/AQL0kBI/A
LoWmpMsOrjtzqfL+18ZXU8HIHinmR8zcTjhhoo3pCe6OTj7jpzbb1eHmZ5nPmr9g
f2gaf3MXa3BFjJOaSm8c3QbVXEVhHBVD4j/5sNdMBnIT/ESO9cQ9YZUzGohEYYdN
An4Df4funXfqJY0RPUa1AYCeKkp5frP9ocwh2pZWX25lVhWwqYdtEkpLu3dOGx9/
3/JnRTO7OrUyH2uF8PaOzf/8hweW02vTcNw0PmZx/peZXZ1imfiKBsSXTXbduHc9
U4H4ngAyIeLV/s0kcjq8K04RCbqH2UTWUDW0XPUXDeZxQaQlsH/8GEcXQ1o1+CcS
kN0Ib3KIkGi6b9pxh2nMrKdEUTbHxGa0etKm4Pr7vHZr9MakI01IJ3Ety80cXo6c
LkLtvTa3g2Odbwv2S9GtsAB8C1Pww6TqWO7Ivhh+i+DGLoyikSIhnAo1nmfPGWo6
2aR4P5hVFmNkCHcMBSk/RXoUjXGEK+euR/0HBUoBVBG9ZlYlAbu660gQM0zYxU5a
D8OEOx8Bxi5h9KCItK6xqscKQlKhSf1odculNjjGzawTTb8t0WbEVr3wmgCLidGh
ONePY2U8bI36YebaiGdefwWzPpHNhUMk8tDvEoeUMLtwahHcSPEneeGxrAYeF7uw
9gyYQQhkaAntOkQssRrEmfZBk61LU/eMmfh95qXnwkWx6GejEHzlceYG7C3vunzV
+v3YmgxAuuMXrycJyb/x6YOlNyojCoQsuGk8hAtyTuEptjzIFeYstotdYU56Dm1z
sJayjtV9339AC1wf05pfRX8jaqcfzHe1wGebPPABv/JHfhUrpvZKUJ2k+d4se2+3
Jl9aE8RaRatwBhvBlZpx33LN3dlUrGH1f2zNadesitqDvwCEKab25NiKq/SnnQq0
1zGa6MUcTlmm0QACFEhjSGDQVfB4wKcl/evy8I52VXHhMXf6lamRW/cgXXoV5f/W
wKnwu/PsfQPS/FZ+FaboIrnCuNrjiSjpgRZFjIRxGXYUHvSOgnIrpz81ELKmyRg1
PdTZYrC0GUWUzZiEeajnTAACH7txXt5pqvQkAZQ7RovUGVy+MT6nr7KrM16MVkSg
emYs118Q9IAfrFP3SGy3sPZ6qmdSofdDVe+81CiBraW2RMLVr9YNCfOqOOpSm8jK
Oo0fsMVIiFcVYAoBaDlln4CRDrUea4RlyrTXO+I0YW0jeY7bOrFai7miZvCz8kEk
A1Gt8AzLoVPyU6xvIQUoe2gEAhIr1FvEJBDOqqiijxtN/dHI1TsLCMvuPtSY/nRj
dX/muaX92AQ0dB0jn2UZQVbRvcPtCHELvrz5EgeBgZodiardCh9K8kA0yavKrLDk
LwhPpUj2CTKQgHqxcvWMPiqiJ9u2WXoHtEMwngp91/Fr9SYvE6YfMljw1MvEhEyQ
0bdJaP0K5UWg4p2BILSFypvW3m7d5Aalgp9rOIHgDBa2SifRU4p/F87+vGX0riEf
g61Jmc2YPfDnmFJP4EZ7ts0VOjWKSrWJEfZKIQ7yyrLPEmjfO6+F1jInYXiygUTr
U3ViXmnz5M/8o4STBGNekP/pG4beM2V06vfwuq82JxyB77fnFQ0e3kD+MlRPcwNX
osUdjhCwrD56/kz604i3xBVTThEdNCObbM+ZWJSl6h5XMpA8Qf5PhbI/sBhu46sB
5Tclr5SKx31qx2PJLZUY791qlb7q9NHnACrHznooCbLiZPiHbedS5Fb5xZcNdb7w
SZIsfiRr6cCGiH2kJKoB7zhFatkc7GfvhZtm4cpFT14J2FB5Ypi0pV671h6DsyOo
KnWfiBBPvqUVgFSso7YvMNqhSH59PSQv1OJFCzSldy2zmCuQKCb3xnKVcQYfedL+
1xJv+JSc4eJ31vPpYux0K4dQ6vBY/B8O2/nRtm77NZSYL9HJ0Xvwgxbo8scgHzVN
qIPbWndiYZvx6lwRdTA6Ad/FIOu5VMIU+J+f6DMBgisogrRFKTXwsnetsCPjDfai
9E1iNHOOUYt/Y4pc+1DWj1oJIH28ov3pnNRWNJgZz8zUdaJZLNqLntJwm/uaQB4y
6wLPo860JwcyuhT2JA05Ya4LnQEo5FtScIJPNz6zo2OHKw4nxUvf60tU21oGLwKd
8GT23o+Z8yVUvtQUTpQVTtCCJ74hewVYFGyad+5qF7t0/MKGsrVpHZiqnowJFpNP
tKMvfYYxsG55PkHQ5rgzESzBoEa0B6WmlfdbyYTVVgOWbdBCSvACRHbphf/j5nq0
4N8BXlFxYW+uiFOSW4TEz/AxrLqRnuR9pSa2SM1CrDMyAeaCg0f81kPzEYliCyOT
GrZZKQuXNEirP/ghEaEJeRGg/oOg1V1cYBFhGDvDsMRckiwvkNCXNMGga1iHzrLI
PpbFVBjfCpJAEIXQB1wctrtINFgSEas5f+2oDxibrHCF3Q6AoNeNpw9Fg0vFbhUs
v/kalYeGG4k085fR+1FR+hAQGCh5BmZBuTfVfjDNLJJJ1JggMqGldCkBHfeh5yUi
SyHtW/40wqHDceDvzQBrU0PeQl2Tyx74n524hPOgyrifw/ypt9leEjNTzXP0eMbD
dHlpF7Oin+taxKXIdHNySevbXdcBBrEZlff2DptBwD/T0lAztj2k+6W4J2YlM4/G
X5ZGUEk6zsTzl/h9Z/qU3ll3NMrKI47SZmE/mHWOIUkUwxXuzXl1Iabmlh1Fnpr6
A3fB/0tiWH2lXwKx7unf/z/j5a+o+jpEORiC4DbSo8ghjs/R34TYFArJ9Jg6yzKi
PN39sDH1OBbGK/a4JLxFH6gjob+MdedHm7oMk75LqM8jC3WEPUozYZSKj9Ri7CZI
cW5rRTCxWXNzo/2D66u1oE+78C8Kp3d3J0oN6TioUqioq+kWi10upMDSqAUOb1bS
pdLJ5snVBZtp+UsTi/2OcPzb/8Q67sNdWOly0cr2FEXa5dgYdy9/52mhF15uybu5
lDAZqdzI9lD9sJWBUSM1WMYETui1WuK0A45U6uBBlSGZFHtYeS8BDR1Trjo8Ey07
2UKwe0Xr71ymWwVyqt5R1XzLeCdk2DDCrW054+xfddhHVqehldI5Bt/xskIVI5gz
/8C5lv9GanPGCsOt5FyOvOiDVu4dMUT08ynsXfeNoMxwbHWnr6+9SiDtqlPXTsrL
3UzuLb1yps+D/JaeLJC5r5tg6woJ0971vFDtJMbmpkxHR+1bPcPG/nbAPqi5XWHm
+yv5lO/3zUcUn9cTh+ouXqoK23EYaYlUkbUWirDebosA+I47yJrjfzW/tJrnucA0
9pEYfyueyQhia0xDQ95jxPPAN9Q/L58T792+Op5W9pmcYTeovuQGbTHxvE7N1csR
XrKnjqnB6SmYV7c2b38nCLmqK9VGtzfK1SFfYuq2h3MstQVBY0QjWOsWMnQXZ4bH
/ZRifG8l4LD9jJDvViZCPk+7CV+gACfHM2rAFzkQ0xQ8YIyp5seM1lH8nOesc/3K
bKh0I7s8JDMLO8o2ZS2i8L2MUHzYdt5QiQXERCmmOrAatLOKJjt2Xu8SKO1aebT3
XoY7bKu6zvJjJHbBTuD883jBsO4sfpyawTllfgfss01QfC1Oe4dQHG9rwLa+A+Rq
nrlLwhsUX371mVTykLBRAG7AqsZuUFxn6ExcVqjE4tQpi3B4byJ89f5DbDbq95o/
+wQadY2XAaWvidxmQYchCYRU1mR4jL0ZKxszywa7VPlBute5Aa1MObO3yyHbopmh
3f4tViEoBoNfe5q5RuFLB8LNt+s8TxaREpVqgZ9fGJhqrqjltUYhnjWas/dCyrsu
DI03Ex+ztQWgSADrQvyTNLbiqH14LP4LhOf2DlJfok3GrNQ/S+SK9oJyOWqu/6uQ
PFgfHJUrX3tLGo1kzuSJKEg0bo16h651ubkFDTXIUv27S6d1Tmw1zvIldGjjemIj
AWFrkpmv3wsscPQeqq0ypxixfjw6mZW1/dsRmVGY6bwgRDg3k7SDoSVnxH1y3Lno
h8qLAfat1SbeBuKA/viov7yEwqLbjqB7jNa5HyOihhTdEmpgOcxzZod2hILX37Yk
zRzg+6F5Pls1ZUBFy3LOCr4AUrwBCYCGTT4ZvYmJGKA+RnTj/aF5LXEkQCnbYdRX
1gz07cl/lcrOez2URZ8P9FFrnV3Kcu/8JBDIN3NXqwtlbbjDsbIkAVxJrGcKU/E5
rERdW9YgIMEpQdQajao4janhrMcI52uUbHGkM7kuDCL2pUa3b7FwgC4gxDkVHhNP
qF9GD1HROzy8RKIa6bHhclI7YgbDvRHotFq3EMwNj5eMqgoRoIjsge8mNVKdfhZ/
g+0QQGkaGWsT+jZkaNzcFhM6LVLgAEDRE2eIwA6+X/wu++5ZIHjPzGF+rwg/Ji7C
Z2oCt7iSxS3Ae2+cnrPiyeDtnWXTn8+etmQ7iG+8jNIuercCzdlJhNNR0D7jCdWy
itjjqEJZvVBZI6c56LGflb7Wzgl5LwNKXg2axXb5rBfiVGvFYiTD/dWJhvMu0FfU
GM+RxzXOXKxaSbeNCUfIDUs9XyVlyI660c+MvJy0+U7lN6kZaKUHX1cHpe47uv/J
06kraosqSo40wkLrH9ITNhUmG4D51lVIZoYN0FvYcsHriWU8L44dVIqZDgMCMQf4
cNh6Tm2ABYyCPLbvK1Wt4+rmNwwFTO/wA5742t/HDIFmZZKHSUP2/WugkXWJbTCc
IH4y4kajldv1LDGutz6Tgf60nT8S6FfpupQclh+vmt3f1pSFZpejAPoLSw9NSjIo
+Lm6Umzd6THQWPXshakcxEcnWFVCx0xjqMN4pZTaRkpsJLbGkm6nDfbIr0y4HxHm
GVdO7vs1wbiEbnfIJU/86MjxIRHp9blZ3LPmJFNy58SIpk0qTMLRr9XfB6LHy1AT
NS3KXe6XnPQJ24ptDDN0XPjYA9u1bNe9KwJ+8MSMIsn0bkc1XHWNT/WKqi25y7/c
Ma3ZCJj+xF8UKsohUeQJZ/CtgjQc9TOKk/s1znnKEqVCEFCIYf8K0MktvXgY36yk
ZrT/UWKmLeJdPOlv5aIs1GEUqU5yJHy034v39/cIuxwWXbLwJ4fQauFyVP/3nMI1
qa87CRCjB1Ps8ZTqO1QCKoSFUSu3KZ2jCxbbf8SeodrL7OT7n+SxZV2ryWTr9bmU
jiSywkg5fXvublWwFTn9qqgmFE5PI02RO5QYZCSpV9ifTUAM+C2ZAhqrkIoe96Yv
x8dJD+3ySzI6SKzJNIv0+zhWZAU/3AofmMZO0b8wDi/ZbH59DHjGzl7I3TbnydGb
7d8MfP1/FH+EdlrZewsz+Wu1zm8Kf+7juRh8rRZ6TuTMsZumISmMH0/4xz6O5Z4D
3IGeOfHVG8FKaFncnn5ygqZkvLbm6J1ee9Jkfe5qBE51w1427Aii/mRnwzV9gI8h
tOGeN4TrgvHBgsxC1GXgFQ2DBHn/KdpO8ZWA9yNoeopn+QH9Gam378/xU+f2JxrD
vhE677oFAtZDSrz/hoK05V55XrNLosUb29p4Y3ofIXMjWhX5ShwJL7pbk2ahAQ+d
ln++1uz1e4JBqu/zDX8qwuqZF6WpkT/hq2e/D/lW4j6sBzlI5oDfZCURA56nD7z8
t/nc3YpA9+/fcp03f5ZmLyG5XB2vrkbjt+NKQVs4xSz6SSinUGbIfoCRhNpczmFA
KZB93bvSv1hAqkLr5VCIkYj2wR28ifmMzxtkDg0p3awX+RcGmF9EYCeUxLY2dPBj
bAk9ZJ4ChIaZsQDRI/nOR7sGb3/GIvLaip51kbHo4SiFA59wpwOjLzKShoiaMC0B
oSlSc6sp+g+DS7vZFnawv6uXJqVMQSdIcPxMRwBM0ye2bGncz8DVlr+pv+4cDpgh
HY9nLo15zBsWMNAksaHRFvt5ny86hetGgUPUuL+ugfS0sQLQI3CpyGGnOHge6iIW
dx18WK+zRcihjmCg+JD3wd9aUcY/Vih0ZA0b9Xfxe15OM+m/EvApyOAskGsdbj+D
A4yRNeahTuvkolzS7b79kYBMfacRiYrs3Ci0WKZRtU9ZbXGy5WlBMwk/yLh0G859
eDyXIJmW1Zv/fuF0oTjzQIv4r+z9d1oviqvji1JbJH0LH0b0TepADnXcgf0zMWbW
ZO4iMZOOYfO0j6rZxKbGqgHew9WIm9faljyLwiQkMK88L7TofohiMefiUrsXOT9a
0Y92+1sCI9QaQVzuGzdw7Nl2xQ8ryxVQzMtD5TZXAzjx7x5nHq1uD18oxp4SI++u
A01tHi/Ke+y170IllPWk+bSawZBA75CrdODjFx3QnxZ9LxB2xHPLZbYZi0Pu9GiW
GZycm0KLQkz4l9YAovORlJZcNnHKK3IN3mx5YyQ9mgXBCvMRdukD0oAQaADWIz8z
/6O++CJb8f5hGwO5fJGMHdJ7AOd5jQpM0WvSQ4cmrtoQFTYSCJ7bRtyOQSFh1EyC
8MSolXN0Em+wvNGkYxVFYpWo/GaotIDvU578zijKHZvA0sK6adq8/UFduhbH+iCf
duDZnJk7VixSrq/obBz7+4zLVoRUzR5QNjl/OHTG1Wk4WbHkIq8sG8WW4qmVdQu6
EcvVGBPLXAfloe+wrfPETm0bZ2n8/wSqboLsc8HO919clRwBrNUubHw66yBwQXlw
aCFwJ/H9SeIbmuf7xdUnkL754k+U2OQwijBee/tV5W/Q3RXPgDLUd6UEH6qZzASh
7i2X1cFnEGjIhhuLHUPCAivvTx07pPqF14U3eOKSW4MOvy6WXg+a/nNZaZbi/cxa
mJK8FvYx4KEZqhaY1fi6r6n/APezCjGXzce/O6nDS1V3iSzQA5GXYwWF+6VGyByQ
KdF8AAHAjEbrywqJwZKH+yy4DB8EOozX6A5+DRZNOBq3HAShuD4LAEb6yZCYGgwT
fe0wJG/tMWPCVVyyZknM5vyUITY3Rv7eO6a4+SmICgNSQvpw5kBfmCeQfqW9rWS1
0NFIYWciT7srxJSZl2R82tQitAG4GAzD+xYgv/yhiONeXXFVb6xh5DswfEG3DGP8
ND41M+CJiQha628/ZdbQ+nwXxm3ttlV7si7Mjbcyp4HQ4o1WazowvsyuT41R3jW4
R/Cx4D8UCx3xtNCyahehLTYFWE7pYQjSqHndoVItto1jCAVW5MNkjvqaZVQL1Ulb
1pQOe32NWRWHdVvq9evs0V7euv8+xL9CuyMOLRES9+th34nqRK5EQSo38D+3fuGU
SYYgf4NTheULnmst88fdG/WWSo5IBKOUSRyVUf+Jir6m4016dSbQcnjjLvK8eezd
2s4CZc3HDh6TB4QCPJXWCWOsaIjUaHfr+/Dhux1lk5qRnAaslSZmGi7Ed8cGnoLR
yN9IJs2SmbBmTc6jOVtTrKY/qynG94qzNWUNqsiTOWs6pV6NAPLAWa4RaaVUoGmF
qC2pSDpI3Wv5h9nIv0SL+LHaRxgDvtHq0Lsr0ccdVfwbtO+1NcqyjeoFEvmWH2SY
nTN8jsdV3gBzsU9000N40YOp4w55hNIo+tTHbiRo5lt2scMUQqpKQCR93E3AHoi9
CZQRYBhV21W/kNSVInAtQXBV5LP57Mcg5PDU10ZJEuamjjqhTTQc4Oz9R9OVJ2nK
DuxDDm2g3sFw1mbO1e9I3rXTHXUChx3AtPJDnQ5NRtyRKU+2pPJlSjZILp+mlsC1
3olk0lUSN4darDr/D7/WPgBGrPXZ+AmikEphP1yrLCkuPuvSW0tRYYW1G0jlUyaO
sVgSD50+pnPnswK6AMjU6MD5vDAA0HyUYoozSNy/J4cMxXR1cT0ZuoZc/rJX4JBM
a5TYNOkdW6v5Ngr5wnBmPZrF01OQ3LxTAAZ1DVTRC9UvubmQvN08woz+QGndVE38
A+VD5iKNOvchaD7euxmqagh39+vIq1P+axwqIr92L8QyZLOeKwArpmtTBjxWf+ik
YaoumsEODJBsub0OAyhv9235KSYLe6o5CKiPyW/6sp88cVndOccYxBZOfSKTGXy1
a+lZd2IwP/mugRHNxqQVzX7R1W1eBQrIQG/5ho2FrXkFC+04Q6VGYDwicLlb8Pjy
HBAv0JmEUeMIbadojnxE5dF6T6lC9Yma1Bm31MkvB17eIUpj6LHn6zv0VVzroOxO
YQOG9bjc84UvTMy01g8uKoLcrFrmKqKTzsQqy9sngfYHsG2aEpVOle5ft8Th6GnW
CJtQGQNQ+ZpDGlnqexIU1t6uqzecnmesvfLTHusmwkDJMcUlz3ZaZX0TfCn49+ks
OTMfqSYUVPuNZ6aBbOuzMQBm+jxWoRRDcbeBmaXZwWfIfLEXFtEV0E/2Grd15dhs
V22UE7hxSFhkx9rB9SbSqWPog7MbbRhodjI+gy3f6KNKVIxOKB9/Nn8kRAERfG60
zydVO7nL1HVUXB7WShTACGQNKZuAvs2tM1tmmu3QLF0qJo1nKxSZdoONVL41eCxK
jCXermKN0+PCcPnMYlB6r5hLorMujizP5mZbB782dQe+zx377+1pIJ+3o8XTgP79
ZK1a3v5u2cZbvYNp7l+sf/xGuGiZHv416tmH4CCI9P1LqgKvp4X3Y93Ii7qnyTbz
iIOWxbSFrOoHaIrvU8ZxT9NLhto3/Iv9Jd9B9Ooy97EV/VlSPoLdISeWZweuqsOK
dN7LBQPuH7jn/J1UuaFVqhg2uTaqVj8H1qs5rsHNs9lNWQjCM/ToWI4Ut1zLq4Iw
u3AviRP2CObwUNWcu2ODsMznftfkiOD0cG9oiLpmBEFWLoAJ7/cu68uua3QfpoyZ
ERMUEEvwr8l5pLrJlMyK37bWRqPMz520ZwObxhGHkud2KcfgSvbZQY3EFTBmSJag
g+XUEp81MsPpTVjS53Klfpq93Vpf60Cr3asklDCWjFXl1iPsbMeoklCXFIkc2CJm
JZBoDKDzlS7K82lIBATT2JEXMuVz5j5+G87G7eYahvxsrOkMKoL+aBMDwNdjOAbU
r5brqLu281VkCGHgcX74V2HW6QfG1Po9TrocSQlbCi0imIJvijGK8lwIP5dzaA8u
D4xef4x2B014feu3YK5Q/syDRRA+Zc7pNCa//ePG4KY480iuLgM8YU2toFxnzOU5
ggzB4JNDftdWz8UzQZHtcEKLhL7KmjY+U0VEo36Wl4SuO1vF/vRZq+Jtnm+ya+F6
9Al4LVL2mXOP37ih2r9uAsxyG/BethE67K49O6pngxTPNNTsP59Dijm+WCHY3LGm
6Osb/avYR2mvV+vg1v6c/zf3/mMDc8LxdtH5y3pI+jKhBO+tmYWUSJOy1YR15CqZ
/cWHDoJb4eLJ0MUoHcxKiY1WT3T9vlwJ5J7QN6yib616R5XfherMnnuKx08AEjFa
iI2iASgyA5cn8As5rvZ20Y/5WSXlTBkEc2+pLPKkK480OlZuJ9q/ZdbgGU0WSm+U
deSJmaA1HN7gneJfbboT/KdzKr3nO2G2XNt4Tkh5kFRgjLPjOoWMoBlvBCeI/NJL
WHWPA5UsRdYzSgWh71fX0jfqIKOypqQbidYmfHQ6JbwAL263XoCZl4KzNT9ZKaiY
VayT1+kogjhqAmkMZ9zYVIIbRlG6AfvUxAVS1flG7U4l+GUTtBLaQ/5vi2v+UvkM
+ao/THTXcBZ7EPGM6DvBuatsrrPvCzMTdijTTIAecdAXPiNDJa+jmf92hSW8WAyo
14bK9or4pYzQxzgRmnLwDy6q8WVDA37Ba9xnU+E1+oJlaPYl35cfwrdOJBwbOUqo
M39usKNa5atOj3/TPw2ftmxnWsxfNArsm+tf1ddCtHWbABN9V9qCYU4Q+gEo1xbM
eWD+9ViRHLlVS2/7ej89Wn3zfJsgpJYwaw2yzJI5tyQ2rerLFyuxvJMV0p5fRXYt
po6MsZe0StglC+KUJ0wfhvRTVO0rhDiaqVvU8mb9JTxdzJF0dW+1r5YGyAcTINg6
qHo/Mg+99exPnLVvV8C2QcIhBGDWPnWf01Ie/AZh4aKeq6nKPuelIu5H1cN7BIHB
w//RcVQEHoWq2dhzjt9mCBmhd81qXpWlVfjhoqgMxFWFt+zy1fWp99TW9r91o2yB
A9krEgLV5hleHmrY83xqQFkHgJ+yYp2sSb3Rkmts0KivWvCD6uSLW9b6aj8cJmUt
+PwIO1A+Bb4WE7DKjwjf63tlDT7E8V4qMMFQsPhpEr4lIoIihUy9BwvjeQ3hBhVP
ioH1Fm2GPlN37Z9nkmyp/kn6x0MCPrALwJEDhRoIg2uVCV8S2z6mb/tJfl9eqxo/
Xype1C5nlpuf6V7GRxGAWzlXhaCyRj/Ch8hRcH4NP6ENhr59DtVEQhg6/UU/toIh
W9MBSvNa/YYgbT4jLjPIaDS3aVrClt+FQAV1DXKodPbK51O98wTK096RE72GV2YI
+uKWNqTUlmgagZaz/QI0pNb7vmfmmMQV/2EeWMsqU5ALPVxdcGPXWDXI7KpHfMzH
dqgBxNIjMZi+OqpIpSytLN/psEKSYcfdsKTdtZrj66b4YawM9f7l3+iutPq4Vokc
/rqjScdmro5c+abp3R5T0iuahyfo2dyCqmrVeUeZ4wOaVtn3RixFjmMyi7zQj/ti
faPw/Ay1PfWX1bnr3cZcTbO0SXJMwXkBcambGzNYkKxzfPysaqryqIbbrBEjcdI1
Gt7a/uvxPewBk3xw2opAKPaxpjExCiMriVqrX5ZYsQQEhFG6Iyn1EHZs3BXTZ3pN
TraDtdfpylxPBUaiLCH4rD2HB5Q2we4JFms8QM1WrLY+MnRxRLM0RtEuft++eMp8
o9i1OkKDea1cllJHJIm65aEHbPGyx03ElUZ+wj1UemCJgMCTko7nQ7V0X0C6JgIr
Jv9S7pOPjcTdjxrTJIa39ZSgS7tbNYkbM0BzKG8aVpy70dATTBRYSwRYhsb0rwYS
3wNxNfZK0aVNpV3CJn54sEieplcpRAmHr/OHuMOIK1Kza4hRan3mg3rxr83BpDHb
Wq4KW9zIMVRVDATRZSl8mvP0kwcO6w21tnCI+OQRP8t2m5H8XPQRLvyAfWDrKSwT
Be4XeuEyCUHZv8NLVS9t9fRnVRrfLKhCq7krtDVX6urYduJDu0AZq/Iuyd+I2hGU
DjkCx0gfUx/jBE3cL5jZTOipqt4+yKEij0Qc5PFwrIUCh+hgggPyaHlYCecf2adM
FIlr93q3pGK5kxS++Kl9MKdYb/FFyijqpvTS6cRjTDaXlM1zq3mj+XlRSNxpeWNV
Q0ZOLMkajUVgHyeFZRlJ/L0mC8QjQisbTNlEwUHa8BXwH0r5I59AieN9rEZKkljo
6NTGxI2tRk9r9uqfPUYs32mr/ohVeluLic/JQpTVsCDW2KTQwiL41kQVwXJBNcx3
wuT0IAH2T2JwIrPnhRlO6rv7hQ+N7DJ0I3ggP3w+Pg6hGTXbuod4Ai+kTNLl4Sm3
5yV3SrA14I2OByYSqpH/P9aKr7+tDPkMY9r9R1x7cW9N2drFt7kyIyPrkMRMMvom
0aT4jWR0hi2U48aKfgbkCP0eEiLt4Y8PON+pOKaRpwOh3Yz2s02fW9w/LsHEIHDH
dP1z4P3Rdu/WJXeXNdyTHt5rtT78Wghw8gC20kPuE64F2oL8ghEJZyqBRX9AM20r
6gqPNOcoZB5AG1Tfv/NdD+o7zo5/1XBUAQRuaK8mZAGrnSjmlQh/a2S4gH2XJA3z
P0OrkhNx9elyM7XB9uqL/Xw+zhOfi+B5EymxM3xpD/NvtfrGNi+wsav9CTBXK4LR
lPoIRXmSVrRAnsp9we7LrgVYGodTkDkmBVPLkhsoQHSiXEkpb2gNSm8vHvHKrogU
RSHgC4KtXWwvWPRPnyy8je84xMhpdRZkTymLYgD9tYjJXMEPj2U3vmC+24J0g6H3
gLtPxGrkbo/q9pEgb3YD6NLx9Pnxzeg31uPQ3RLLhdrK/nJ7V4WjxIfxuiMCkRkW
PbAGtlXdomgzTuSwpbh21jVzRqC9e85J1SQRu+tgd00rl2ECTAzz+27NlTrX2CLB
ZnV+XiKljKieIXOhDd9GQxLivlZvmVFW5q7G9+MEYOqvUBNGHvpJrJanT7nuc2AN
G9GjmAoQWreg4iv86fyKhVrRLl6ag4wswk/j9Mi0QeyJzRMmxS8fa3dYwBoFfp5f
PyFpdRQ2QaF9weZdPJ4PfRDZ20t62WmK7/VMO/e2lhi/OvpXzGCu9OK83M7TJAMT
w2QqnFHN3DWP2YuXxqvYvMaKYS7rcItpbBwPkA72A0wYMYOBhHxLIHLfiBhelfMb
OvRKq5Xh+Y9MJ9FzNi1Cuc0FCGWfJpM0NytFY3JJqOkFpFIpWe6Gclsgjq/gmbHp
JOVdpAx3Gf8JY2oVEI4Dawzev/dQrACfYBmVBeHS3PAhEOJd0w/S6M7XIEJ/uFDz
//sbZYS3M+iqTra2uaYJnhZsPJardmyNcXiTftgBz2gf5SPoVCqfPiHjoK6Dj9cR
PGcyB+yYTcArSLVXKW2aUhsZGaoczG77iM7mEVvv1ipHF8d5hH7Kpn0lLaOHwK0I
jV1ZG6ERayjZQjp3khl1bEUQZbxnlUrjqFVt0OhsYdz0JIXl27R0Mrh0oAOiijic
T2BfNIRgmldYpvEIZjWiWPXWZ/LJjXpMmqeak+gKjzbUPfTigKYJbmPorZh34Bkq
mtKvW4DJHtDn22ESaQnMhDviD1RbUCAmHFWkUMlSDfT74QRiCGU43bQ+MJIv/KBW
z8J6j07c7egRPSXtblf6UbTqRXjoGJ39keBniw4jz4hdQ0OkaG3+AWP/urbIDKbM
OnuROu45fphSGVAZ49HCaKkbNqaivF9fG9pYU1FI3Ql/T1c+yY+PhR2VMO3zkUbG
I6DAup189wZnxLGCBDGxn5Fx1E74JSvb2hTiIT2awl1JYgEl8ATW6hRZMeljnjqP
Zpm8A7CbYjUCT43lXcypzTFJNEzgj6H4+6X1nm1cOPrTRYnudB9Xqien05vTw+QI
DJ7f8oiMu6MnSMvPOjCnFN132MxgZpfLxVb3b4KwswLIxlKCXO6TEKzkFH+7/Su7
aCuqqw3B36rKOMBkjdd6XQuMH6eL4LN3dVb6xyrTjJwTXH36pCy7UXzG6jTwaNtC
BMxwKV2y+vMmn/wpcIuzi/qfmnnxKbHq2QjK/LuzW4c4vHJD+yCTjqIOZUiSoDLt
xXe3PpDpbrC3gVOoCd1TwRIdMkilodGaMMVvWJkWF1nDTVuAHGzKcygiQF1uF9Hf
wRwgYX4bmZhwoswKmJUg9RZuBXXXc3TfUi0BJpnMIAPZfZXA6o3Oy2c0wQzyg1me
B917OSR7RBw6ieH1ivAD7yuv7BIofENHROkKrHFdXx2rssTX7425ZmHMlXBu15wy
fkfwdiIxwPSXhpn74EXyMKL8A9UqAf3OoRDL509pJnLTc66bFzU8r0pSDk5cw7x+
GvZSvalflF5sXJwI6zKswvZOpA0ID2eeeg82vTPSm7UbtsewQWyKx6zvSrGoq+ZE
S+H0YI+XXZpec6I22RBBFPcFS8PjfZ3Sxp67eOS8SxJOq43jSyYlCKNi8uwvplX8
tX0DaoWlQ7h+CttKU18WH2jykRaynxasxx0qyyUSIA5zZG//+yTVDa+5VY+ginsb
Rk/jtL8NB2WVYxS6PQkyL/44xK/b77y4cfgNaM2UVfScCanC0+ZWJuHF1jeiCJMt
mrRVErmnEE0I8vGKYzecWossLYFmZuZ+Q5tMSO7VEzIudpRDSboy7hcNqHTvfK9o
qKbRdz0M/NCGXkP9hCwsXzAlB0GWKro3r8jp57A7CrxwkOeeykYbppLZpKBNDl77
XNgq0aJX9L+oqmzIST62xNcskrZgEx3+dsLIxQbWoYB5APg4TAqULu8kq6c81elc
fNOiHgZUeBI5daNshje068XUTsfQmTKe9LOm+jVDAqLFrrbW/W7ICpHUkYiKDhSy
dJngKow+K0z+lYS+oKPm8kz/f5mUqZA+QA7/jGJCXT5vIWv9yBHSwY4XiFqw7/27
18qSxyet0X+4twu5ZXOyN2HWwh1U73zjjJERAqzusuwQduqzHMTkTtgG0rfif4XV
y1N69M6yGU7P9QSphJLgjCyU5+WY6VCoxJONJlQxaDLdzTnsBqH78fzV4918wNia
vW8cJ5H7gWLDjEL8gwawTev4in+x16GFylvLm+XMGKsaYw0X7CDa5HjujwvTR9EC
ydgaSzbCBIrCSUkQX6wR98gsMvuV961O7OaCmoHREDmv9KN9L8yi8jlKtRHS3tKt
uLF7jqiOwUIbkc0cA8vi1cw/SvX012jkm2+pLw/sfdTOJ7YKJixj3YL5wrapAtaD
9DmuVU7rsoPZPHvq1SUUjEsxKEX7ghjgDjeKDH3x451B1EkFOwSiEqk7lD9kiMc3
2yNeXUlpEtvPJn5vVwzKB+VxwRdgd1B5JENjZJqsppF9lpc6Ji1lWCTgWs2XP0cU
CfZR6lQBkTKpiCxZMXRw5iQi3Jk04rkiojMnM4dYWW0XzpV92v+PRdJmafL9XuiX
K6V4BkjbbPxsc1wCHPqdeuKMIpbz4EWWmud7tIrdQs2kOuQMGBKl1DSK24DkQJS/
2aVSq/2xjJzuOxU+K9Fs1k2N8MD6dT9J6mAVHw2dDZwCEoxrTnlOvhfQCx+PaNoY
qMHRuzxt+sVSzWWb+BfxSgBKppcvXsaUxtzzvcvFXIwxtMz38ntcYBFdGp8ihHBI
GmEtxQyemnX0+LnWLUtaAGRpYFyFe/97TN92IdABMuqHlu2keZw5k5HNcXDSDn21
8rPozVmmIMxsJskc4COdAYShhQhP0zSjTNuFSmx8LDP3bkenHalIX9dVPCMKVdkQ
k7T6p6bEk2HGj9lx6+Wke/gUH8Tc2V+y6H0veWHBtcV7eY2JHDVulwIPiZHSn71v
HEWigAgzyXc3vhOtULAbDwbSpLhtAydNO0RqiN7Fn9VkV0kKQ/FS8IlLUzDYIo4B
dX1fkULx96txczK2jHgDehYq5ElFugrt3Cei6N7oOD6Y9N3nZ5wbEHRjgNV7v1wz
1LcHM5ycGGfYSlcMZFVc7CtbVaCZIquq9DYAbVa4ePcj2jpjjrQ89PyRaUcA4MaR
puDrbWkcNW95C3q/8/kK9z7WbzeA9PirWhrEKJV5qOehliUs8cm/jyr/SeHLqsvK
31nh8mWePAsGgZvCa/CjnPXc8jQPXmQLIw8//ucXrsYgvdyuWADL1CcQzA0b1+mB
+EfPBafgvty9F/NvHRVOYphen737KFwe3wkFytwSDrNQqighU1PTbufFFqI2FhuK
OuOim7JBsp4Ces9nkevRgau8MoZRRf5KE4vD5D0iZ7Ky0iUmP+a+18XpbrKdjnw3
fDeYJw8FRKQhY7aQlUrGAJ9S5Nf8LJU6pifLP9fiX2wke4oqSEcrTTWA1/p9XXve
rBVqDesSfSXH6picuNFLIrzLB0X+aokx/sykp9DVsabarLc1tCPcUsAiLEzzX09U
daYOusMsXrDY1XYdefXPqcbJII5q0ekYpGwW6rTEwpqwgW0g5EOnAAbe3uyH9Oh6
pTJ+7sObBqkkyw2nfn57fcn+tZYws4gly5QuYAFB18CeTdJt6b0xr7ry7FM91Znc
SOH3YntCwExfFkoxqm50PHwDIkHdlJOHhg7D2nATfXp86WILb7TuDH9hpU1kHFlS
lVHUaifvjlgWqrBTGShxUI1OvnIPb4Z2NwB5RWz3Lz3QTpQ5JPGCGrfbJmI9fTXu
az+oAw1II8+IZhju/Ur1W1WyNzTZB84TvMIjwABtpJ/8Up34mrkLoCoWnFWa+ZiM
GIWCIJ9I1gkexVW10au9nyDMBoHNykMJ2M3+G/xUeXCLjrrpRgIHVsv4jqzUytM9
q2Y691PK4N1q+pr6+HKRewRLLkXoGGQTfIsxcqaiMu6WiZCv9Xu0AkXToUb9xQmQ
ECp4gPeJ3gQoNPUTgMQKktgGWavn1g1S6k1i3gmr+dGoGx0xL+LS2pFvEtT0og4G
xg62EEpPG8xJJecp5+vcW3OIWiHizrLRD3qJcuerj8sZYj7fxmw9+WVsM10/+GBR
LLPQvQ+k0BGxQ3H9GIRrTEEmtPlXBOXNpCJQ4SuB8706oPSzZCxKUGy2Vvpx7eoH
EGMhWCPjvp8whGBZ2yyeWupjUcVyQaBBTpeNrarj9kfYWJ30BDG47GCUFe7NJgSK
23AqzutcKISV0QwG5sW9zesUsFITGmvdKJ7X+jkLKhSP2bXhC849Kd3n6kedQMX1
qZqWyWlORQdrwdteYsmuelswBOxKBoqSCJviWmhP5h0n1Tuz5838YqKvIZ3saMYi
TVSdwYddEMm1qbZg3nBXtd3VLzT+vH259nYQmteoBBpBYgrcrDRDEWwH6dV2yfjC
nwwY2wf6KVzmfZQmMSIJ1Nf8GFn6YvOYbIRvLNPel7+hnHNfdikI0d74Y00UqHcl
J7PO1PWJ4eKGqj2glW0L2mQLzHMnWv48OgtofNdWV/YM2LZTk3jr76eB03Hdf4nk
J9xRjOjuxoWL2PuJ+rPDyEq6wt9oCFylF6/Cb3789jNI4DO4RWFWcM3PT4+EpRuU
V3DHvHxP0RhPTVplZSIjbv/6DySZR29YmUCUDDKUn/W/hJwDacRK4faeBMafWfrT
mhawm632ObQSSu2nrYQoqWIq/+xlfwu03ff5DI/9MsmoMtO32HpKUFAdWLV7gMU3
iZ53p4LuMkW3GT7eD3GcwePC0Adh3343YVGkSsRF9pGBFvWQafOvlhCyypMVv/tC
vo2D7RKApPalf2flmRK+MzomIACN0C9LUdW4ihhmzN51pRh/ayoIOD1QPwgwxZ0V
c83puX/232KyMDe8ThIg+P6Tim1fUALsv1Qqc+MNypYgTeWmrE654usFwb14IzCy
fZeogDYX4rKyK5GCKBbWQtOoYPOeir/6SQEWButM3iCSwkD33vgBvqfYiIwcAibb
PPKyu5aY0uplDCXG4xF0mh8PoxK8twG0kmBugLYJ40K8RfoyYHxPbDRKrvDxY6mN
bT7vXdJjoO1IOOyKYwrCqUQPHM8AuXVI6okraNFtRWOzHw3WpAUiay5Vtu4YDY3U
iBySehP23if7hRjL7EYGaXGghRl2M2y8eoCKB8BsdmeOiW2VfZD1gSvHXP216feD
YFU6mBbSicB51ohB3EAyi57eObizs/Xm/2S18fAisE6p91YLzU6MSZsMB07yyUWi
/m3MPH1hs7Cw0g/W4AYs40YpNy6Ta2t9sZx+Tchv6srj0ppb3fyjBJ6h7/iV8jcN
l051Ufk3p/EUFupHj65s57XwnSzlEt6vsyu/bTR5YTcw30dD/XpipbDvYCGCm0/U
QteAlWUl8FWbWgiR5MVUoUfWC+X4VUeXTygkZn+lsc23ns0MbiK1K3nbiENrQfTG
iN/NT/sfqOQFzOB4oCf4SK2SJsEJTlkPSkqs7YosZHp68d3jTu3Fvl2V24QAVCRn
XtrEmGPYqrysVF0xUwqAWtWabbiYWs7+v8MtWpMN+JEF2Q+NOYKwooZjrWtkcnFb
g3C6pv/kZApXn6DZenHJt0ssccNs38YNNNfpBmPbw8aOanleCgI+bdSgo0CNvh3S
1LAb2cUMm5tAnIXrkl/dJ9d+4B+2LZuC8kf79yU3qLvTEw4V70SCRpWZIMKq7dfD
vRyfH4PeftdeShYpfZsFPwuPpSjW4zz8FUOUjJ2jR3cJd4F5rBVoBEJ3g3ChTM8l
XsnU2QcdZTd4xkhATB55irVBG3m0wWaS0khMPCyX9DGwS685erLqP6QhpJisO9QM
Dbe9ovWP2jCuBku+Yuntk76ncHxiVIeynndg8EzJ0dIbZb/EACZfgBgceruz3Q+q
fjgQvt4qsVDq2fgoHWGlFppXGx43kDpazp6x4JJcZ27XDGw2POma4u3THZbxKOcu
cMJx733/0FLRXfohBbNkhdw6ERe/wuGNSXbCzJ1e/wSkldna/FtIilvsrtDb2aAv
Bzo9AU76UAfs9nUPleeiGyBVsiVZb1GAV/tgNb3CMVx3/JJm6SspmxkWbdZfk0oO
4zwcW4okzl89wUMrqbFfvpOgl4mVVYEbFI70JyPq8bR7jPnRMXv3oskIQpIILdwZ
efik0ACrZb1dBWZVUAr4zwWKIGiOGdaM3yUPHKRXH+g8YHRrdrbRSP1U9z3R+MnA
TykQVqUmaNcaoRtgLny44E43BMUBxNiw0fFPw/T9AgUbhOp/4bnTwLUseGfnSZoi
GWKUgPOfxYBC95iPQYTfXCw5/Vi/0th5np8GKQrSJ4jb7MrauARe3u9Z3zZnv3bs
mHUZqNrBlkzQYn3CV1G03f8OfRS6ZHM0VxLAxke0Cxy10PSDztx+8urjac2CzYGb
mGnylUYlYAmHHlpG6Mr8M+Z1rE+v31cUV2figfc1qIVW2Yr9cO/Fnsrn1NTepHbj
hoJv8E68kcX+kcDmK3LQPBw5k33/w9R6CIwdnVLuPX+hW3wy5WEcFW9TwfOUxZun
BXB1AYluds2RhFEjbOLOThJTn5tJV4qFMIWEBz+NfrYuJWhlUtlJOAGmrT5jpFTQ
R/I01Vq0vz93ADPf4cWp2UlnI5yPtETf4AFtoo5ujhlcvF6P2OVaShidzQG9d3zH
iBXWPUG3QlzSMhmVdYF/48d/9BI40pbhPW9XdYsp/QEG6XvkyHr02S+8Wvztz+kg
bIr2V43qowbmsnUa/172pLGDuPBIGlNe2AdJc52QTh577PPgFh6d9Sq8PqFtJgle
+tWHNgjf36gb9Ur1GBNZSsE5XPm56E0wHBk2OIPNAXdWpLRFwieWqneRAZoE0yTM
0A5SSGhSZjVdBKu4VzgBuFjMGFegdbd9gS6NZk9alEFSGnyQ6NXhf8rGlEbXar1C
UcDJLa+MEsyPIVCSKmhQYsPNX2Qsh6BzdJvs8sdQdEEyBO0E+mUwMG2uHxRvoiRf
cbY9W7ZJe7SgatHPA27e8TdtffuluAp6LxHfKILOEPMLHPKaT4X+dh979KhjyN7H
GB+bLm5psfAcWMBRgEvln3+W9Wl42hB3ibLVWM8b8mTalU9jjLBw/B4ck5c8wKPL
+w6jKRbLclYXHFyAmaXD21+zzavfCuL2EC5Qc2KNo8RVX+VonYmWAafOLF0Yagin
MJzpNtr1LYpqNmH1hnao5UcxHFBsMGpOwGAXei3lRFi+UYAl7L3MH0nlfh4NHBle
E8OqID/xrBIFdjoo8ff4i07HC/l0KWNEa5KP8hs3HiE5WolQgHdaWir/CZMouqHn
Sp5gId5PheVsyEWAEzK2mVzMeB8Kcd3UF0RqQ8GLxztdZpT1GbNHZtI5/UrDD4pQ
us4KKDvsbkebJf0fSDUZzICheEXLRtyDhhysQcosh/jO5Yy2Zr0qrlPu2LQswYr8
ds73WJHIg93JKMPZkADY6J8PtFLp1UaBint9eFLLDkV0/WOLwVC0MwSjbVPDsi4C
Ei3aRibKWGej0QWsnyt8vYYeoNXX5Qw9ggJwyxswNRz1Kc2jgEPbnGFA2cjdTkPb
VhNRWOdI1bnIFCwQyf5He6nhOWDX0yk60u+BQt6pkkjd3Gmjnf/iAfpSjAyAH8hx
9iZ2aOwe3IYlypgFaopuggto8FZDDtwInez/mEQBlLMhPY6iN6MnSrW1PMPW+y+y
XG/vlmZ5uXJIoBKPVLAY94Odcp3oMW5jwbpwOEyNgK6Yyh2PXWt8uQeHluFwfTol
KfQ0TrW3nEy8A4D/1rvfzvMxFUVnQDWpcuRwDGSzF9x1nM+v8Rh8AvyPz0FKJDgJ
WAkl6aKdAhe+cwARYmvOzHu9hnCPF2HkcFmr1CEcrU/AeW8HJI7RH5xmSqxlP2Gn
6CrlteTUj4CcnTdmYmX7ZOrI4fHmOyOlzELN5j25sRw79Jy/ZuLvDYqUoEeYijf3
LHnL/4FxKqR1AommWxZHGZHmXKb2JJoo6nh5pdnA7BhKHDdrnhYl61yKyMWlkhWy
rq6KULlxqytE0D6JjzLprmvUdNpo/f+Ydk2dmt/JXeWd+zxyBvUFr8LKnkY42jF7
vLJSjzoP8enxPPlp/oF4Zvw4JrB3tV4PuFWYYLQ997K6uSEoDES902ObmM3PZvUn
BotcVUIZnyKvn92WzZ5BHpArKIQQ0rRhIlbWY+O9GBDdkhGjiov3Zip1O0zE02/w
SFAgEXXn8eVnO5/+011G389TxKqWux+nHVa/Dt/9TQXGH77NKhp6sl2FS1Kgyjge
cKE46Y6pBAWfmHSOtoSiXjxkszgqNUny9cFlovcSSBVTaYGHqAN/sj8ctVuk6ejY
SlWAuodkcW5Zacwmg+iaUu/4pOz5O4tbxfo4sA+Bk2CkSgFpA4WZqhiL+QirV8e7
1Y2FCimrF4JgAKezr/0eAN9ztsvUHTgSN78s7ntLiIvFyERLbKwfVuFsdamn7C2S
CNRojihyDhOQild64c3b+2Y+wAK6Ddil5eswevBKkr/Vl4zyo0voqZb5gNQvBPio
TJ1gfrD77bpPKLq/ZIS8JgulRNJSxkGpa//8BZQJ1Fgi0EYutYA2K7bxIgrhfcUf
TEBfveP5hjFEeGWuEsdo+eMrq6PHOaIOKyEzhIy3KEHsLTWhaTamhliOIcnmLV6F
Mev5bj509RrT+eC1qfA3NzgAKbn531GHuxR5zDkSe4HBSKhKqhieGtKnBR/k+YJ0
19Ni+urbgEkZkcz8MEQmw75RR5Bzso7wfczMps8BtrStC+do8c2dQF5bqRe/xMpL
OTJD3gndmQM7Ku4LUjd0U5yR5khschQSXFTjvYWHHUk6vqCdmiRgp5l7YCm44XAL
nRE2MOZS9r/Ih7xfDqFt9JmtqDFJeeKDDVK/TTIdM+hPaxVnOiM18X4hYkKaZoVA
AYL3kseAZMEFZVQ98Mv2iu8H19DC3KLOyIFVi/sA+49uJ4R7VFDh1iHBTdPmXihP
9tyaiGELUe7pnYzw1I0AbtXTClACZOrD/Do88t+4Q/CGKZfWbRHvruwmj2Q98e4q
3h4C3buZ6/XgHeSLcCZitffRKaqvAMzyLGNwqvABXdEcXknIxbXGjweInY1TxQ4C
R227amN29r9v1juTtnMC8x8vSa3bXl72drWYrPSteEn9RlWdDxhDjDoMoo9DXFaq
ZCaRjOFhhaR+FPtmvyYypJHm/PEvkjcR/OaJgbya1sTSUuP3mBp6l4RG3khH2vuZ
dXE2xPcE3vTZKiiBMgpgjwNRoKxSRXtRhS9K0TF0bJxOSWPgO/cbw6f9I9AToONc
twnmrWScPpHv0jJgsBhi7t31vhNpZDMPMtYTfq+0Qk6lut3FDb+FNDWdOWR3O+ze
fIr2rmeNOJcWZoBE0rQAGknluZPNnftNw/QmlBpz0Anrx34IjAMQ/CbAwWQnmn/P
qeyGoyVKX1k/axmrCP3revM82LJT6yqh6Le8nNHEVJd4hZYRHV/a44Hq+VzBFhHN
9yizYWALxGG/3WFYwI0160nLbLP1nQyuRGneL5hiMzaGhDBXNSs56fHWRU9EGRmr
iUgkC7ZCg7cMQwT2dG86Sf6+UQ2jgSuvO9NRUYy4rfrqkx2Fwt5oedlFqT2qm5Zb
dakB5aliAgbOLAeXzRdDD6qPn0Ku7mCbs3i4HDk6uewMM72KZonEShRuYxleK+AB
Rhv3TAVLPkM6LvyQUd339E5Iqdx0UH8cH3QDCCXMnnnDmeuzm0t8B/IVUXcZxsGs
ZeE2YumXPWjCRmG6oZvVg0sybSXqYLIueebMfmYJ8BSoJxKTnoIHMkyizJCxgaBH
VMdi1v/aLIn/YqMITYiS2p+MvpSWdAu9mPGlzl3YVel5Qg0PnLiY2lU1mMub3WWD
xg4oU5sDiCsT4X/9WV+Xfp2+dWhM/PtLCzH0xcDwYdWOtY9nvgPP0sQszG+QL1In
paYjPd5XpHWcNVQ7kkRvhVlJhIFjwv70m8i5uRjHSCUBEweV2NqiUCk3aKpmjhSR
ErxL0ECxp9gJwnuQ+k19oZbrVaSR4Wcm5zYwqAXRj6080ahr4s5TEfi0qQe1hCSS
B1okXGpgunWC7jDw18fDnaJ2XtEZLenWHKFySLMqHZtUC96Ez0MHXGn6bObW2f0E
Z0rvd7nbJDKPahMHWutfD2d8aSnTticWjEnaNt5sreCLTPhsNlUlVm5ssqtX+X50
Xu/WTjsL8ULqWvjsL/jG7dOBdy3vrnjZiRkiN5mpZhq5vEHHyEo5UFftZ4zevgc8
o6v0RI8Ljvac7MWRRjrtEziaWBJw43JeGuIECaedP5NsYXCYU1Lvu5qzJPM7wB9P
7RGGZTe6Mf86v77DlG+xYlKqPZiCFst9BywLp2f5x8m3EuxgS8g0D43Rj5PZ0hT0
gEEdO/C2BN8/W3GP27STOUGS+YIl2uBoRI5I/CBrLvGCoUNJT7eOqbYqY3ow6JiO
sbluAlDvhbi78ZfL9mM1PGHx5SFJHp3jzeS3ScqmBHfgx8xNERJRxBU3Wp3jM6YF
c51d9+yOi3jrXsl3Is852FPq9JSKkuy/klAPe9GOkXJydtefKSXA82EoaLUfiimB
OMfblMPg/CbmIFKuQdE6NyYEQ40GDrVslBRfWbRO9sGKTHktyHAoUVmDCL/IiS55
lysrYhCTlPitioWe036XgJtr8X9UWw+SEUvCVCj1quAw8cSdkaTFtVDCZLufVdAN
KGEgwfY4T/2r2byoM3xOYDF0MxMWIDHdfpBmXzRCTDbyNy7K3dL+AoPQEBEYY5be
U+1gb2TAkYPABCEtlw/IhgtxB1K+4mtquiunZJ5/o0fGPD/xP8Cxp4Do7N5KCYCj
BEieK8PfYywnl1cfuRVakVWP6krfSC9pCCNRNkpVAcxH+C9FaMFCgSft4t447EIK
0RlZ0heahZOJp63Nz/KKFIXAVzLewTkixzioy+9JkScYRL+GuA/ZkoOppAcyVLmT
kim0XCyz0hv5czi4vPSipVPTjHVsHt+M3IOvOebXSHBo6fHAvP6gtFatcpbDZ9pb
NZWJ8sE+WpU78awnlpJFF+HeUOjJtfMpxGgKAU1WDUQ5LsWypva/L8lTYoEzyK2S
BzWLh9HsKt8qWmHWZbeGPb0GHReRfadiWfeAridAgtJk1TPyiR8BjlweapFjPyz8
uC2/6h3xCe6CeKNgtBm3iH5wjDfpMhgPtZMwqA/CoZeTBHUp3KGbNpYAIarD3Woe
UFlraeFcrU0GY9Gbr0Adz0399pR1x3Ql8vSJWM5mM6iHG1EbAJgej1/u/9WNjhc1
FhhausR9yuFGnkyr/vZ0kpJGsX8GmhsVb00PeK7glp9nfzAptMv0C1rsHaRSpUr0
pPHnU4OQl7EUDJ0cgqzssUjsbZVWft3JsZsz52zOrKwywm3UVAORgXZP+mya3L8Q
q7JTA8hBXgJDmhVlqNKvZnvUCsRr/RO+gWvIFD3J1IImPhb+9SbOcQO1lTSICgg4
vUfYT7N1sRGyArPm6ZIlr6U+GSF7EyKEBgAhLqpGU4FLg1uMUSD2XLdwxVDUYClF
TV4KFG82s4PEEVAHpQXE8Ui+3QsLrWy88YZ2eEYQEBRyS0RQ6kTtaht4GOm9ilRt
ZvzCBrf/ESltK38ayxoZ6gVobyK4t1BIgPYf1C4dc5N8P5yjUFMT6MB8dUbwOuoO
f1VSCssqCC4+NpPitWDz694dP2u/I6B1XkvEwl4AQhu59vLVb4ashIMhcmKBWbt4
pSN8HzXrlHttdnULuIiwaidaUIkGh+uqtGFsw/O4Yaoq46j3X1aNKNkMSriVDsMj
uwrbDTIKkt2nei9cxKQUkHHeCJGZd6sR4juKIRb6yjW1xZy/DkwCzTYRpj1qdTe/
XMTOvVDcwgqM4HUv07eI2bqJB4VgDyBjorhb8cFMqfXSxTH1sCg2smkMYUywdHdL
6dlebJWGvg3JDZwHhEhXDk9dnSA/riARve3Xkpx6LNjLAnwdjHUniO/7gSrC7cG6
T8GGP9BOwqqiE8rTYaOKYMpwCDsSlfxwUoCq808C01z7Qtb4z3AyVbpyLYRmK7ZV
YXJq6HQV0icw7A9ebFu3gRVvZFjM8N7zNNki3HDqAq0Y8shUzEC9hdIgkCqsUo2B
KJXu8LSfAieRs5AqkOiJcqHdHllU4/T4yXoujVYqe69DO10qSm/CJVzku1YQOr2m
+BHVqHa19GJyR+fFDzNiLj0OhHhU4D42y9ZUyBqpHrVWdVrh8YpBdxmoQJB4TuNq
K0UnPx0DwhRAUuUqOJzTwYjfUFjTd/siRSoO0Y1SOp7WAiT6mOdFFLxUxGkfeFoo
lrWM9Jxut8FboQCgySaN/h8Cskq30MX0UEK4Q0Qk1GMb4slLDW5XxlvCHPyfFEZn
xGVUQbyzH1HKfbETdxM3C1VwGpN+PGhKNbK4GXFpQBbD5jwAIRhlYG/GTgHRbNUt
S+YqiJWLhBg48O5FbZuxp01MczP9HpTHUObjpJETPbtkr54LZjNBbd/6luC2hEz8
DyctuKU2cPtZcqLtLyJ04A4QbUXC0WmX3f5AVSxpN36eiSLFYtgCvtJBq/wW9TTD
Tt6tYQOAFpzJPOoM0eRkENoO2VAqJu/00CtuGp36LxVh7/CF9+lePUX+IguXMn69
xb6lYFUPDJ0WC6LxqFA6/XDZsFYwVz2syowCGQlkvqtvlcRJOak3KQgsJcwl/qHx
1A56wabCt/h8MCNwfu1owgzMpIaOtAbYTJu+oIIiar3gHAsz3eznWubjSD5ggxpQ
5RsBoCy3d80adedqAb3WAZQLngWBFdFiPKQ0RdXdWnSKn+6gob0zDorWIZrmhtxp
Ke163hNNAok2KrzVXHW8dQ0FxXflqpfewamdG1WdPbrKj2J+g4NpQhUgeT7cQX/y
JyUKVQgYErVKPD/eTCnyZ2YNTwn3qHcu/IV/ThG5KZk9yh53gZ3+CC1vJMUoKMiV
HYWN/I0/xD03UaGZ8YDlkuCVBZAjMJ3foI6kIdFPKdfPIsYVT7ELzE1xRalXgxRX
K4j5mEcgFd8h3Vv2o+NJEaA2EUbMBCj8p7kakYMZ6N+ZD7f3GJHUTspCTTcj2ERJ
tCaK7o+S1JQ9GByi+AjbFlrf+R/r8XrE1t3e9VgbzMZxeNFGKDoUVvIy97jyLX4d
/TNF1B0MU4mToND7F22Ry9CflOFvUZUB3N6RgjVBxHPxRIfqs9/KZfFzXA5Qy2EE
DoUSN4C31czRkg6oMSk+/hN5pt07/y67QoSEaNYeI5UyZQUq6HVrNFSSI5eQEOQs
5cyO84sV1Ri0bY8YlVLu7PdyIU9kI7b71Br1dQju/Ol6Bgx7CktKrydMdXNTpyQ5
gB/2bPJKEm89c0KjzI9lWVk9QKNOrNW2E2IJWHMNLE8W6JTXACJaJUZJGPBkJFJ5
+tTR2yL0QBWzHbDCz1UHb0uMEuKpYjIhNOtVj3eQQaam6GTz3fF6tT+EK19aiWiE
oaNcdcOlNrYBTjdO4IU5nDpXQ4b1e287Eycd7lqKYXoyvS2XjKGxFUjdHYs8cs6r
6TC5KcGBRcsw+ZGiJtQMGEeuAApHJerYw6SocZDHDm26D240dV/aliT1wVmfcTnc
aqjfHd6VTj0/TcLsA4G1Q4pzYgPcT8EESWSYgv3xcbeMGnwkNqjWeGeHIPoKG48o
w8v1WzhtbdFKzzlQayamoqh8ohJtj+DoUviMCb+seauwfZS9BTtKRRa1nFuZB8rt
9tf2VMkV95uImUxi4ADn6rafql+V1vDT2HqvnWZwy+2utLADXNhYFdwX3LzjU+42
BbM87rvXG1EP6I7GFYwlYmGWDyLXHxw1oJNxY13gZ9H40pe8fLXjQXtZI+CCT8tV
e5VC+unU/E+luhYc4hIuxjCvvenkI3MYeFtTSLrBmCIRk0h0K08NBMvVuAeVIMMn
8amgfvoV7VLRyEiwVZzsoo8YdcDWPFoRJjF/7Kaxj+LnR+LS4H9FLXTHIvlvtLWU
9hA31GSwph3tpDlcamK5hDdaMVCOs/1bO6hYpx9+usSWxNMEQAdBJgT2BgUp++kO
APQx9ZFgJSdHZVZ/SrQZsUuI660WCfSVjA4Ai9nCoULuV12cX4OdxLzXTD2DzhRe
TIbHLGABamggRZv7o0wILYnPoBhId/N1rI2kkiZYMDgpCM5Pf+O+/0uzUDU4xZAO
CvRVo5f5GTiiE8JDJFdq0clMsOPlg6Azcbo4DVwh5YXNjjDMRAN2wZtWam4KxZss
l0iabd+4h7K+dNL7/q4Pve4dokHuKew6IAKPQ0R8HUC62L8Qy8pQ2Uz+Tb+ZSQJ7
hQt3HplGb3uFcxHBmzywrtdbh7UQ9hz2KCH/+6Ijk3Hf3SjVFfMVGRjzyMtmeCUo
0lR8npb2TYAfyFwQVPrwvyFgQ5QPuc0uYHmFVH/rBQH/GdWnOBBgm9XjctN1o84f
wTvidre3TLnvK3dDfhVwMWmd5ennjyjIjPDKxGBkRAbLh5bylIcCNx0i9CRuyugJ
M9QWQrr13LAWDQ2jj1D/MMJfOxvLbD4vAKSqAP3cgcvIrX1oT2hnldo9bSwJBHA8
wby+Iz35vMJ4GcAeFROgd/VxeavyPH29utSH5E3VLjszkjY2qUsDunxYqbZHlMwR
/mCTEkNe5XAvZ60IaF3OF4PU9RvjhJ2TkFSzObDVRIXThA7/53nz10Oq//9AB/YF
6TH8dFOoH8kBBDsP5xp8GkiRjNJ2nUc0eRsveVXluwj1TPieCObCzPuZ2ZfvgIjw
ixOSBj/pokk9JWG44xBB95Z3R2etGMZPiW11zZUUunrbL/yqyTpTpLFPjwjYh0ei
IZhAVp2/q+Jm+XpsPfdK54guTOykvFb5bfcHUBjWxpUn29GkgY3M1ZVGI6wa46+a
yUFRz33ra3Ar5spoKHk+UUV7ayL+CIHryx9UlVjiwMKBge6Jv1P9ocVO0MB/cPSv
RTqWJ9lZ++QY/IXHL4bE+GsKhMFy/1yZTMOJ9Aoh+W4ghDdIflLxeHK2jPjthFFm
XjlwETodUoZX9bQFBzLfYVGOtQrjR732rGl4BfeDw0HXoarX9277q00kGzuXTknM
mXDL/jWdIWwUPcLcEGa3s2jqwb0A1r50v6p62AsuSV5RVjtDy86m7IXpBRa28Co+
V/fbQQgXMSUcPSwViyWdi2iZQopwqs2AvfTGaZyQMbHeb2YG/oeryYb8iphC3zTs
V1MiZniB5pqiV4oZrcHU7tgJC+wlQLq9z0wLS0HFjGbWcZffhGDoKv1QxtsIlKYV
iwjCRgJ42UG4zUKNp00K1wb92viQgDhXfqHGtFkXjLRrxbQ/JpfLyiQcsb7Q5Omi
bq40rDr+5h0RgD95ela+yomXzyzpy5kmqGpERYr3YJ2p1b4+2I+MPaE4R9VNsV0A
LkmjHatXMrgjReO76np7lXDyoaZGH9YXKAsW5KyVgmx4Be51+QuvJy6R8P3Xmlya
OuCCF8sv3l8k0Il0GLVlPuPbx4QK9DpxDowRIwFSBHqGNKKHpFhYdMEM8Kr19rPI
v2IxllorLMpHpmxmxqS0PVPlUJFfPwn9vAGhD3GcgG+GKnXaAPARKbabd9WApL6H
zMAh3q/xlsaYH4BYq0Sj7yJV/LZ0EtCZ7MWQ9rBo9q+OjaMDVaEdtWMrtELsSwS9
RVzMi4dfcmFmjq7XtOa9ETntqBDPEsTXA+ieWT2asmj61YNuiSmdZU1E5QNm/zZZ
xO5HnXzcJi8OD9+EOS3Yw6aqRwbDkWRHpgu4rETzWdALJO4S9tT4iAOX2otalu2f
eeqWImX234G5pmmieZItTavQJAgqwnV4bHELaHam+0+qUXHPl1vpAgCtwroV7NZP
IKVu+9M/xazn9Bf2LWuBqIe992MULgMjXarr/O0Xhecd1sw8hWIfJ1uSCuYt+ac9
Av+FGiwqwqI4Jj5uUC9SfLsAR5hUoYonCiECkl+kTSdkWzw3poJl85QFyp4m9tNo
Nj/82wvTr+ejW9BUBRVslRMBEgSTpYkbgJfZRdyWs6jDbPNeLsBC1DmFEyAi6hfj
MWds+pdAs6To1fPzZZyDq+JV76zwDxLzwEkFcrqS28xHNt/Jfg/UVjzE4c8SBJNW
2IDeSyybUwR7EynF8n0TaMeBzUF9yWV4trvWxlrVpzO481rmuMUv74ji+kpJ61QF
noif6pWg7EHT0wETAB/wpsMK5B9yE5Vyh/jlKM2V+nt/7n8VaSaS8wAt601LETwT
nBbcKtKiriFtvm/IJFwjZJmFASta10o9fIgp2t9QSTi6Yq50jmgdQ+eqJPf7kpxh
M/HOPZbBhhT/KzV5pPZH/kTSBtXE0w38vQwDwdTFX83Es/+E7msIrixOtRQsoZhN
Wptetcx0QqSefitZdj4usmWiCUOWN7AyPQytGoaotEeopBtcO7077eEyr8Al5fxK
tPUTDX7G8UMe/y8qY1sM0WXm3Zni9WB08hGTxlppfNOszsNNT/V+DFdWDxpwvEQk
SW8psHKDmCIHm1oynn59HYaBoi6/b+unIA/q3HiJusDFvuJ6iyrBa4I5s6X2Q9/C
IVtETGZmONghnbLcCHtCo85caqpZVwtgAR+xoUipnT82y30rUdjoHiuVvhv1xS4E
FUhgJE4DZ+p2UaGPOj3WN3pDT1F3mBX0vUBeR7Y1kTN9YylQQq2Bt64CfoRubf0q
EoGu5MLuIWw6AIK0vvKWIkHHtB2Pf2rTINg6OGlUHC/Pcq1NYLFeVzSLEQD58T8x
H40y5l9HeBvEwM7vH52/CfF292dhqqMV0snTv4S4mNGfhLsRrQpXFWjMmNSxgqLK
XxTm612JI48aP91g4RV4sehR4YmsIXYMS21W5ybe3oQjYAYpD+gPzqjmEUKMLq9o
8cl5vqpMvY99wPbQ/uQD9fCNZebUUaghOIc07bVt6FQmgZ8lPQ1w0E4ZIKcWTjGC
/1rjteqZA9c6xLH/vo8rfeKDCOfc5RRbxZGE4RBLJwNK0U6e8aeowieue7mbQwCj
/LGlHGNtMnR7o7Ypz+qHXHlj0Ol6Zwg+uJxxxi/anEKiC/uhPdGZo4HngBo7Uhuh
ZOWDs1QKuOl2XvKQTIoyMq7It0a8eV7ov55ma6zN+OrVNy9sisHlFoN3W0M5pRkb
VFfZ0bdbkhaVeMLkmn3r6Y/hdWkkREiC0untk5hVlpkaNu8QNrbfpKzQ0uSwRnHk
wt/V8GKn1tIjTpO8xTC0XtvpGVJPbBCIPPqRCwgpsfhsf7Zu+jHWlBR8nIggiefa
BFi4Hqm1FZrvII5bxr+0kg/lSr3QxCsgJix1ybod41dWI0hwEJXBaKykEmpWoa/h
uRwmaoAY5CCOZDTavJ5KXllqIzGu1zAK5eBMHe50kkG5NKhUXCdYLTOzlmsbS29G
C2+BI/6zLm0YiIIndnsLI8eNuguXSgv36GJZzO4Y4TdruclQHeYbjLV2ICmwJ4aB
uwsJICfkfWCRbuOs+rL884FS+sCCkHkyaZxJQofeOD3XPEOglvf5BTZSwrCEQmsE
M9GS8ecbdlVR+SHgbbU+KWiZVqDakqDMBfXrA2Ugjr/Fala0e4NhJSapK0gIIV1V
0ToUDzG3+EnZmvglyM5qH3q6A6FIDgcKsDrYDWiXrOcaLtmMx8qJvQZlNkIqqxeo
3g4tlR9eAv3vYk1FTPApqCYHkzfhxzXys8yIfJQWXXHNf/qzt0aknj83vx/xztp6
ljni+m/RQ7Eeo8lM1rNI6PqtecxOS14uChyLo6LVkaaki6iFNE9MddCWm+wKOQep
36qQpVAXlRfKrsmtp6PNA9l+wRPgF46YEQg5QjCX+EEiCYsyjvhvtwZ++pVSzAyJ
keGKGSbNYGL4gjxmIlWS7fw30buFIUyqwvQvEMUz4O4tk7LMbD3+5oqyROthqeyQ
hkEHEBk/0U+yGeF0TxUA/Tw+cI13+9dJ25O0UkCLyWhFzfse88l0eq2ExP1S0iU0
EUDo5oFt+XY8uRBMVtrDQ8DWapE/CrhTpPJfXMtx9e8kveQecxi3tSTMOMFIDLnU
c5ZMydGCqJ+LPfl2f9FmgBD58lz7TI3cWHdvMfDgrI06w2lC1aDV3/57u30alJ+8
FsabRk4K26m8O++ucrYLBoOy1JRHU02aFnC5wroA6BZTJuBonLFKe+JwKIeUjMD6
nZvpl3LwW49vWVephkFVfAtXIhY5EomMmWjV8Bkg/Hh67TvOtBU+1kD/91TUq0Lx
UrbakzVwF0/JvLEDTsEUBPhxvw+aBU88qbcgCDbqHRutjfg1L13HCTUCBmf3gQWf
Jor3MiurAKNwXkHGn5cOXqx30vFJ28bJHoG1dRbNxaUtthmrUBJV7y/THLkhGR+H
OcaXZrt+SfHMu2AQ7cuFUxDIT9QT4TgdnU83dMG6hRkWRsNZAKZYwRRvcYqunbUT
9vCEcprFXs3Bkjq6LhZdRljMg3B1cGcCVxs+XuFJXbpGJXCL2v97NRioBx9w2Gex
1b5SLdDCOCjUCaxarWw7gqe5bxE/z6Ee3ugrgk/6oN05aW9xI6/n/tU6qWTc2/B2
TLwbQWugSKZ5gQr9MKRHZ7oA0cPRcWOraQzZd9EyNEUMfTHJy4A+MtCR6G3dBhJk
dP/UCJnKpnMNHbktLgvnjPN2D8NEbXGaaCOixkCbN5P0DU4AyTR4LAnqY4XiFUzJ
d3WCqxd1M+eRdrA6No1wzybuWM4lFbDLwd9VQdolgFadDCRh9yLv2EVuJMtqYx0I
gsx7/d58BopbHQz3Iq3Pfs+QINZW0LORcFSbRuiavPW4ZjveHSwc9sFqoLLlnwEp
8KIH+y8U74C4Z1D9MzBviE4EsZx/VkLyVBwVmGP8mi0nem6a2FGO8WsTAB+0n0Zp
voB4L8JuMANLytWvLRYrZtqOhrgvw8J/xHftQJ9iu3uMl9qhwSR8Ng4f4cy+H7V+
5c0powiMKV7yhS0inWxPhmR6oWUaO4+IhHoY+EC+D5itayIafy4xOBW2grwHQYU7
6EQD1dZrQJkTUXE17rHJsmHPXmzHRynkbB0ftTIQg2hqcZB4hj3vX4JOLXeNjg5r
7ijdTTJNYfNYtegILvdepFqqKR/ll8lOJNv+QfznEj27siBWEGoMZTxMuOdDYoCG
yXi48F0eqi3TxyNP7JbZ0RMWydnXXkWMWrKJ9rxPC9A5owDiNCNWxLs0j8BIaAVD
aQxSU2fO168JCBdy02E+QgyjGoSgGyujmUK283YTk5nJdR428x3G10ZZ6ShaheF6
ZXFILqcOhCoeRu/cNEUtNQJPidpEwkUTS1Z9ENGHb62Dvlyic1vzP0/rGLoAeZrO
AIgM40pIClCoRdybIKyFyvXkczDHDehXaiSf+G+BZR3IF9XNSbChzL5i56SHc7sl
XfSY7gosZXw/WtQFqHpqksNvl6ychua9dLM5Nvp8Jxiz84XUrmJ7k5xI1f8tPPHM
8aC428XWV2EfyMd1vw/fRazXjn/AK8aatue6tLGYRTT4yb4bO1GSsmtNyRebdujB
ZEk/v/n7lt0hMWlORiqADRkkWrwWk4DBJHzDQJiGyTub+wU3tLb71cEl1hao2UMs
EQc1f/TepUuz/f07MevoYv0SVKAhJ5lgks6JoCQ2SfU9W+zr+Y066mpJ/DsVZYUE
kZ//zALrvuRXBi8XPxICmvZ0HYGqySv+/H+lGUa6lfhkuXlM4o/wOwnDzQJOIbHi
iKcbW+RpaoMAmeBWy5hNVqsANCCP3cVRxU3WatDKgPQLu8xcrmCMNAxhHAt5Z8oD
NeLtzHxZztIoNPn8qY7aGsrruKLP49yOtX7wuocIJ/rYcHdzc8ag1nwXvJqEQerM
ILkgDPz+4+WcNb9VkJM/5w4uzdJl4UOWjUdfWteURNhdc1thwB01roeETtuKAhsm
Gblu9V3BLS95bMWEOlgouuFag9b1051o2KYLF1UpQZbnO4nftknK0pPQjXMOFT8+
PqiIOrJM95MeTuABDBPJwrMNh8Eu1Plol4mxbeDQcE7HUobh1kwUN6HmEtEwyuLf
ZOyCt6foe6Mif+diGvdFAN8kXkLwLqhe+w1H9fGUKODyCbY9JsRRsJs4Oy5Hx/j2
/Swwjld27ITppeuc6xSXRjOhYtEJP6Pp9PUwu2Lq4WXytB1/te0lYo9JniVbLPU7
lY0qFGtK3gJ/HRSlXpqu7BCrU7/u8/DAELYNthM0P79GihrCQlNYTB0N4yW28UbS
Wyt62ptlm8Y58MIKw78Q9XNDrPLvREl6bOqBlwpvPZoa4hGgVC5ua3qRJ7xfw7ld
wvhCzrzxWBTjyoCPWb8hDU477I0TIACDZPrxe9WBuw5y+OcrOGWD1dKMiNpTjsai
1adf1HSrsKgmYzHbAg3XeLz2YTeQ1dadbkJxHSFwoAcRCgTBtVm1Et6CLFwwXh+w
t30wF8G1ITXiGYtMhLEYzrrBn8EKWV3Gt15nCrCrrSlPS74xwnFf2h/ChES9fz1h
585gpsbtkZlGDhom/eA7JOU6MIHU0SGDEMvu6Y0AGBWE4lnkGEbq5+z/mAUZ6BaP
YXTem3cf4mxuRRCfGrfY9wf1LuwY0s9FiQo1qEjD0l5LxpSIbNFGNiZbll0u7dY9
yTQLM8wnynNZ0XZV1X25JHng+RJnQvAULgNm3L4l8XnPZb6ZnRnM04pXAJkJXMBX
IGed1t/jALWZFlOOdlSgdtLyQ7r34jshva+TJ2/MW3ohw+E24LslTyPeva4t6g7k
W//iaexkLpr0k5Lfnde9JqKd68DOzbkbVItWC0lFtRfxse7p2cQOkWnkoUkuFOow
7UrMtkwVP+swSeK2d9ji2NejePG9sbYXsL8+k+HYdrKBYo7O2zfuEhAVN+wEdo7T
e89QM+WZX2WmHHS6bwvDYguVI8zI/3eEC8hcPZRjEm12GxR+JuTnMfA9/jqCsjXj
7h7VMu/geuE6nOgmQUtiaqNKFVVO9RMMVPZnf4kVvVmMQ/cy0IEcXCyPXWslZr1j
aRWdpy/zLvZu6QRidXA4fRdfQNAAeWIKUj0AyQ+US4DPMZLGBX0z2wfFM421csn/
ZJjdBOvOfH/ng31LAP6hOcKurMmi18Ro7rDcRfb9A/hcDZh9IVdRbCYz8S6CJOtq
32mOnMyuhCu7oSykXE6u/gRmNdIwOrefnsA9poI/Czb5cSgVnQQadouC+MUnn4so
HA3KZPhygcNWvdh45OrSmF/EqJZKShOU3g/2PCSy++A7uLAF4QFNPETC+yUhtcA3
DotLmTfo0ucC6QPGSSa1nNeghCoXSWwo/Eo4gBlMVd+YYlmOT5ylTKbxrWpxhcne
fD1zYySR+BEKQNP4G9X9cCSZnduIdVcGh96gEWxdHSt3pBznjK0+mO3xNFgight4
eIJVR3G8MSFkiOZGOay+qgWd4mZqIS9boddOkgvmD1XxYU8FRaKGuWHUP2txr6Ot
mrPxG3RlvTFq8zTE+4jmUy8n00UrLiBIRQDrLpo1IF11ttpBwW8vfwIz+3cR3vFt
lU6UttukUzW+uvsDAzy7Z+P2B4uamZIrEsUhiBRrlUZlUTNT1OFOKgUrRsWt5XA8
TMY5YHRkPrNsamBBNRXeISPEZEYOemDYKbEe1So9yOa7fMnYVSY+Q2Ftb1BFuXHb
cPQTbzJNKKFHhRbzJzGSnDn9sJgtTFCAaDFtT7G3MRgBq5LZBB5STZDeThXmxrW+
iHyvdJN3pjW3qWqcU4YF0ZnRkRSOiSRyR+d4N8ua7qA3UhG5vnhRVWNggOzC0BdX
fhAs1kFOtPwZu6np8lrt6oKblvDKkE9uhNdieSv3lxWIOhz6l1/hspxrMQ5QB8mj
Zsvx2ef5Hdp9vtgxRvg8/STdh/xOb4tA5EfQK7ReLEfrpbes9zi57aedJQEZcbI4
guEjcDKQjAipn8jc+IgB3EOzAKlNnYkBGrWEwIKd02dhLlIUic9aiaD+4yue+N1n
pJf2VAFfDCzHRVFnU2DgMOlxt8Cz8oq0e2ws+zutC2pjksvYBeRO7eoKweeg4y4m
ZklM9pZpKCJLd2/KwfZ78xRHYTlk5/2yKWLSTI2dMrTIFtbhSYj0kUrpJPUjUYKo
YqnONnqYtAFS6vDEMo4G9EHnQPllvbwss1a9wnjWU9FBWqyOppzk2Ua6q/Xo9IR9
WnOgfiuHEyQUCZKaVAtpGuFJ+fCGMfIjZ5joPAsUZThWeP5F9TKGyNMNRjDB2gkB
m5oEz5lG36SDXC3e72D7boa3dPuG9tmy9O2BdYkNqtDqEuBqatMZf+tNtB6I52u1
Kt6ptzzXNBFt2PvFtT6/VkRQvKiHGfOuDGwHhSgEzDl7gH9TFip1bRObBA+/umdB
s05fAvZ8tKwsglBBzdrHQIw7b5uT072dvyu8JzwrELQmbRGkxU40KWi7ZDVwDT/r
TtDOtkFFaVl3M8KfyFaJNZzgzgqIKAAqAWxdHBKKH2QXagLJMlIdlDGbsN63hhkM
9FbBBCBtfMQbB7+Pvp2nkoKgFBlNip5hcaSOMVIHLd8nz/AFsw0cXUFMyBaoiRnz
zy3ZwrCaPud7G73Ik8vwpU+5UKRYROPr+KiVE/O+2wLX+6EQ9ngwsLGlIc7bwaxV
zm90f7eUZV6GKc2sA+9gh+MRo12NESvE6yPaSg4gYtcExgbgkJqpss8qijAhmyPC
VTJQe4Y5zinuiTj/0doMSDcbIsxQeXcxEeDsjtfK5x83MQ3x5fqjvafejOCa6Nd+
Uitw9s19pQW93cr7tOvXJ1xzKlStbfir9L7YbmfI5lbFyfimk1oPxBrKR+Z1dMzj
y9PD9q1FTQ6o8C4uLQyiJnPFK8rloilkUXzT2Co7WjDBU6XNzB/FqGRhy6Me5y3I
PZEPKLacZsw9OcExSqLrnl8s4xdPKN9O7OExOeUufIc9ihOfpKswwUfgS6BeGLUc
hhnodauXLU/BmD/4SlH91gVKbeR5kCKegz7UoR4DeR2KpB+YT1Gg5N2OhlEDX1v6
xZslueZikxjHLldZm4qdzUV5K7EItjuqlHdjJdEIOG7nNEgIk6I4go+1DvQjiZ1h
fGHp5PUYVTvO7M7IyXscIEMkDjd7mzs/s7XABzn4FouXJCTHoEtFCwMVXlo3q7vL
9NFNX338B6vzXVNbXX2D0eM82w9GPIXYr6xkyV9u4dpat/trgfklrIRxkC6dYXqM
Cpi2Ijtbs5hUtYz/Y5rAzU2KVICbrMR60WHg8lzMwSkovPBEln0/ki73U3816DMA
tfcsZQlrGFqqYYAK248LHQIrwtTWppil6feH4ReBNrKtLJkebCSexl3e4u5EQvdd
Et1+St35SbOK9BWvyn35FwfAZX3TXN2ZkvjTyskVPB5lT/q5SVNpGc2lZuJJycRl
8ZsJGkiF4pZw1HuDl8lG9SDBLMrNErIf2Azo5Ip7Mm5L5Hq+xFHDylfygrzEioR+
xlZPT/kTvo+YhUYu+9xTUeRWZ2L+6WEcKrKQuy2HkDNHW1rneEyjXrKx4QLL60ow
qVXrvbGUMO6QvM6uxrMeR+c93WDagyXnCoGrzz6qzDDscGr+NEdicjPQgx7KTixC
ML6RC/e9YiV3vc/8U1K0N4a9bVRhG2n/HAzR5+Au6nWybxacMfjALnzMZCBvYDzI
alh9dg005/ChIt+ZkBFV3LrLdx1Pli6yB9ToyHZfvRHpIO9qkgaD6AFRN8vcVGh9
kxBqzB+U2k8xA73T+OVohHQxFJKbaMrnQP2rfRx7risXitiw0wfjH/7iuKUxBmoX
QwwfLJnYtp+Nt71WK6e2CoQAl6sfVdvnWAvUolqRRpy0ucYsVfRlFB+RdXQqherp
wtZzxmxhYwH1CH13NMFcqaztwgG2myfRgJDKg8PVt++O3eMo53BY+RFu3XZnAhTq
76aODoG1OLKsC5390UQf5IzUUeYwZUe8ZQkJCrtueDCSrFS34dOLTWg4asKIqcGA
N7B0e4bzRu3rMjiMg5GvspM/wT1UF0/iCx1GHhmU6gvsJgH03xIaoviFh2bAfr6R
8AwkWqyxeJdPbl1V8+3X5QxootKkIrTEyx8zjvAi0y5/maubNKuPw1KdG0nkbjlq
ClKKY94kGk1VSb0YrQMR38jCRHb4jiVdHzQ9/44DAQFJKOvYAndJyaqgAGhnrLC1
7wEewz8x9h2XPfUvNyHHxgkpbwHjMpfRNSOnTeoi6Z2kY8RaAcle5HUCoWNHBPT1
K0I3uOqV6wP+rp3tU5sEf3vDzAWOqro8PZ3DQbzJqzs0fXkPkaEddDNYX92b32U4
YaXPLrEogaN/Uw9LCDZCWsldksyrHPf5VEeo6fSod1BYkwiKfoFlUaG1C2k8IQDl
+byyXNzF6rNUPTDx4dNy4R9NuhISdTxsLiEGzJX3JQ/2WDFL08BpWK1q39C0Lufz
DvXvzmB9Jvplfjbo1UHTV0oorCtSvzlngpZZYri237K7V0pf0VQM46mvuj4ogqt2
g/khXTmb8gm8i1Kv9ZUZa9F/OyzeBVQHosQyNTeD/A2YDvwxUVWfEWVXKvIqxlC3
lZCFgjGKR5b6TyGLxVuLRQt39BEE0fNWqcCbiEI8OzkEAudfEaYXvFEShs2AVFEe
6PUqJ7UbKknHzutDTYVAwyIAAC70VG/3pzbPT1fAyYKhjwOPrVvfe/xlI7Gqg6BP
/deNBqBqYkc8CQNIhvhaz1QSsinbAxMtsFqwGy95ZysEeZlntFN42GhkVRT7yL03
O+TVRPWS3BONMY5lYKrHRojzgHE4SJowbYbkmEmjD+gkGuoLkoOydG2ABbu6BiuY
LrFXYs0PTrybpgsEjagYtDTfzCYYTUyoAqTnSyz3Ypv0u9f0n9NUtlAcpR7BcWnd
5cjLoEdc/Lq/LX1+y6KZ2j9aYe2BFwHnSoolgMnqvmY3pXRxtbvU3ZGaXYLgUrKs
dDHfBDcsUda3phgdI2y7Cbc+UDno2QMWQaprQShn9f68FBRiwfKLqRmz+SAe7T70
sBkvb18Mgypza8xHjbw0IhjBdlG+FN5ZCoEsvfe06op8yR8+GuxiZNvtsAE7Einh
05vTGNhZ2TsWWn6DDI6xHSgmXpxRY5DntqpyftufUwin2jAXZlhern1MNrTqbGsu
fNVguHjlFdXkKD1OWTkbV6uoTbb3XfJfCMUHRC5fNmx2ePghSwyppQ0fTshPsoeq
YTpfE4Z9GPJyjYORsFzaGR0vKE6IYUAd6ap0gCv3NdZbHWzEK+ZsysVQjhcEYC/e
tqhnRIuf+Sp8wWxnpaW9Rpd11ViL90tyAFORLSJLa8LgWuzpVNqG2yWB9YrABoAy
0uERDrBTrS8KMZ9TCOKa+pIDMpR51UonZ6AVICyVNkPwYFz9YR9y3R7CMRRF1u9y
L+7zO4OPggIjdqUueJfNvNHuwwJ20qYA+oomIJ9ctZkOy3dIjgPc0Kw/iHN1L54x
2XXzc4DsWqwnm+ewEcJIdKnwzgqJ40bXp9hILU4IiJf1jLAYZ/uQhFgTeR9errsk
64MOqs9PB6Q6q0rgo8wISYQKlyhM+S4fXWLVZg4qMT695hRdPKvjYCYbmSS3z/Cw
Ncw6Pe9Tr3N4oggRsDl+lIfjZqTypeqkex6FwgnFv5Wml5FwnucvnQepiMmrqONC
bglSQYGUPpFVz3EB8wPhUFKLkanO/+3fPHbyVyjQrX1rtihJq5XP6w8joG2JbEFF
XHlJai+oFEAAEjCNOF9pZgfAUiMijRLH0FSY+0q8jko7C3ABZz9zfpf49YSnzC7C
gwBTMXlFLQCLGm1Qg1KC//+pkq0qFCQZyhuwejP+6bvJCq1/Bk1YZRff7O9HdPDB
1z7H/AKNZ7VpfranKCIJ7o0Pj4r1Y3nyIrHAFKncdNj6/97xrUuHhafnvNM0MHof
acNd9oUlii/E3ssYpD/vvguRNCZwQINsMv64/x/2Ts/EvOUxDNMV3r+awfclq4Xp
bUarX7PuzEYk6J6j05u2dz2ZNNS5zu8qm0BB/3JBXUdrcizeazgmoIWrMPhoslp9
ajNTsMasMobiIr46skoklJBddGtIYRCJQWacHToSD/iWvVBwDrpGXbM3U22KYGoD
XXhOFOYQK9Vb6kUD+1T0WqK3jT3wLQ6TgBK2sM8pcCQb/e04pNyhh4YLMxfxbX04
kcf7wP85ufnbYKBzi7lJrJYouLIfKGNQJTb4eYOH/DSevy4P2Wi/q+8m1WG0Wd2u
MODJ81ZZbIgM+a/r44oqn7iCKf0ugIgDho5aeo04RNpO5cCwlL2/dwL+3p9+Ys/B
gX9oBWv+cjjQyEN97WUBRqY3PhaXLZCzyL5EDDzp3IOQAjvvLoYL3PNywKNMIJae
Fw7+7J8acZbjV/XM3I1cQSobd2fHY6aOB18slRIpXOZcXPLr6rtf7kVbAxvLDoR7
bVenStCa6vvbBtbabNGBVWIacaFLf6WXz2vlNVnqKpuAEdvHtHc5Zr9ioO3cAi1z
U8YtupQzD/VPnLpZ5+d5Own4rPtI1Z8oV1t8EQe/SRuIT8+C04C6v6Pro5bfyonx
kH4YGd/ridswU0qIkWD+8qimVd+kgJqQTc2z6dgiLo72SriKDx9Fp2l7kJtYXJei
SaTm2k2ffy9zROfnE1SLXnHtrt6o+DE5mZ581T6QvLe7/3Ex7ho45BK850c7AoyH
f5cmF0Z7hmtdDoWXJfBh8ozB/Ky1o9uNokMxP6h1guirpD0TGZC5XXETDraMGRgo
ZA+KlK8PTKB5wlnsX2PIM5Jx/i3PhqBmi3yyK7GCUkCOPS/Bd7VLvD1mwNXW3Lqh
3VVeJ81pm7ghrVC507pS6k0ilWIQwHawJK5xpY0Rm+8gOZYSDL7ypvdKtYIdi+oy
IsoR1o/ZT6rUOtUU7mqkr4+eT60Bze7z25ZXHZA+yjRM6OAmShixQN+Vj0X56msS
MUo68QfVsjNcCVAa6OemTFOP8mHGCv7wUkWLYMjD+qdjUkfzkHJqALK6pUtLPkC9
ozSnqaZaJZguWoW2FJD2hFmO/EomlN7LCvp4sEvTNYTGKnhmklmFUZDVTEuw5IfZ
o4cRDhsbe3ovSTiUUbnKJ8OZJwly+n3aI763K1XH6V7HyDnriH2fkK25aphzyu8s
c0zvAFzwe/l/OlHJuZjkal+x6Cz7QgxUCK+qa84vZrFEFdJOkBDtjqEo6W05f+3F
3PYh9bz72z1PySOlgMfnRJgEx9nu4BwlPPXBup0HIa6VCEwGsPk6ElWg9eUtLFB/
Zz4V/SifSw449bT3V34Ho1coshIzAzxaG0xRymt1cswAJterX4HnxHKaZqveF2le
3mMZikMH1buXWpHfR5tpKLF313bkDkXQ1sZC9exSAAix0w/S+sLhXpsOORK++VXG
xSHGREfeAXgjoZfwoGhH4yAqy4viDwR3JOlNHjJ82FpImvT7cDuOJ7mS23FhUSBN
a1F873lVzEEsyxghuD98qRAPp/Tkc5HRSe/FRLs3Tey/q7J9LqkNqcg3Hdfs8Piw
loE2RwhjtOfV/zT/E22j76XuumrTDDoVpliTPtflMUzo4UifD7CbowdfKQOLDpvh
UttlZZ9AeBraS/FTO5Murx8PxEqLFNROyf5iZsc1qQhInH+TDuVaQ+IT/zxm5kO0
iHIcJfdP7UMuUpppZ1UlqopqQTyRPOcvVFKokeVFVbckFw/jrdArZv179BwhlttM
5lkWBd9YQtsbnYeNPMhF95F7/zl3aVPkay2eOb4pKCVDFcMLk5o4bjFzchJqkXUB
MHIGBUBwzowgXtlyU5YuYcQ+Eqw9X4+Q/tHk9xs4mVakSQNQ2CBqKlS4y+vszD4q
0Dsws87gn1C1hHezwKH5ZuJXwcLuDEBJgKfrRpVceG0cqFoybY6mMe0btCAgaxEN
ReWuJIN35HflgnB/nRpZxSlDqLkhqE4S/BHG7UkkIHDmQxb4zwuSLJg/FdDtU/OR
MjHobU/aFAc7HJ/G1DoW7jofIglvZPutsv0xQGVGlojsmPDzqm5b6EJh0duTI1z9
YF4fzk79gGPqJiRZgWDKaCgKScrQwf91PvuM/FQQNg/6MXaMzzZVMPKP8D1qp0NS
+JU2Y/4pefXMu9A8YsDB2bJ8z5G2ZpIyT+tivdSQZ0amfrIG+ECsYnKMM3Uo/kfq
HoLOigXIW9Jhq08U8+IsNghPYWwuJiNCtSgiAB0FVi5+4FrPfQL4rl1Pd4vof1ZX
YBnP0EG5vwQaiOa+luoUWFMGeuUVNEanxCF5NINoIX4w83wt4W62DL1c5hAnvQLj
NrvVBGFc/VKlW9xc+1RcmuD5UZ4oN7ouAQN6eFjnn9ofeYRuqaOkkcmJAKPMe2mz
DZtovWfc6cJsqsb+i17CnQJMEbOiTk6qJjhghBJ4H0FC/kArUcfcGu6nY1bdYywc
nmfvBAo/m9qxNqUkp66okuaIoPKpk73z3MxvwrhHpY3+YMLCywlQJOLZM1ulVQWy
Fg4o6EedeaD1XPrSId/H6c1QxxO8PN5IzAAj50geRv1wi6eIEe6YfdzIlljfVIRc
1eStMnp4RGubdh1xsNfeqpTxMyHeIdp79qVYe12eHoFKMbujbZz23fSFVNROxoDH
k2rxEfJmjW+bjszaIlGloDM596tqnVAe6P5wpyMVLwLS5Gl6uOHZsgmZDGC5Bmpy
GgbGzDnOGvGWdkq8NoPnV+ROUyQwJ3wlDBY45FxfrI/ql7/wHEvEiS1k7TGvgjc8
sOBDdg5XRQ5DPVOYmjiYOeHGpcz7FBoRZuCHcX7RTeBZIqquipXk2s1uAFzbuwPW
3MNjast6yxRrk5AfoDMLbq+6ljwCfIK3ECjofAFSAtq3PuNFeCVnkMQBhRmh0sWd
O2YwIq1YzQqL4yxGPaxigOaSwFwiNqO8Fc/NdsXWjB+M5KS87NyzlakLJ4LEqre2
7tf2tLFPogGT9C+XkUexsOCVrY9HY5rMvDSrX327YFEDF4PAJkRho0SzoHZ+sWy4
CHaWuBMv0BeNh+46xxnUp2pKwRkDb4vVhg9ySAc4XShwVWsztDjNFaRK9RrTst5M
ncOWjbfq9tnQ9+aRYSSONt+94fOqOcuRrDGV002eCsQ9g441T/vcvl1++WqrHQAF
pZ6dfpgMWPwTh9+hPdLOl86pQ1NBBGA2qY9WB+AJ1Np14qbWX9ASX4FHN+gnUxtz
x8nZy0Nk116rpvAfo9WcEYyUMCUd1hUDwCvWQWlnVE6BvoDSLJSsaIm+7KdU43t0
uHUkKZaj8x7QjfCC1KaxDReFPtNDUh6uxLkCcttz+vlHr+IF5OeuAyW4303cmlJt
Nyxp0Zb1O2WPtFLbH3tkNQB8SF5KLPuEwmzCyIWsPcQq16foiuU0XodefODt2GRT
7jSgY6fd2w8nv0oPJejPT8aWEvY9tzYI7u5TmAgPdHd88AceSD4W+0n8P1y4Gz9t
PvP8nB9uvofU9H229AH0HKK+x2b75uyDyJNxHpJBf8lPENyoMKjuI9CRmv7zCQ1k
ppFpGlxuFtRoSgL6Jmdw4rYemC0FHeZ2uYV/jqbyKNEGnfIVx2Zko9YMyr//n7xV
10CEmbDAqb9sAHCzXg3iP3UTOznD7E+FJDIxmOwq9MYtls5H5wuE32SbwDkLEtFH
HLi77Cp+Y0c0WP/tDAm4sFRzJKcIHKnXdWpygSU7tl2J5o9lMTlruWfqS/elkykX
rIvpRP+WsnV9asFoeIlket2cgOBQNXpvwF30P8aDOKX00AxUxVO8U+EgvAuVYRCI
IJXoZJKh46Ml1ZNoMeugJqfO1KBnJ3V73b3ZIm1aYAsOEGfpRbU1CRfSHQlTd5JI
g6u+QUNvU+nGr5UOt1fYt6wUaI2ykEvFXDnOFKBgzN6s3f030cMXHjMVSZ4cLQ8P
YLaljV3BExwYQdSzquuUrbOx0CXyGcv5Ga6Nu6J7D60t6cL6MywTfRwB0WHITQMQ
0I+DuCwfzKdI6ofeVkKPBNjmr2MitI1VMHD0fN3gelkQAn3SXppM+7N1+Mc/MnXy
lAOQmuTQ5RJcdgeEFar3hj9APBN3UhEyZIy4D06SacsGBU1opLRtsFkLSmlfZ/93
cwxszok7Kyx8NWFqOQSYblvDoIjz8slWL9GlbnMlbrT8N5xCbDeN4qqvmtwhSXYH
et7ClXbSH+kyahgoT1DSqq0PsoiMMXLNRc0WUNAkTCOC8A0d/UUsY+VTmxanxMuM
rkSVaYl/f733IZP4uNMOCIaOB9R91iUPTPcXys3C0uZPxL41fnkKgiT/X54//JJ+
mRTesHowOgPl4gmunwUHtaIeFF0BX5E3yT3zvdLSJp6RQXcS9bQ6HM1iA8h5jP5W
gaxgwRMCRQtFbqagVQpp+MmxY7I49GEf9adOcF51bfxZ6RredtZANSHPDFY1vqj6
CU5eQE5C34yqB/DdlvStsQNON8PuxUsUuFHyg5yFt9nmGjM6e+pXIa4GkVF8EyiC
bLG4gFukf7I0WwNT3qD+oKlVGFHRob1QCcyfxfOxv3RhDLdvo99id2SciQW8u2qG
N39MepaURw+J6kcqjYXMcin5v051dSw1VSNuWe3tgfqZa3LzruBd5IXL5rlb9QpH
HYjUtJjK2T0mKYeALnP37eMA5y97KOGqgLNMP3NBukUcGp0gjE9/sDGPmNPggx62
z91hAL2cenfwdlRrJcnruAemfK8xLtgEjrgVzXsHtJYKSbsQl48PoiYcXXQJwLWw
O1A9HrpDsINQ/s+oPP+0yixId49pfrOfP7LVqT7d1o81se0fNiD8zKo4S35lP217
/eY26x4LUOBTENRWHGJYP6unCIWbZHCceKaHgOjPd8Xowm8NfJ1d5623PPDIE4ns
r3DUWRZUg0L7beVaYMDxC6G4YzvVW8VOuBZoEuuJXfgxkr6NKrmeVy3qA8Pq39tD
tZWRXB10LrX6NAqgbqFoALvqIBiqS41+llAKscjzGg50LnGDCSdLGFQEVTkyILco
chC7XfeL5azFXYLRYWFnuLRjFjl1sOGaWgh4bs7Hbmpo9fa6f0AZdNUEIC6Cmorf
nnk4toqVYXCNBQORTS/sHPUFZ2m1MlppCWtmu9/m2qkv7Zs2oSFEiZokaycgEXN/
lmdqy3vrfleR9wbvXpbT/nR3maTWJClMdZIDGG2tZyJBgmtOBV4X+QpElh+m1p+G
n5mXbt7fxf6xDeM36TWRmuWki2gCjUB08vo9uyL5ZfOsr5oNPJV/C+LoWQX/1pF6
7Q2AzyQIEEkiTBEfj6F9JyW33m1v9FzXxLsWcpYot8q1HKlCgr0Tjf19pqoqWf3N
9HDhSjP/NAz+/BhLsbNe9NXkfHlzAJ0PCYYGHut9Z8WoZLqMnxe1UcFQtVAbjvUq
8bGTf25dD5WBD9lh6LU7QC7J1r4HjWqCybKZ0DPwINl3zjwE8W2NrHSYGEVBB/81
Cp8Qk0+8dPCFodhSbl52ofbLmYTtnM+TvC2F5fVVp4Ec6aNT/bmFHuhVmYBNxA2o
U5cO48enFrOAQgSD9y32t6pj27+gQCfVU1QOqdNBvw0saG45yqqvxMc4I3p5kwII
pG49g0GkfzWmleITRkbDNepZ38F/pHl5ghUGTF+wTHOJkO9jIRgUajS07stYeHjL
0E+x/86rExKKrNAY8VH+tmGrMB4WVfTHPSMLcB9TdJ7wjiXCbnOn6OmiyKMqIh6k
2Gbn0rbnb5oF8DAuD6TsvOTzZYm01XwEv0uSCxOmCAXKrZOt+n8Hx5gvjWEKnFLx
VjE3EN+Dn0jIBj3F4Pm1PFI4Pqy6Rl2sKnEMuz7y+1akzrR7KYRv5Ntn57LaM5Rx
lGIs+YO6EbL4gurdBfCikwb1t5IIg1ndv1tiJkmaKuzAS6yxLekY16hf6DoC+v0E
cDbCuyVQGz0mbhaG+Y6qjEzwwqDV5ctV/2LkYvlmhdQSB3AT+KQ6O9du94coEOoV
AzKGZ22gFoKlDqw47yQ/6chHwIDmHxHxfUdbYZMzFzqtTyGFPCPhNy65oG+2EzRx
a1sx7msC1sq5lhfW6QfbFEZkvydU98KL7gLkRC3cI73JYuSK6vTfHcIp/UG3Gb1a
cXTdGboSrHZmMzQ/pzzeqv8Lyrpq7wogwD0FRxN6s46BLrMYYTAejR1zU2x9FkUl
4MHTLKpQf4d6TcZCDGoXvP3OZVuHcbkXGXkjGe8qYMMWidCpE5122Xh/DmG/j8LX
HExFIgfYZKtczXhbyNgbYDVEtHwZX8tYpw2XxIrawng5bgi1oGORRP++zZEA5gq5
1wmdV54KgIX1TjYGbXBejybRLsp66TB/WHdOSQmoeG8Sp70z7JwRqWoJ8ix2cW+I
yN8Pbmwkz4m2Plv0nVgD6P9vOR6NH01cYcBNQC8SNNq1WzEJoS/x6KffumO4l+kc
KEiVzkOIwOcAiO5KQddgCUKL23bdo36OAmFFOXp6zJVuzrBWF6+atc4a4xZE+oug
dA8pzhRlV9v5UujbxWAyqFOHuXdLx/UVQJY1JYGoJb6UWMAh+/UabP31s51felmN
SV53E0WlIl55V1tIoeLOHeNM0VaHICKmgCO/rYZmsQsaevWkPtuNFUQkYY3THe0n
Czt7LOdMKXA3yD8hIr8dkNAEO+I8xIm0yATTcTiUamxNG6dxm3ohNS/ltAvsolh1
ogqJEFYYQjY14rISZjGDnqLiqWy6k1cwzWWeBqLQkpXrJQvbkXBjiwRadzlzVBqe
eN7nwo2qHyyc3RtHO1tV2vVnoll8qT6EIaSg6R0gv4XCsbOdQwSNJeOiSCqTX+wI
i303Hm4tZ0OymcIJyjRUImhejjeesLPreJiVNv8Vhc/WJVLLY0y4pWbVT48xiIwx
51TbX3dM/TE9ov0twVCpkRzFNc+Fb/xU8SuC0NElNsP4O2IEkcPA1XZvE+gUImtS
/Ml4jcDIkZO+MXveAzJh3DxOIxcDdE3c4cIRsPc6mgcoOtooJvB70G67HKxJEDJ+
aVYyR0stUSfS7UVDM42tm8n3ctwHpTQjjntPWK5T1llkHeH56yYZo/ifU2i57sPd
8jXFVL27o9JV9ZUg0BwmcJdAQkDr8usI4JGIAivsnn6H316BZQ+4F8VKnODMrlld
0Krz4N5BPACxGVg8bQDW9Ug/auxNrhF8wDzcHUiwHM9z7LO0MJk7qghanaEGMWr7
YEVc8J22kp20U/nDVgQd2/oCUz5sMafNNG4SPoZ8M00ALJjA+4GP6qePKEPzBlq9
JqQX3zlBDrmGy1GjydtUFKazV6Yy36tuV9HDKeErRfGHpVOpXJ5I4EENrK4Qjyye
6tqZev+ymxw+BQ1Py8tGzdslWbgZV214mtueeYwMRleNOk6QMJfhiunGFafJkgaK
1aX7xiXQHZGNEtvJEQcAh39dpp4UE6wxU9T4a+aFw284FAyBS+JLWH5UlwuNmXoy
IGQBa6z6gtac+d2H5289Zfbg4cPZHZ3/mnBaQUGRqWXjV02XULPX6L1/hP81BBTd
edFF0uC+zh3E+Ryz63Y6mwHgq12F+HrOrR0CVH05YYwxWuk6i1TVzMAkAPm2u5cl
UkI7E7OLMGqkF+IoDFBUlYo6k8Iu+0bHPrVnd8T/dSQSLoVdj8csZ7t1YsS3Nuwc
4XK4fCIOLTvP64p+GDBQeALMtJxyyRbMZaqGy+bsU2lR5Y7Ml5v3r0uD52/bf8QK
fWNIFsAtdWFmfqtYOyJmhMF7fD+fVF3iVMS9eOVkCg9BBwPEgnHI1kERVjzwiCdj
sBy9UVnz1fUjju8Zac9qbIouSTvMHXq8eowx+qABjfFS6iyY31h5RVhEl109EFv2
lkGkbmJqmBn6xEwkPQ76Ge6at64Rfr/3kuiTBg2e707WSIM7o0uNnKUIBq9nrmNB
uUgLYc4+bHONWebcqaQ9Ktl1WTkXW5xk72i3HHv1NTFAMqaZaCLD83HpHUNU8zhE
mYKYYqo5x7WrZOvsGBt+5sve90RmDqMDrADrS12QSiztxfxDG/+Y/6DLEPfNkLkQ
VBVXnqbHaEL0UX47BueTtHzDr3O/wsukM5Kxa7nXHzKwWrHo5xk2ulILWjtyxDow
F1RegOru++NpwWEe28hciwiZhLeIUgX1DXK8LW1f+pwI3DgliA3+rc7CMD/Epnqp
iv3ZQcZHXj1U9KiZ/T6V/fHT7b9sZrcKKd10Z0j8q++FYgF1x2EKU77gy7PIQWsF
tTKE1CiH8fU9xnYGIBeunNkBPXUB86NQZq/mEmyWUlE4zdq8wizrmaJpTOtNlj4v
zD7d0pojrvsTHQXC5rCREdFwswgRTJOuftOMQyfA/kOs1QIaahPA+i1szP1ds8NF
n5Gjqwg6OwuhPeS7aAW7fD6T3yUQzMMuVpVpdDmjcLYsaw5b3icLnq3WANd0mggg
XHhuNDIMyD1LYRiYFQBUwBL5S/8wAvSMrmA1+Tlka8EFMt/b6B09KsuDKM0vvM9g
/9xmatUhteW6xl5UxARYsv61vIP+FhockMybxeHzfZCNdFMCe523rEE+tqJaSemK
k3RcoPhiNdqDg43kN+DEEC5PYWpdSSFQACFrKaGPK6loRnUAPbM/WWDMHCiqF6c/
k5kESIhpKY/K2GOnc8zFa1ifSIiv39iAEpLmLtYlC8qzGDA5OPWkD8fZ6G8RLqrp
2xX0ty8UtjBdnanN+LjewH1BQh20qpsSrlhXuP7D2IrYdz+MBUisMgZC4bWILU1a
/4wyckruYnBUOz2d+a8botFGvCoMq0kmwf1BNvBobIWQmHAXIINbMmPkvjAmA32/
/rR5FKoHx8m6neYIjhgR99RfjU/jZ/CuHOtidueBJdeoD1oY2e6uOfv1g9IAV04v
PlKcpsx7fxVkji6JtaJ7BjVOeKfYxcVDQ4JpxpeQoH4Fud8wocvG/LErWdQraRBi
UgEq5dXSipXM1vHOSTK3ISQ8sh7eLsSFHAOCkajvOx5s/jQ2iU/Q0GwZj6UFVnm2
JCaXvuoVeKdSgRGtuObnmSZlSoUWE5yBJqrqm9nVEAOL3iY3Uru0iJ+ZIvUxVir9
zNR3cDTNBqEn7jMI1IDeXJKrwcgQquDcmwOiWBLqSGPqg+BzM5s9pILg95mQMQ4o
DC9NCLhcBTNOq9s4kbm19+PQ4K8LzN6mY4e8nI1YFxBCIWbCLgkVBu82dWNA8lCW
FBW8lEGl9X1WfQv18ErWCS9uIWy9uDKrKfuvd+TomsiM/rbO8ogk5osfvETSMT3K
NeikDJVQAp6nAikqgc3+FCIRq5/tRiItal/xK1lxT9kqYRa/Eg6vBjvoQZYF8j24
dZRZFEj5Nkf2Nx/RwYgn2IuLHg6amNkjzyCxusWtPPnwHlBZTl8s7ND7KThf0VIm
01C8FIRlh4e3HMjLTYQYtvTN0Eyr38rUbP1qY/MjzGaTIvHErXHqMdxhUKg9k41f
I+tIcTaZsOj78AmKjZwuQSdvt6uADgBnx847Lj2LP4DBQIujPmI8rhsd8FNg/e3m
IwT9qKMN8rpwaXfDXlXpPrKnZHgeflfgBluPYiEWPgVPX1NMBBrVyld9+6h1eQm0
+QeuOk4CTMRzpF49udFrZt9GV8XhRMxr7DTFXTbbtA53WYISr4ymML1dIf/AxoYe
3v4Ph6IZEB99uxt9qxAtlr6c3WQbYGSvoIc2+Th3VEas8LGCH6mz2Pp/KsHrL0CP
SmHbkKy3od3xnt+uEmFDQP+PE4GvrY+0wgHJOWyNwvaoQljKycJ+II4e8jb+4+bE
H0XveDvy/xbKJ01RDoBeuzb2v+1LmKSnECci9MMAjWeqfovPEUff+g+nhAwLAPZ3
MYyWUgbtT+fmire8IDsHs4sZw7GBqSSok6IS9JtdQPYkHbma6d0CGeSviPvHiE8J
7g/lxlwHGWYozpR5pJaT380P4bLhbnG3y3EEuVY77baG+1ZDyOC2uqSxdkyBNyrv
aqGV5Hv1j+/dOI6NzbR8Y1o75TRtKoIR0ZHKZUtc+w39oBUWAMZCLbqY8aj2Iq+1
BWDK4tggg+LApMuf1rjlhPP8gQArqlljoPdAyOuAD3icnpSuiTuuNQyaIgZE1L6x
imyHmTGvY9NR+u0Or4uP2s9j6kZVn5nm/p5N9Kh74smivJAJIQWTYIJsI50jkfxz
DPoqb8cSlQPhapU+5IqOZb/v0PytSggdnxvj9tRTibu25ZX14ZCU7Cp0BXrbG0kV
9INOwnyZzHpaaEzNeJq9rCcQM5rrJwqAf51/UKsONZBctnRKjFJdV1lwGmXMdnOI
37anAgn6yikrHTjkyLFj0x7FXUijyWM4SWn7D9JPhYmlF3VZVLHMBLRlPv6iNq5u
2nyVLQoH5J01102x8lVxGJ6MCo7/gKStJ+evcuA+rRz7TQYE7oRoOdMrbB2sT3Gs
ei8YmXRcUZJwzxlhKdWW+RckERS2yUyqZ0HKhcofFr11HLliDf6Lvx7BukSAi+/t
O/nPyris8ogXKDq2uWG2H5nRAJY9GG/YpXfv0QvlI/wYrZM+pcmMkGYNd1VHhFRh
q+7SGG81/ydEupyPvDoKX+zZfa0TqpOFg8J41MibGK9q2ezLqFTqq4ovtf6aSmMc
Pv0vrZbTap2McgInOXr2sEo1xHgXduwj3E8cD+nogzmoq97HJK98VQEISgWGd9xl
qb4jAuv5qvcPxncSNMUBBixqjPoXkj0SyazmtI96qYoiVke1ADupf1+qsNHusu/L
twr90SghLwDVMvfL50QwAPm1qSiNgHVUtM/eNr3UpEMmJ0TrHfzRu7AnIE+DVU6X
pwXOF0wE5CTvOpMdfDKXS23/Cryn0a7iP7SpgC6fAaOfVZCCt5jBog3uY3N+Dkq2
kpbmq37DeYT0jTy9HJUFJ0TlcCobBl0AipBUD8WNFl1kB7Yd83Aa2e2fyfLxqd4v
gPX39aQs6iu/leUqo9E3TuEOPRt2enVCoUqT5oIJPUW9ipLB/mjKZp4hlaCZNQgN
IH8Rd+kPpO+7+345E8dm5SDSZuJ/hKeoIFLkmQiWDV/rQvhvFWGUREXnjvbfYkEX
rQk4vGv0AZyUKa67kXZ9NDjndI6IRr26NB6wxBYvu5q9f5sdjnSC3Jqm2JJe/ERx
d6W6MVZvy/LgeyO2jVG6yrpLIqXEiXhCyJKHDHwtaHfA0r+GdBEkOwuHWVri3xE3
2g2UHbMXImGSEQvc65kOEs/323Ov8+LXMnprUbE95o0BOAaFKB4y4odvSVeZHKs3
V7x6HASqh3jLTVknbUjK2Fm5xBIUXd0otcsjK/1SogG6oZSgKt5s/8QCd1LF0NjQ
UUJL2vncKPI39wszhO3n8r1qukMNn0EQVguw7aY59orzcBgekJpGytB49LUM29rA
I2J4APlDrw74DYrEDmQKZEtcuQGkBsahIxB5KGy7DrRH6wxXJOSWXdF+yn+80yQH
xHb+TiIP/0asi+pEVcRTzR5E4Rn7WTKh/F8GOk5jEIZmr2HL1xvCE48QkzmoEidM
8dci8rd8HAznZ71ElVlGSB9jsi3VUqtOJQhjUhVOQCkCV9/3YRbpg9UAjMQdWwhM
czzMghAYjpU/v38d//u0ZtIykoRpH0uw7mtBBteVvfkDrwDfAtUAIrn5j30yYByh
K2Ohixnd1oWlrbwzfK7vc/C2MdiwVkT3/G6c2bChLhCJa/qH1GjxaMyk74hkwx5E
8D5O1w01R0VFW4wNqLIScVnq5MhiHS9T/eaCCAJBNt4LCDXAD2wLwWI/G+nWR6i4
6B72b3jAArEodMhAATI5B03jnr8xVsxocZThNsUe7IJ6D6Awjva/y5mHPjMJ4b6g
LrqNLlsZoM29kowIFlkP+OxVZttvUrbxZv452tsOqO8XQWTwYcyODbep4o0Unzex
g+E8GRGwcIHQhO6Ln9sQWDr8F+b0FhE/Wn7lEb6MUL8QR+BOgui49mZqEYSUAvO+
VL4UF1iVkRoaq0kH7pxtmY19rxA2LIoJ4HcQapOLN7HA0aBgKpQrM/KJpvWi9PVT
BZiXIgoapmU0L6Y97ZObQ8xbVbKBKXSPXiY8AkRf8vWhvj16gNtf+0oSwIaiq531
6c8NvPLTaHsQ4tkhkiQwM2hspbISknql6e70H4FUD28s1urb9OysmkH8uvDlfnZ5
15xOnrr7wdjmU3jTvnirLVmkxSzIl0QLbEROI22i3GnE3KO1poq5IyAPuZTbx+QR
BaeiedPjj/CMZ+JblIAnTAnN9JakLkgfgSVeGHMQF6BZIBA/5ef5ac/yg3IzQ9l0
MylQoMC7YAH7FBpejqjvSRxTxq/o4k9yvjyygdcB2GAWsZG4AE+6g8JuwHaWTLko
QwTuQzfIW7I3ZHZi3l28iJzVTf0tTTxPE5Duj7qvCctkW8+b831iUYP/X67fKFh5
Xv/0VQvWF+0vLn6S4iJfmMx0MbB1Uw9OZ+1EAnguICAdfkB2i2EHTDlDuvgTHknD
gg0ky72N6SFZn7TEsIa/TLzSFSmvUKppEr1xMUwZHOkjuIcK0x1LGQD+F7zJKiNE
QBzAcIXD7ac5B5oNRfbS7MqnW31E3H1JH7+k3f6N8sjx6q6rXePFH8DxH/f+bFzC
325WlYdH4BjifINz+5Ucgip4HYyRTMtK4dwW72w+TXqZUeWXPLNAc4frA7WYzwx+
Q4TPRmLWa+IjUN4vywW6OQHjiSDvDjC9w5F0anR0zDSldVbAob0xYxBsVP1YE5W6
f0Q4eKnXs/rEhqoyTBGsp0EXFVyWq5+xETb95p1T0ZtHprcirxs6GlYDlj3ST6Sb
i3S8E004gzg6RSY10PDotehns2p7LZCMPkv+XOMWX0CYqmupNEeEJ5RgQaNCcP7s
BLv3dJwu7eTlGZL2vCYOFPbeULUtvDzt5/Vxrk/REP6gchZlx1WdXvtAPEEaKRrn
AYaLnO6IKQFwjmn327sqOrizpQjmT5CmOQiDJ+Y8NpKy3II8t5Jtq3MHe6VloB4r
6fHTzmybvVfTLkqWwZud29kNqATg+6ka+YIM8j8Y7QVAUAdf1iofMqskmvSgEJr5
7+zp/lGhFWezxhDYk3fYpOgsid9aBFYYnMvySViIWhHw2xLfqhZ2yQQFCsEM9Q9I
zV6A71L0qOFNYKlzmtzlPZoqFNNWIo9oSttzInbwIacKi82P5jl1XaqoMOzD4Gu7
bfRiG5CFSpVhBiuZmJKj1ydXEFyIaOeEHKP1E4KKMCheXd5v6LwHpkugjO3nzZ/n
ybPojQ3iT36Wf7LLNYZ4+YgZBhwzEHbYFSDBAAgl/f7KRmCEPkXPSnpCS16ALchE
238q7pez5RwHfrLzXTw0FSip0JlHnpn6sa5ymoF5XYdo5SPq7Hv3k0wIG6gSSIU/
BVzoKUspWyXIQ13sufmAcPTGztbChenTp1scHqEaddZDhBXk0hjUml4yFxit2wru
7yWeTZrd7UpeAl/6oICHY3pDPM808UwpIHpjiwiOkJJMvAEA57RBFxndbYkY5DS/
SOE5LulL5Xx1vByLQJDsMmXZa9S0OXf1PbnOxtQMsrufz4BPmtWB7SIPvLAEdz1M
Dc71dDl/iUDxdxmuLaUMFZR8Lu13apErbTTzZ/uw2JGQ2dclEGiuOgXS5aD0VpJZ
voPSI2B49MQb/8v/JBxtAW+98QvQb/2huyPfHTRomWT8rvbCEIWYBfY1UQEmlOcN
jBi2aLqS6Dll1yHirhZ4Nei8ycou2Cja7VFdJ+06OJTfOU9adiop4xczxtpCU/Q6
k4KniDR2X+BEG96JZC42aoflOAyd6BHi5rCVUgnr/QmK+yi+ezgN2v0ngP98XmcO
YFDvzm0wS/a/MNDw1aSd+XoYFzKv3ek+i+ZfWI/30CmLl/s08NL5VrVZTVy7kWTq
dqh2+ZPVEJn8vIZA91xaLl98taUg2ec+KPfI8V48P/FvAur2gtQ7v/tRXloY0WrE
fJS4PA1CRAnBpE8eQOye8ZT0dhtYH4DuUSDcpvf5Bu8VBKB6NvmHMC8fgNh1ahML
P/mwgkYY7IKdZJ02OSVBxYiPa4UnDjm2JsK0Qrer+q1Tll7BP8x5UWR4pfHBOpPE
1/K1yU0HyB2n470vkk5BPlqpYRBDo7FPb+GKFOR8OVyt5lxLzfZ5RUWEDqUWcYyE
mEJ1iErLUhXd35eV/CwxIleNDtU9m69jqojyay0fYf4aK4BprRCikJFOx1mD1WiY
Fk9mU4lMz462KWMXSST8iqazk9JLmahnKNDl8AP2Z5hiOB/1h75ZwY0YR444kSRT
F35wOvwOYSzzDvyLcvGUKePoXQ0fg8yJ94XSDfYzMKEaLQwyLB183Wq5CRpbA3wR
Jb5Y8rs/lkWUYF3V5W3VHRlsqMAteT76PIcf3FWFTK0M3LyPQVgX9RSJJWvtmnaH
5PldzI5khecQqkdQWsUDlvgKGruYpNkUXaJufmF1dj7xQlXtRQor2SreQ1qX2/9I
gRK0npdEWZS5or9jgEPqJrXwFok0P3bYv+qSFZNaNvruaKFnyybo7pp2fEDdShzt
YQhgRoxddwIlt25BhGmjL3pN1SmPGrurJ3soOti0xcZ6SI/Spcq1fENy/ea1qpAV
2LUhhJ4qoZdppko6l9D36FS0EBVpKmC8Dme88O8VZPLr73vwl7P/zTgDoX1fiE9T
ZewszmXbBEqFOnGLSOnQUBt+iIUs+Tg1fbx9nwjEyrXZ/rV2SuFZtqC+BE/IS/8C
vQOWA5o6n1oH/pXd4jWalfIv66Avhk5PXY3WYJ+azGUUv1saFico4CVluvs2dqgw
jfAHnydcU2rTG4FY8BWEQrcxnBl9nepDYBai0UHpS81R6UnSBXashz1aqDdFuY4/
bComQkaS8GFWJPuu09LqzfAWGy0OWnlfnN1Nk3h9cIeWIBOiIYkdcTMWyl7SFyJS
cL9ubhpvG4u+m0aRvv2FUGB/jYbkyhIvkT7TlaC+aYnjyoxxsWGYbbmWljmVrqyE
7q7fbaxEhJZspzdUMglg4M0Vg0QuSOKv3JNs3wfukh/UMo0wzGY80lIgFaKouo7T
OIxojgqT7j6nRpfUwatt/EWnmZ/RGHXRku14xeYQOrUU8h1AUZcHPhqVlsTX1p91
Onz5w9vOwYuPXUwBoiEobWSvmWlupRWJlqW+G9Swhf/3Es9Au8j1rFA8lc78rWTU
hvsssg3uUXIDdKEQPBXQjTUl/LbPaO83qer30jbX1nQClAf/hOyqCJ0jgUFRmlDE
dnhjqzzSmTs/CylVChQXn+8aNsJ6wFiJCKSPSRaVGG9GJHgM6F3NaGMxTBdVj+Nw
lY8nQBMXNF+1pZgjYE9tDf0ZIMSrWRLBjeuIAvMGBYfr+hwCfiyd15/t2NGX5/Mu
z6iSZ+YRTeJnqFTlLdBFo8UBkXPefKWe4aPjGsV0iASAv4FQRYzyl5gHAvL1guqG
Rj5iUeCb0ZQ1TmQrIhpgQSOJMJufwRm2NaeJ7TL8YcvyATbbLq57spAaLzKpE7In
RS1ptfhu+JMi0fFduXMlPlGzuGTpd5YLA2g4O0VNdFs/u6MjMOrlXNW2oDQiQp19
3N3r3PVRgOZvZ54xqnNxUgdFwBvpkrU/SedqfcZDjX86Ja6vodW+hbDL4APP9y/p
zOJ511SNrj52HK7M0t8C03hO03FPsBIhPpKitc2GqiaCf4Sk74LRe/y+uc4WsGiG
xQGxTORvpZr2eDKb0pLzc+7CWZqQgVn72Q3rIR3FmsBmFx0V3CAY8vu24PoiBghV
x+YW6fumdlPZ9Blsr0kptyG7a4kQJfXwacAGqK10hRFtJfcDnKzvXnQpki5IhQh+
PoMlDz9cFD74KyjOiQ6PnJG5xjPbBLlWmwHT8WPqwXEhjvLam6Mmf0QulqevX+Q2
9j6kMQ5ZVvMAHQrK3ptFdObZOahIyrhEsFRLLCUxzio4LcvMsrK6MfU3vubiX6ty
Axhczgm2v+tAZEsYlBQj7215xO9vQdva4GJT6bz+X/TkMx9GX+Xu4LV3qKPTikDi
QmdoiclIOgq55QEfs6Q81iE7CDZXFYFgKkjTdR7H1wNy8hmGTMJik1Esj+kWEb5F
EPOoV//HE/3XkR146DvfqKO7Qn1wcI1qCJtFCD/tiGMpMnwrsxaIrMj5RvupleIJ
OQqepoLl0MIP6gUonGc3duzAtY1GRTZfUP9WfjulAozKY9025DfgNrVmWOk3taDj
A5GAP7lPKzjoZpbkgOvf1KLlov/QwK/EgT3M0w0ZtrQZMBPQcyaLEPv8H7CWDYJ9
a9cnxOjbj7xx1yKbePpEVVDY7RncO0TMG+uIupw2ebPSb5efqJjb91p8uFjbcphA
2PosRK7elxHAdACefQkKW6ziNd9uIgvDNRjfRDKQOpDhQ7bJ37ORy8wr/sJsL1Bs
pv67gpmrBqKsrahpykCWhHzAOvzIfgw8x45ZoOSFSEUuEp4XnKvyjkd+TV6iRupC
S4ETqRT6DqVrMZfd7fFO8JS7DH8CnpBHH+dxIOJ/Rh+a9tDcMN5U6a5cHHE2jNBl
mNnF1XsHOe/X33Hjx+zIZk5pSbWWOOinnHKyQ0GQazhCASKfiaePyk5HxCqJr8Bl
ieOeygeIV11oOyNmt1ViFcU+yxK5oxuyw3jE41JBNn6RM2Hjf0wGN1MN4TP7/WiH
+gD072u5CvAACnAFZPX5Zv7yXJL1d+Esk16jf/shsb/hTZlCgGbCRjcRVE9A51y9
e86I7iZHADO41QYO+18d3RRSd9Q9AbNdNcp3uAWn3ucXdl7YrXGcm2akQPhC3eFY
6ifbnOoVCSAVGNXbES7FxeABBO64xBJnIf2ihn7zGeVyDy67QUI9WOO7M2c/dxCm
ylXhq1wrP3ww0vFv97Bbisk+wQPLn3UvAaBQTlT0QBQts/0KqakF0N6GxprFQUTD
bF6upxnux53mcG8WaYg8RfPY8qmhrvjKmS7A+AuuhsTrCyr5s0Cle5azFXg/KOdX
XClp7tyTPlrrib1q6KbiLEL614MDUj2A4JvZtf5nEe7aVvc6TFLl22Ft0PsnuOlg
GKyg5HH7xS5i+X/tO/+xxZOFf4uwG/Q4RDhuQ53AVKNrBaZsjHCzrPzG+Q3wprNl
WGgfD5sq7Y+ZIw5jiuui9hg/tA0CiMsUK5bWey9dzeI4JeaUitKfRXQGgGu5vtr5
2NdT7nI+nwVHUftSY7iEGdGzC2ljtcu8CHaKMAXTv2fFOs9eEsPml4ZP9MN5AOBG
dMF2pu0+YC4VrBFEOXR1ciGdJGlmzM9GU2J+t8UWtMH3BWhOYRr9cA1LE9mpll2g
Vmrmbrnri1CI7RX8f1fA05VCUhiAj2VuHkay/HO6dEjlJcJIQAUF8PggQGGPEeA/
UcNMjK/cVhCJu5gCAGge/yxm8CNnROpZLlVzcNYZlfSEXzzF5h7rJYgV3sjTm92q
uN/q7+eUPQQEFV+3Fstf8XJfWrZXyXlDtWftvU/66QGYpyKkgscLz9zmGcFmUsIu
EU/OBNoCkAUI7sDucRzOozg0XDWZ3fbJHuNW0Qv/+mNUPos77HOxuEY0QMeI1Kgz
/QbcZGjaYU6c1vmsR3gqhnx7lnKlwGSPVrAeDfObzX1yjqaaCE3QEhgBYEqblEqd
9eAk5c2zTSS7EvTQSDasFqqsonJJGM3cqW+hRtH+CLk4uwE1H/qEgzrk6bSiCHRg
bDeocy8t+HY996aZjBHDj58fo/TDA5qx7L10S3JQyx4mH9+Sqbm08X06wQAopJsL
u+LXBfGbt/jUjI6WfMJKC+Mq2MrfkwmWKbkp3PeB30ixKx5KSQgylcOWMyta15y0
aYNE330jAWdKvKJinnvHj9d1Hg9kEKq8sq8huJnMkNRhkqNntejwIE068QJGEK7t
SUrQCuyUrB8PiKy/RXIB/w7rAqThMu3VtEslsy/XESyqSfyyYqqmWWayooUdbwcV
Wo1UyAiBDy3Z2lj2tMYCVAvmFnh7VunHTHpIIYre+VsP0wUYQrutZTul+u1lZ2Bu
YQsWKoGCAa4AKF1dkoHeap0L8Ew49sc1jD51ZLKFlXdYaS5REkLdAMCeX1Duk/DI
pWQJFfwxllxoDTab7mCENED9C1jiVoDVz6z4cqsDxYqnThWCNzsdH9qrllTjE0Kr
amDq22sK27lipcGISd8rqnEFf6CI01extQ022++FBwQjDcvojhLeN9njEbkY/DgW
PUy0WWqTvyZE1ilfulYKYUQHSUpMpKtB1QA2VfMnroQhbGB1QZHjY2/sRdWnso+5
oRCmavo01YIwIK11UrktGe88Bu5VoqAU+ug+/8l4a/k5VHV1e9m6++wk3aF7c09v
M2O/PYsY/oHrax7kEN2A9Qu5HtUxnJiWx6Na2fw1ZMsdrt8juoP54jBEhlmQaWDj
1VcSkqA88p+sQd0bdf51zW10KKtsQTo1+vCjOVfOis2TY7dAZ2RoLEXRV53JqVnA
id7c1J9fS+TSJrJ4QSGWQjT1E/xrqpPrdAV7MW6SER/QIr0s/wz8jF23UaGLimoa
cZNOuSNtHaTAF3BbGUFwGmCNB1McWKvRRdXBkquM03xSrS3DdkHYwQhl5H6yFqwD
huN7EtzLwG8xQC5r049tnfGJFslbevE5ldVqJOEfxT1mU6SXQ6gxgrHh5iwgQd6n
VM9xX5pt+6KVmK5zbnG4sDv7U4ZuE+eNL4ZLCXuHJLUO0Lqpbk0qS0IXPNcOQ7LQ
WNsVwSVDE+/xYa2Z3yKZY75YM4exsLaEYHObes1cqn7qVJkaN4/g37wfJXuiHojF
Wim1V3HALI7AXsl0emY/4V1hRsKrog/OHx94izev7yHXp7M62aAwI3xcqm8yE5a1
hZfObeBq08FgQmbtlX4A8wq/Y1dxrDo7wbuPOtS62dmYPcvt0s0O7L4a0lPeWY+6
gFkpfFTOn/4OrUBWhhbdIlkp5L1XjaVQxh3xxQZ6zy2FANAmGLNOZ7FEcE6M3uPH
Pd3eZMQcEhGlFK9n/9YuPY94qt5oaOh1YdWOThW+LQcAXNdEdX8Q87p1nFfe35ql
HogzpJc5lZTkpiEJ1TV+uUAzywAEEthn7eVRqU1ow1Q/aZ6E14q+NrcBc/zRXjeG
1Bi8PN89VtceNVkYDHcgklmsnuXQwsv9fICVqKi6RI9RJL6Q7Vdhj5mNl4Ll/u/D
xGDPVqezsMU8IUq48fmVy7/eWgJ7ccHuxIaSHq31FhhJ2w8kL+gJabY2xIdmCw/d
P7NaS2HojUZqiM9S10qofnL6nOHTtKsgtCbawo01PUU3azE9HyAQTLCJAbybfhuo
exIG0IUfV1ElqZYAVNqcabjkPqLvYiBg9/WBWWNhgdZ6+JNVN6XwYwKtYKmcXbzh
r2oqkUBHDKbW99mSV46zni/vb02c5GwjOODbwRRzDHbiqHZixsBk7GHiUpdvyqPm
TZ2H4XhQdH390cso2BMWFKd5YWtiseeWpyM3/k2HwkBQT/na7OGH7pW9Rquc1hKd
xyKC1hqysNglh5Fls4aoMIe+vIZKp9SlI2SE5b6rQ9QAzl3iyG0wxsLEUMC1lS6g
zwijUTVSA3wsF9Js2iZKJ8K2KcUSxYV9lAAdIm/5URo+MeL0xwXhQr7XFxGlJSmY
2Tt3UaWi/MHm1bwiefH8K7hnEQ7NfYYg8GDbpx6NmIR+OGfWLvbnjyPZJPUF4GQG
ZaH66n2uiyDmQz6mqiuIE2q+RvLwk6ADG7g4gfzxoW28TdlZkJ5oBDRWtHOmKYsA
LilIO0WoYbt5VY3fcZVbWkbSPQCCPI6UPMOZYy5udGl7W4BMwy+6Rn3bLnlNs0W3
SBlmxAXmI84pQwvO3qMbV6D7hsnOCch9l6smYONzvI0GgoxHKCTytlE3Ux4zV/pX
NqFPC3neZggVe96TULFlwDc+sTKH20qpJWKALrBFQN9P942oeFAxs3s2UcSn2xb8
8BF9L8xnTqZIRB9veVkh0wwkEyTXvKjSb+PZ/5WmYxmEnXb+rkiD5EW4u/Wyn8rj
5488ZpgiPP9qyXAoHCVPBSWixy9xLG26Mz0pCJc89nsC8zUKj85eCmzRfmJRxbhu
zqyBYem7jTy2gqasMVoI4UTuC+kQG1bM8LJluL6inSqiDAwVrWfLJMiYrwapgMjR
GHu6AtNm36TWKCgzomrp7gCIMwksBjs7qRRWWC4Nm2tVjmjuXyKbwYPEt1IMxGSH
edCQugjNGgBr406B1kiMNbCiEp1Cx+Doy/g6JIo2XXvsepoMJX2DRoZhj9EirVln
fYHWPYv6yArrJCnWWmcgJ+KmB6Wc4sUshJwdrVZ+o/PmW7TrLOGxgYA3vyDgDYS7
PZTWouU0EMgRjnv+gVuOFfXWM/Mz4kypAjFT6sOhkyGu8M0kfbUF7EzNi8c0lhg9
Ga6gbDSj4cnHhIyZREIDAG5OpHjmK8CuX7lm9HJTfqmqIND2292/1hkbexSGNGgm
A0gr4ThuhfIFE8tjAmB//dIKm7w4akM+HLQ28ZV99ROr3ObSPXck8/hZ2C/kjah8
iKiQDYAyxXPbGM2DrtRIdY3kqjrhokVPjYmJC65M4SAEcvmdKuKmM3j3alUXKZYj
ypK5ayHf/r2DNkLaSiAYGJIebzyvSXGIOD5K3MxHi0rlgFv++cTUvljBc87GRF8P
cr1TIIA7LpVL4aPAqF8F5Qz6onz8u4nBV9vB2BdvAOSuOWqpJSumK3YuBB7I0Kdt
JQQKM4VH71aHl8azqNIOH5qzOT9T7Jq4CdE8LIYD4wLi3uZx6cviy3ZBkm/VX2kN
n1tkSsK8+kIrOtaksZU59b5efFa9paOvhvpD4waQCTnU74jXa0jONfDD3fpcktgY
dBBK2fPAXPMUMf/9PLT5iTe67qKI7R4rHGLhH88zvq1pimt/WlaFgJXzCLNRqSot
rKm3nJzoDdcfMYNwpcVijI0/ajPKw/yaEvuiuAC9ormt5Xw20kM+afZKYLGawsEv
Yh9NudLrkGUQZ1QI/vkWoHjHe1bQDLhr1PHVBl79/Aj7uLQ6u11JlQAr2/cPD0Ma
2m6WqWg+mza64u03ix9zhLLTvN7pQmaUUuFjGV3y6qy6oFjcgzIfKbzV3HO3hKe5
dRTG9qBUA1Fwwt5G4VlVLO56CchWVeLc8KzezjKQLVKScyzDICiV4i6xBR/ZwKcg
X5Sle/BXLrP0otP5VPsuB5Uozh4PsHlI84fgokWuiQC7/Us/Bp2wt3ME3ZPhtc87
yLwRgCKQX/x8n3CwOhWwu1pA4uXbX9Ns5+mKX3B42YFrM/16QGPE1xYPpL/ZEQgp
/lE3K9DjjaKuBI1Cro0OXa8yckpEE1rm3aw2f5ElJjZlYMZoKFyzNABn7F2ZyHPP
45n7jKOKx2S4xAp+pn0EDEyLLS3g0PWckIyMquWwBYv7QzIU5il9E8cUYpdXwjlv
Q5Q11j7xhFjnuDxo/4qITMo3WYQUS+lTWV2WZ5Kt8PSRBH8a3TS9E4IUzFCVSE0a
UbdxV0A9NEsPF0yLDTKIFjC6SIYzOUYyBT3wbTkdb9bsL8p3FuaXAzytAJ93HIOI
ajFkx/H/6w8n4e47jx+rldEwEKfep9uAdcmUPO466AbzUOviziLTVqIGitHJiSwC
gNFUO27LxHj2+rkSUeFwyHhRvvQmAYCEsHXvladFtAOksUsPyCPUyVHEiMQIykdX
rQmpd/Bi4smGVAr4s74EvQWknPalTS9frkGHHrzxL8OhPkv0bKzOuZcsvdB54iD7
Z11pK8Q1dnCgMpaa9N34ktWTUCVDmN/S+sYUnb21WB8nkSDCuasikSn6rhptecmQ
cn7UXp0z28eTvhYsgA4JrZFoxgo9DTihoO4Pxd2cHT7+XppJgDfXqGH4McWaGDV4
F+SPhMhfAkjLgmZhyguNuJmxNHoLYrGcTvlILEA3dpMKlk07ZQAQo+373zaN6jkZ
Tzr6obJ1HXTzmHbLOcNCDEQQW4k5U8m+skuvDrLxVfz1q9tl//V8BfrHTKzS89qU
HWqj/CPXAz1acOBb/81bJj02jOovJX2ZONxHLaKkndqexXsxK0nTZ0+R6P4xUNqI
LpPwlC0DAwagahHYhU6cAIQSpx1eO0M1hIV/wKz2VPpWGDAesvdROG8qU/ux4Lgu
gtLkaHQx0vQCdwnWAqc1W8J1Y3nxVQh+qhkckxm2CP5cX68bPNPJAFBBag0KQR+d
nvdWo5UK5vR9XyuD7sNv4npTojLRQLEZ4C6NSr/AW0KQqGqXKALLUpVvGRfY/31P
EBWI+zMRaWAxo9+4z9xiDtofdVxIKfz8VhtkM1s4b+pbJ4wa+092o4Y/jrdHQf+x
GWlJ3LZIj8AYTPZU7woxsZz7RL6y+X6k0T0dbMHhj6dzHXWtXqKQx+lq72c9S727
bvdhN3t9aFs0sCYkC1bm4P9ruWebpMflRMhnc/jndCeXIh/VP020sl3GMkibCy0s
91RU9TAAHtMR86jEA/Jt8EwaAqa24DXph2eWikcWw6G44vPFtVDXnlCjrCxJwZ63
QkJbTZ2VOdJiyVKe0Ee0tQkT5WZTnHP8r4JRU64QXYAQg8YSmbnCXmAEskU4caSN
J6HoVQN6UTv2o5ZUs1AJvKm/dx+n66jhWMN4DFdRSLBulzK8a9oxHeDpMxNCVgrb
kAJD79V4jYCiQ4DpWiK8fKrZ6Rc2bJuzO6Y3TfTvdb+4zKpmkMQeZMEv/Ct/2oO+
nfltd3siz73320qfmbssXIwtjj85DYismj12Y7r0bemkkOQKos89EHe1i1B4E5nX
C1kHT1TXqa1KR5x4eqkPDz9pWD9b8eBS2PHJnJk8xbF3J1wRWyjJjKGoGk5vZExk
DmBHAMHDHoX/0Po1vtoCE60qvmipSCtTWtYPaafbBBjPeECG843WYGrE9IKWZLDO
QL6V7tvFplLTxEJWZ8ihgMZ3sczrodySxsckmxmbn4Mgq1OpZqRcQfL/DImF9P47
2nNMLQr3+W/rx5Irh5/rEbJCfzhLLf08cRlY2zUdCwt/KoPuMF6fzyU94+BwzSuV
GnPApcDucljnFvM2N5e1bcxWmpRFby21HSXCR+24oryRya1Q2E389+8X/wEZb63U
UvbMLlx0xPZUZzd42Chy9QHkstkZ9SJoEpQxPg1alD/YHcVEEFuMfCXo9WBnIg9n
aZjiqgEdN6w2eenPS4RpEPK5fsx/Y7V2jlJLQcwJ+BKD86+Fm0BmYJN0DuJrX26p
7XXKxdWo313SS6TvrJhP3mT8gWCsrANp85KQBtbDB+xT6y6UZZ+GEfNKoy92GiY2
wnKu4I6g/o1Uk8dFf2/d8z5AKS90GK9RbEYDXEFHxvKhW8MWq8sS9OwFEtaiqKuS
uTfMLvS6qwffKnXjUH5gUkyBHSaVi6c0P4L0n3EB1jDSppGfUPHkeIq5L/fY2eEi
9FLnxSsn+hIU5IPV+qdsgscPTfqOtSyuXd5ueSJjiNkwX45KiOMTGB6tAsTGLhOg
v5qAU1OLZjtqa/VQOFE+rGqh4oyz83B2sBoujMSu5lpqqR1VyctHmvi5OFMz/9pB
8OuWRGkt8yx/hUSiKEFo70DsQ8oZfe/hN1yuzoX6wV9uFP9mVF3AT5t3eGMMcdTb
2TfbC6YVxxpjV5qYa9sXTIqnkdldH5A9d/HV8ZKSpAOt+dGET4BN7dupkhfsYbMG
rdE4QDUFNH8u6DlvOlGNoMtXe+bZOmBKEygacd/2STBSW8Gut84epkzlRncaUHJc
VJ4zKtccMWDQrMfuTTL7UWPWg2+e/yGWPb7KyhgqVos9dwRFqYsAG6rp3uqCGfld
Ifpw4XYGYCOSrm/iEF8trkSoD0CFwgnRDPWmhq4epxyjG/LZtcHRWJw1U7CMaDEt
Xlti5ucL0/QRVmlxpOjQh4om+6iUg3hXupk4iUmT+vdCFilkEBYQwU1tB5Mq0twY
tkhSNsOPBV8Mvbxofv+AiyzOGlzFP/arGPHZrj9QOORZQCAUDBMEm+OQWdRYwyrD
RoOZdA6HylVcZ0m7C6hIi4dKMPrRHNLdQT2P6u53OSelnhuybIC0OZYXB6EYUpq9
QkoPzyFrEZi7UQfC8O2IZXc0LjnSq+/VLw5K5Du4eW0M7UkwdrVbJ38ChAtlZdL1
bg+bN9j87p1QEyqGUTSCCGKoY+0wlyWKV/0H36X2rYP5g3bSlvDhMsBQjT+xM4u5
WzoCljJyTLLdfWXH8YvxC7D1nPVADUBUIaXU4oFuNGSTzaIngwK/9VwgJJ8//hwt
DV9KaSfdO0nsPusR+j1+qtb5/xTFEwaDkHeg9lEIOe+WoCD7Uw+IwidFcJg73xjw
O2+8CAWeEJZ6D5j9AzVetoIF4zOBY5rdLeUiJabyx7tyREArYrA6J7lolk1JYf+Y
biR5TubKOxTIqO85wFc7nHyKw8IQjY06LOraln1EpJLwEESjAXJPFDJFMZ2qrFZt
vi2OjdeZuosq1N5lBcBMYybldCJtzMBphBDRvjSa61bQrjmzBPyq0GD+BRki0D7K
sLgsHlqxvUi4zR+EmLw8H1+QmM0VHe3p2pQeCCU0B3XTjzPSTAD/rgVZKWWD0ChV
fBING/0JTnvzQnPclaOT8nHH6EMnZOS/cR5HcOjTpxDeYbZIA4mziXKkRFTLN9A7
u6utZORYkRDw6AF+3SQ6UVpUp0ZRo/h3xS4YDptbLGCkK4pZTJskes8y0Ht5zn77
B6ArRnUhPXr/pkXGOWPx9r2IxmYJXyZojBvpG/SeMG3sZwOeB6CMfuMwlXpQIZoU
/2+Y8QWs3BUnzy3lAxSAvsFX6BOZfJSUxfir5sKAA95E/pnj/MaClNkwMY4TGlvn
i23qGNxPlLfYtweJPZ9Zjjht0XUgI4MdMXas+FQ6zFAohPRESFvYRbic3j3J5+yG
5L1qHg16a8qEwx/SooAUYv1EPzfKjRw0DGeY2SdcPlvwBcmnrxiPdPE6zIFNt5vz
33vVgBEM9PP5xym3X71Fq7kzyAErmnuy8W4DC0wdDf4Cg2lRrPWltmSI7u8nylx8
g8AKy7jvUbI+zUFyrcMR1QGz/mrAZVJS00Dfyux9n/ljlf1UwjbOPNYREEGaq7zd
pc5S1h+qQYiyokrr3J4owd742aRqyAlNpB2GWKiQ0i7mXooEDljYpBcJq3STdDTW
XpOgZtKy+TiLzUHqDMv9jlvDts2WPxFk1L1xKR8WpI0RShC9mQvEuoZG3Sh8ek4u
hwoyQw+wrmoJ1YVV7ZP0nhHiSd8hrLWZjdjdTMSqO94aC5N9KgXO4jmtuDbTkwt5
F5lDeAvT0t590Y44vIffg4MCzzEpZa+tNyieX+VdmKgtlKY8hhkegJsdqilxCYrx
zDoVRVrR8qRs5GnNFbKL/UoKUFx6USVb/qZhcT90jhvEByZsbz6I4pQmn/a3r97b
dxUQzo6jjZaBK+qDzuFLxchessEbq72uQ+mOhbvgz/x+vpVoPIhkgF1tsUXvUgxd
969AzpjAjvxafhQ0pyuJgXSOh3ceu/GhB58o1c58Ps8R0mTq57Alv3FaeBT3x9H8
upgbzkYHKidJWPH4cPYYqWDSlIgjfJs4UShzp9+1aGy1ksRRmjOWb+GwK2aRtXsg
c4sho1kWNK7kfq8It7Rvd8VFzZuVM0HRNuLWh7v7MJFzj+bi1K2iPLqrC+5IX7vA
OFHRwFcqOdyQudvXoylQ/UQNi53FZ55JpWItbxzaBOSeKQHzr/en5DbEB5xPZgQz
EeRQ9a48jQKtImKsgf7EyDDJKSRztfgQmIrIdnlTmxhrvwprJDg6gH3ssU9MwXWn
AX/6wCoN0pCElY2tRlrJMthY84+vhSrAFUWjxm6nYZMiyNeXnemXsgqOTtGe+9Sv
drHakITVcnMtRRSbSwD8ncUVELmdruze+I0LRzimsHKuL1wZYnzzGho5WpLzf7OS
Hxh9na46GA7DWut0RNZ9Ij+UgeeYKCrJTNlUt0oJBvfcdMiSHLMmrrrz5OOeKcl9
8qr4UzXq43dk5p7cOJO04xlb3kDmCu8o4xHv1ujPX8NrDJbhBBJLLZWQOk7xCExL
GVEZMe3MGKzrLV6ejUIHplYvZivOQ2WZEzARyVUNMZ4NhjJMCrqY2/GrniB1EjgN
zjdGrPC8rueuXXY31AGygZLTEiXA1NDYHG0fpTTjVqU9hwwkWYZ4zRgyjqqtZAjE
pCqCbJtYhqTTX6ZsrqthTyLaD3kDMx1ptmxWcjHsSg6qIO2BA+xnBFbORGDY34Fl
S9qNgWEVkA2LZiDJhji/p8pOG+xgn2dFjFaf1f9GYM1ljk3jCPn5tActjQHlRSS4
jMyMrJl52mM1sARM3hLFOgXhhnaRk4cP+lC1NxCu+y6SmjNEDn/UQX104QQeQubd
XrZ0VZa73UhCXOpbyn2x0IQoRerUblZwZUpSDJsj8C6LzVTEXAUV/RYk3wyliK+J
36KzvmbTuv7RwJ3Qk4AwokccxefAJdvieq1v/y/TK9oAXAKieZ71HIyX3gjBac+x
Ija/zCsIun6s7qQvG3X/fGZclgVjoq2nvw78CZrvus2ZJAdP5jpUZyQBFjlmq6ZN
Xf+DVOkoo4GfA2BPzeu1HoHAm5OPSz+PyKABc4T17IV7KFYPQF0LOlLZH/j/kU/5
eUl9vpmSNTRKwTWs0TkxfPrcDP5VYyVUesTa6oZX017kXHEv95WG//Wx4vHMSNm+
AcI8pEXPYjKjryR5djOeWLG+pd5djFfoTaBQ+SHlhWLFdjPCViM0jGjc+ceGJTRC
AhOe4B0hxznhqHp+Gp1Q3hDbACCXGFHnG4q0rkdxBcLg1KHm+viWmQAIbKPfBiLT
O5nS4mpKBq3YSj+OXlypPGlqokOvlC3HqnzYaI1MwVX6Mhe7FM+7R6A//Oa4JDHY
yGt02jq+RGqJHja0Y0IAfgt3qLMHLLRRt1a2NzFPitSPBqsVUAeeSMQV9c62R9SO
EjLX9kkEKrVlEVy4sDf9a0VlUqNxeDSteFMNE1Mz17AcwprcT1RwA32ZeBtoTC0s
lbB0xJ0/KssrdGYHHJyA9HV7d60wuVm87RnZpeAPmZMwP6mbkBud1RNOxVOu9kIO
6FNjWcC/qeKg1B5fqDdbjhM2ZYucwcKvgtOn6YR0faAkUmN9BXzvoAzpQXS4xoxc
6dzB7Ve/YjlRGuqV5+FuwBHo37do6fwBzRgQBKwu1dEqPSZIAV686w7PGwoS8p0Y
TyqSWu2S9xuEXJHloxQiHy3KkqfWvyzTlKz/SxKtUVJUsDdC+o8XSiyJwIpeacSa
DQJnKP4ElChd8ppOdTSDE0QN95agS1eDK3+H9TxJ6Oxp94W1MNWRmezmZsvjP/de
T2yprhkTBiiK62cqSIFrjg7vqSuTnOLtAryrrJSlXbeGi+DqhcZ4jr36Dbg2LjaF
cokKJy7t3ofguk7rIQXtZYjHnBFoM9eZCGRc2W6MDVipe8SPdzjt+0eWyjmz3Uvx
KpBCdXDyltf06Ate4vymvspL+QwTBh6Ywj+fiQyFu3MO5oEQSPHDgbXbH6ls1dmi
VahRLt/EdgBJzWqvt+23AxJ8AZzxLFQGjdv3weUR4fkLIetz3Uy3mlWgM3ey1YSd
g1JAak3kMNERNospbx5ND90aKCL5Atg+ykm/b1OsaxP4NivVDZbaYJH5yBD3yS2L
dJMDXza4rwiTfK2mucJNIwu8AXbUBBQsTU0icdtftlTJO8JGCkVAJqpDjd2Nb/Z5
1jk46PGwUaudxu+elGswjhvME7Vu0gKVd7HgeuHnMvzOM2uq0Or37Q629epEyIeS
5usgM58G2WpV4SnrF9e+i/TCXko/Q8RlUTO2jYQ0AcPV/fqz9IcIXAIg8nfitVAI
556MR9eKXFD4iHuijb2NKUg3ZqFmKc1SOZoel11jirKW8/HKXZpLe2Nf7jhz6SY+
z9piu8ohomVnN9VQijC7RF2vtcfUXtfdjRLab5aYjzg9xVKixKm8F/TV1zGltfQr
MhyWQEKU58e8gW5glogIgMsFpEyY6qzfBH2O8eG0HU6wRZcpJ1cW9pKwPCi8uq0a
MN75l3iryzzQMbez9X4BK4pRy28WqHnTCd13yW1+h7BOCLvBQ8X4ri7OUtSiiioy
xudVwb3oFDMONEu0J+AbzSecPqT0t2ZQ2wKOI5iyHob60RIRGTH0sw2qw2toJUhZ
B0mK/4FrNiJPyYSS9ltrHdmtsCia2Yi2L3itnqj3KjfPrd86epBG7bnymz8wYzBH
S8T3yKH2KEaRHkol4fq8+cdvwdw/ospu89WgHxDz9zQXEv3tNJbfNCKDA/fl9PGe
sOkksiYkVkuWQz7d2CWkHMt2UGSCTKYvXRr3Fh8+ra1FNyZyiL4wbM1zWvqI20S9
CQ8UmxOvxEvSVXn/IyjEXpigwV5bfHwr3/M8Ry0kdyCSiEGHjSCRETQbkZVw0tB2
LAaBkP/tGYtiO83tETwLAB5EcWc1yS5Qq8cZlpQPW0FWQecFGOpJ2FVvWNtwQiDN
BW3BZBCuUG5av9rI1c0atZN+aECyd/1jzZguScrkk6Agg4chnZdJBxOOuzp+1l99
tbVPmtREwoHBDMy9SPatwWl1Wk/4rPTd6+IrPlyX87wWHvqWdX46T8h7x0MpJB1m
yG+Wo3IeUFlKaklTqj58ZmTROLDxdU36k9X91ILRsJfG1vxNe3dZgif52pV2LzpQ
f8u4BhnseTnWJodAI8a+W9tbOBMjjqIeJ9rvP0bZzAbtXBb0eRDeWU2LEN9Y3ecD
6nVU31O3J04uMS/WCfMLI+OvloucNhXOuWp4RP25rPIFW5yxxeQ/pDHNsN4HTs09
rgHXHPZRQKjl04ZUjxum3SdBg5mLtCip8F5bg5lMXF//dJQxPELiJ5C5OdG6Zav4
xtnrhOigUlevn9Go/41Xg+abV7piGXaVY1R1hH9IL2k0Nlm8/mGJNw2Xhv1hWQ+V
DyvslOP9TpZqfwb5HOnecithrwnHeor9G9B48WEavTcSZeXrdi9+mJlmB1DGxz56
NRZ9QIwzpuU+5MW2sm6mnrYtgWGnZht3TjTtQ9rFsr98oiLqzYFINNtQSw2dS8+k
2ft1mT0Iy5eJrG0uhvjmjqqUqtb3+esdPmDk4xxKLeOY7QMLsFhSY8nHM7P5Id+K
C76YfAenyFK8E9dzA05kC6CWV7B0C2toKWjtJB/E19A04Ecttbp87qahDDBzlXK8
J6cPhWiCgeFZFrVvH3kHs6YUHTfJcFAuksto0Uo9acbq/tSkVWKEHxIxvW1YdjIc
izkusft8JTMiRza0/nilGV5MUca9BD0wJtJT3IIBx1ifOpEmWJ45+vUGmjCAVSK5
IYJ+5UzZ+kgS86k5ZOv6FkclhVFt0bOncPDnt0AshlBlBnGh8vApGK4Rn/7YpARE
8zTOzmKei+JN0ofkEawnBkSeDG0f6CPORk1zZv+3I8FwIUBDornyAjjdBbctcihn
v/aeTeX6Wno2PC1J6l4xeb3NUZ2/A+UkRzF3uXDb4X73UI5/rjYqGrW9SU4xs/7G
J8ThHcRfHSFV9AIvwIscR83KipabFVsj2aX/2JygTbMlQhLzEgyPby8+THAuNR1H
3utieZEsB9ofksh94D8VudRjktEjxPTqS9xkKyfMfqxQ1L7J99B3VayNWPRckcNk
1XZ6/bErV6HoC2Bat+iTwyHIWBRnXIl7EdpgDtnJdLh5Y9SSlO0fP8LZ+t09i5Oa
MF4JZiay+d5EW3wQuOEIXuxDbny3XrJbncygz847r9AqT0NqOXeVzPZ3/xvxJx5J
nrv528D5iYOt2MF22CPedBZ4C6r4RUX8msXak1hdN+QHpG1OpwyHsepS7PWRyYF5
cRD7AppbN2GK26S7EJ0/HY9feNgV7CKXMolH4bseUIvzj3dslOSqaWbsq5EZ8GQ4
nrLGPFycEh1mr+k9neqsorBuvhFvPO+/Nt6WBbiKBNwd59EevsXjTUs27G0UQkF/
lW4AOstyCe5xV2njPh9A9SsXZkvpamoCfdMN4b6bpNXJl6k4yJ46DkpK2kxCf6SE
S8htH5XteyLVmr0AockC9E1tViv574Yz2U98hZ3lGtqP/NdJRbEo2T1rw9uAMzKr
nlqPmafI0UygnMz79Ll90YuoL/X5EIimvfVu1usgK7QKhWM9zsrzLrIADO7H7d4h
pgdaQpmFodHWu2ZMI2c4yeU2aEANld9GpJGLK/vCCqwjPDyGbBIKeQqOjeWQ2YDE
Banp9vAmTiSH7mDbj2PR9eTUjjsZP0Nj3ZtJqzL+9zzo4JlDYQUc0LEw5dSyLjPt
tmAyAAWjLj4j1X6EjyNF8TbPF/3Y0X+xmDLzD58E9I5Po8MLzQx4Z1DgqHiaVOqL
sAh+ORIjHV5AlOg7tMK10XRlEaIYZfOId8eiB01shYCnqYMpXORcFf0AYfDtsFc8
kguUgdI5fLh0dnrBDyE2zCzR3c/VU/wZOO0OkpddLqe+TeW9I1ebPEgAZcM9qCYB
YHdxW+vzvaa4dwUe8xwWyTgOc5jE542lsVLKnStkoVsChIzJBm5PO406+quWEeIt
DSTHVC5n3q3OubgwgE/tLh1qxEqi/uxAqRfXFiL9UiaoUZZWu5GlKSRmgEN5hMwl
PZpyXgz+WP09lZoStOzZrYA5LtUBAUWYnFXhOVyh/yEfLvDjFkcHJ4w9Vpxf+Jx/
BPGkqiyYsRMrpGqpOzrbBtLgCl9JhnnAPpCjLDm9zfUoh8ejmq1G6Wie0q9d035G
+lT2onXukCbvFIuyPJ+flNNc5zW/t6RCdPHcA/xWTjywgADOVxiQHbc5MbPdSRVe
zow3rAxNB76QROngto5ZeTWeVNp7+Gd1m4Cjeh43ohw6AIhMEDcCzPStLbUm0ALy
QIczaUFJozTWGOL5ARvul3xj4w7FB2W4UhgCqg/iCv5AxsN4t7Ac0BQJcA7jpAYK
cq0yQUuH1LL07yPQY9sMCiOWFJRy1kkEcpXWvZS706igwtpaCIr7ro2zmI4NOmYF
8p/zisqdTNl8bXHtYLFLyXfjXbEX8A0aKQck6eUNfkoCvIgR7gfy9WdK53IFyJh5
2awES7yzJppvS0CveHB18rLN4llajkhvfaUYVRMEmi8TMdiDwoc59HoD0BpGJhxh
anwfkwlkPAJk0doOz8pfXtpHi+HG3+U/pxD0lQq2R/v2GiRAqIIW9bj/le3b7S8y
Nlg6s2x//lLzZcsSpbMoCupO9KWaEYKO+78+ub+w0Q743clmubIKhdFgTIS7YhQY
2bDA/q94YutVSO+gfkPPmdvOkjaVwVXGxCcP2Ap5ddCCDMDBUvDG5GW/K+0nA6Bi
GSVW+Pu8eXpJf0PNrTfFhm9b4ai6jiJVezqEcgrilF4lYMmQpmxPoN3eS/THsuac
98aUkVzHAQKJGDszPnhgsPwN8nmos5adR8ieEbUcCxhetJ64g3LAsPDCKo7CjAPt
gOMPlVRaOKlU37mLlsEQYIDz6NK754frBiVwyUG/6qpkiPgOSY0zEjFTsmLbNs0g
rAxDwMLS8vtMAwbKCFVDMWngCGO2Y7vdFh175Oh+aCzlYwiIPU/QZnq8oiEtPNbb
i3V1xzCgc+eV5wVZKbTDlEw11xg0VYCUOV3TuI+BDRHHXeaZNNbD4RVDzroLWOJ4
PIAWRPu49NjbGqMdZZlvP/Msy9A+6ftbpinBzK/ge67O0oALMFP9EAIHbMzdFEwI
Z2clM6Bzj4q0sDT8yF66JKEgZ3M/hFkVuS2isb5OnmzbZk4WQCJB0XeFCZfaHMyw
EWP4WKvohqu+vklZ1thlEC61UX53myHErdZsSLU4uiJXebO0lDAuFiO6gWgHtdZN
J/KDYeAaL/AkDjBqhUxjYdw/6C9U6fs96gwydGq7O5paObQa9KrHLcc3KRmIvsYY
0ezPRjVjg2x8sL5opuVLUBX3YGwf/DPjjX6Gu5Buxir9ADwzdAkRIgfp8wQIEuTD
D+waZlLVhuYneSuSkdySt1pqzXSWgtjrW2mCbtBABfRt/13VGZyWwH9r8hTVcuo4
LJdLz/uSVNsid0gH/upalqPU3mhAOIJCvU1hgnY3vlWyC2Y00f0JqxvSlBlmi4BM
GHD4T0I8LIvySHglw5UQTLageaj0fqW7EiU6fb8Is2D93yGulAGsltZZS4X8HfyY
DdnaAlFAsSxsFfV/a0CMCWJXtQ7MnMpyEC7CKHM5O3Ew2GJoq7wzvopb7Syxwft4
qaTiZznSXbB3FJ09NxCzhQQhj2P8km6OTBUAuJCikaViUlb1IVSzATFFeUUAbWcE
z6rttvSxQP+pSLJpljASwbAyZGPyQ1Efuzj8KGAHbPnHWt9xASNCGeleEWjznQJz
3fK+xYq+Pm4jILOTOwtaPETog4z2aR6te/Bl/xrP+exISN1RhTx5xkbewtNxfmoM
Vs7PvXCsNjhnLylV/VpNX6AMBeHBl1lZ3ILhg4aBn4Nve1BE4Nh3U29Ij3N3SScm
bu1/7ugwbpmhFIyCgTK23vRVWyaUHIZbRAYXOAvfdCDzbOCCMfyduWOZFfDiT9zq
ZIfFZiyu2h8cWpgF8W2pFoIgq5D11u2TNM6XfTKrJ1KwElTzqqwbIn5iz0FTOHT1
Ut6JkMQy0IhEqrNunXvB9WTz/O/1qXZxpwO3bCXgVQDt5347qvGOS4qfHoHYkNZ9
ArCLM3qFrCnaBuvFFFvEb5tkcX1aKYNkqe9bwdRwqSCShdyZFlY0G5Cu//qtw1kV
N4z6Xome9a7mVnnJ05BuXqkYbg5G3qEfiWOGtBm9nyQKbfZGObNOk7dp1j/3CbFT
7qpvsKLR49Y0WcZtmBkKoNY4OjTss5ktHrrf3jTJHOe3TKKmtEZSx/bWHHBHDSiG
UB2ElNZi5xBK1wv3YxzBGgWrdej8tB+XQ4GkBxpZSFgLVfhCZ+71D1v9wetX0sQI
S9jywg4AyrRpYGpbN9Sh/Om1mt73iQ48d72x2NFnF7rijN5MONoukcOJkLrsqPUB
tkqZbjfULY7SF5Wg8KsUXP1WvpmwZTeRx80q+E0umVatxP9Zr8psiXnQUXvAnAN1
Fel27ruuH1njtONNKtWxJhHwrVT0Bqcl10k3QVuAu5/GEWbfn5bNDS6qOD0LB5lq
lcpqKKw7fr8woskb8AoXbxxzyneGg6y+L6Vsdz0uikOqjobwEXQgH1kENGlAIRmG
Oc/s5EcJMQWoh/myam7OqdwqtS0Lxtre9ovy1s3EdLdivwo4uFRdx5EM5fWJ2pPR
dPSTSQsPorANDgzsWZm8i1JxG5aVmQZ+vU5uRZqtp/XR206Inkr6aq2EwKFjaQ+G
B8IZlBzU2bkgDybpxCYAg+elC1JlnzCf2CWXgZqliPxkK8k6HDxI6fEPp5dn3I6q
dlWdvtuuRE+YP+pB4X5raO8wFryFpmYJAKhlXkHCTZfb8+E94TR5v/FMsNgjfyHt
/2sK9Jnn+wgH+l/YyrrFTZydXWNrpcQ0IaAijHgAZzQVCW42HBAJzV4LQVylje2V
6IO0RMsJ88ih0aRWQ1OKXpEG7Gmn3iE8PL4Q/9OGVhc/W1NY6k3/2MS6FGuAL3FP
PKWYN1iGT2bQdV2LxJoMUycHnVwbOOAic9KkpRP5EGVnRBCy+2gCociGp37dq7AW
zHb047o++YgCpHijnCyVhGGhxO1h4NN8i550WJ8AHnu49CHTjHERpN6AU/W6W0DO
3UW72gSDVgw1K4c0idMIqdbRa+RTPeijd7ZU1uiutGvZQQX3YbsKkWdIy9poVPsT
JihRU+2coLxeUys1xwKIUof8YilykCSkKPng/FbbASFKox2+9Qx5OmTUjuwnOxXN
5i4JL2vpSilP7WJvBSCYQM44u0/gvC5pkCCrOljgyMXkzXH77TvZq1L70vREFPig
lWzUMiVCOeMOMB/E+k2lqMXXVYx6mccJ9Nxr551cz4vVnVgrx/Uez7pQXKdXCy/E
RaGP1fYDoadmOLYcqfITvAICqrCIXzsrSyWbNCv0mNSOvr4pgYvOs8FMqU5eXZuf
z6+rDjC5Zht9vZfF3dK/k3+grP7+iCb7MZvgMmHKKc2wBycoVldXMKcTDkLunshF
GcOln9SU/lrSdvDoE1pEQZMI3Tyw+ietCV2IiskrUrncXefFlIwPvMY8Se+x8QDt
9T9i9MM5ojpAdp84BzfUu1Pwbi3fjASWRBkl/t0mzhfzc3rnGVTBmF+OtBooIv8A
+9P300huxh+x2UGWyVrkZRpPdIJaA6JSypVruiDMIi/DXBA+Q8efkl88J//7wLYN
ZncdSOOaP4v4Br3tIgPOOlDkiJfe6DubK8xvs3EJZ4FP4E8YNloIo2SYyl4jr6vX
rXeHiorvx5OSX4zXEKN1wHs/Fsv5cJu9d8UiSwZl18zyar0MgXVz6eyuwYulE7B1
+SEGUlT5c+6s83l8svFJwV4Ei1NT7bezDMerythTt9iPNArv6DDFpcIZ1wKG5wSy
QEWiUeJ9NVyIPq2K5l4HuukUcsDjDNRP15oi3xkKWqPRI9zjL8eTJJzslo513/sj
AdcEXbWKykFmZqn6/d/D/Mw5zC5TqOIG/LX7BgdIFl8CYW9EfymDV1u57JMz6uH1
oa34YtZ3vMJeoMLuCJkNVh5RvRdRxpbDxo2AR7sx09C0r5xwK345O8Zk7dbGBdxp
kjuJQn3SP3bg1eCDQi8KocFY8/L3sNxRBse3G3U4O93/Gd2fzKY4EMZmeHUuw6wR
mwCkbSAHVStE36OXLxNJGCw52irE02rIby0jPmP/Npf9xEfyE6T3qxbHtfSQgo5e
AYqhDa2hYq9AoQCTX/oLtDrgrQpO3kU0k4ohSlPKj+vnXgshgwpILyzGOsWO3oHD
tNSoZYC8UXbBNBDY4cSWIdu48m/P5H0tW62x9LowJHG7xdCg5vaLgJx0GO+GySAB
J2vs7+c2FbIhiLHGHioidK2aUjaE/1Vh9sK+CUZ0kHAwb3Pa2WJU0M6ufdcv8faq
QOSshlmkZQuPFhAzkkqWd5fAqZMKMYjNtcxjKdZNw4x09lKufgIv+1YNCzRF6s3E
ERCcP3jffR3h0M35+OD1mD0AOSOJZJ94GjKYt54hcLtDCro08xVQqYzshgCEF7q1
/K5icjuVd/qAaYhPrecEkkoyGOJ6rsLTJPgU3vTGHPDtKRPGoDETiy9NgLNm1Str
XeqjVzGyPc5nNe48qvwK/+Q6vvtRETWey2KvbbS6c1uMngtIwaVGyeR5JpWy/MOD
aOvQoDOjJPfKYqETwSWxpneqbILLqtLwko1FHNA5/WzAKiLfGJaThQSId3m+Zb29
kQ8VTIb9Iet/InQEnvvpy9o/gQfmKuwsV0ey1cX0xJQF/uWlQvZHZXTT+j6hrOpz
RwcDjmAO5u+xTueJdrNZynUdXw5/lZJIBNJjgkeAKxc6Og3OlKy7yZqXu10mtGOq
GNY5oqZpbVwoP0M2Bu5Hr7H1mw3Y7Gx0QMJMdyNSzlY0ukb11A3Shas94xPYUrJn
Ak8dSkZGv0iW9WDmTFwMskK4LczwZLjV9EbNLuydAVCNIqDHtSvrDvLrKCHAcUUp
Mc0OXOWGBiRlxfj1Mp35ci5F46PXKAmpVkxiXOCoAkEZCw6ep+/mPgewkHnvhNy8
kJOKnf/wGFS0/wyBIUHalpqL1kwaalA6QXsEg6ZKQD8IhhQkWTK1Gm6rHKqjC+kK
y9+EgUZxJZ3lJo8gD+zgI/YwIUD0WJFo/E7gBN6Dpo8N9lljYgjIObKCCGoo1XMx
YsLsm8mMs86qkIznrztZhOGKnZ2GIblYINe7AMLXxV8wrmO3WBiTYxayuZZc/Cci
2l+UNSB/h4KsqUMMcf14UrrJj9y6ipmpoEeRbsxIZs+G30OLgGERGheIJybPI3lZ
1aN6y11LkS9i+UvZMvqxcqkJEjfaJhBXHhV+khBP2KtVM8JMNnM9bkQ1TTAOwm/3
PVPn4p7n7kpCIt4Frlyeh4xTp/jUmuQRcfmItAgAanMeskRGXfXMIzPqowX0iZS5
RLLbUVHBIr+viG+KKEDXXrCgHPxigqDE0xRMJiSBn910Piw7yS+xHka7KjXGHpzm
Qlcnev67GGuAt42M4/81BXiKCkx66k7dlyep6BKZ/mxN9Om3Tge+aHtNIz4uRdE8
JHcfGA8CBvBMDJL4/8yWKo5hVHQ1rOCZkZp1RxI+8NNUXmhcgnGIH1dyoNS33J02
o4hBCkDxCc8n8o/nk5AeuXkVkcQQ6NUzkvEMHWZ0UEKuPALTOYYfM5HbOAxzKDQz
Dur6/EIzE5hdW367r4nQtsNRsXlbyHgXJf1Nh0dlWcbKlxHI0iXxD6bZVS/mvqRN
jKOBaVwFlWVSNhe3pVvQMfezdBfEHDtL0JEKXLcH6GBCAaDRj3Id1Wa7HekQPuxj
xm/m9V8VlWGQuQuWWprASlD1lYz5DsPfZTcbfwCO6ul4RZWso7WTwTCdKuL3uTPX
V1qhZJMTGU2fP110GxRWwbZvAha4vfJUXUYmT7jnwfUJzxPdr3YPoTig7E6NJz/B
fIFSOI5s/7wKwVhi64vmNqqjjmXXMivAX4Nv4YYZpVsstAj+p5n3qhoHHnbh/CLh
695lnQnYmt2/DHlrH61yY7lc/ZPNf83URdNokCxiV9Ex4/HwTfUcOolDJAiuxKpW
Kycc7xGvMefCCbAsOSJdKo3nqD6D12zia1ayGkRqeAhjwsE+SpObx1PCP/mYL/h7
Faa6nx5aR16MMVRWDNIrFdJ6PIGkY8uiMZX8PlkJG0e6m+wIsYv8LCqPFdhF9rSp
YMWPLH29PA+Knt7Y4ahbGdZ6jy6ahkVStfaw0wns/LmKbzZx/l13hr9QQXbNZbj5
Lwrc2BHH+YuVGTXh+IOaEtAQnmqKKme3QJ7WLbHeI20OqhWnbjCGeuQ/gTDjyW3t
iDg63ehexyZmnzN1eo/Twi0WfljJGSb0lSyYEw61xqhPgagTJCRteBg4G/R/5mzn
XU35TFLeRmCTib5EJj3kdc3ol6lj+ZR/tth0IG5XuKXbUSgiDX50IBHunWhODuwX
C1NxTCsn2Un3rISKuSeELPtPzHif2Oi6hQts9e+biCb0J/Rr+bdKZHWn33Sc+xo9
cQUB+Injn5KjYyc/48FF5gH+7GAXEdxPx8sNih7eE7zE1uVH07JpFV39Xdd9Dcik
xYL9w1Fr/h6339jOax5DZlQPI7LP6U1zuVfN8Xbl/OYZHshr4YyXQ+xmd27uynmJ
7NetrVg8haKkBtwQRJ+lI5eY0YcolXRsU7JR+Aggt1RhmQy7hg9WDCpqpOrjJUgG
/MhilkfujBZcWU4XyNyuqOMELpPm0ls489D/Hv8uK5czAj3gHq87yBzHF/XYOfqI
502P8pI2AKCgT3w3FAdccvBJKxsml+bhHox9A2I+7QzXHWy6Okr312DWjhoPbSVB
ibnm9IOK0fFeddsR6GP6JTrkYwAmPMimxUWoe0JRtTq7KyySRTXbZbV0YCVPYI0j
ZW+N3MGhYyEVDp0kRfSo9T4uomxNTmpA1K1G+PaPlbi1Jleohr/4Y4ESBIUjMrHK
0EQvoNGZZ7IIb2IKe8gR/bnjyHFVLIfT7zeeUBC/s+Kd0SwMVGXf/MgZ4UXuwjeY
H+eeN8fIZlAIHxWeA/JEbu9F46mJtdnVR9NRU6shEKMImkr1rUBXVQQo7U+kW6NQ
J0Nt3R1DnE1aouJbrAX/EtgUYNK/5GSFKoKAtOOo1x6Cl3G15ICvEIOmOnNtWygr
61axmZq0yqWwzA2w64a1bNbuwnJ2A5nM4MiL1+NrXcfRaY3UYF7psFK9Xo3Rn4rH
XPJOOlmT7OUp8E/5+XvOSdomA+0gU8TSjhR99FmEXae7Ycxq7HrkGlWbJhkVeC6X
bLM1opNBYeZspRRXc+n/84khOR9P5UHYiD6srCc0A5UQjA6vZzfq6QeOFamYj8Ao
Nao36FWE/zNv8nGMngrx1AqIjqVIL57yBEmxzMMd3iYYDLLkTvoHCvvjAtQrPmYl
U/xjc7GzAwGEt/1P0/jYg0CVdaMwK0CLVEqJKPiZTRkAG4Or4vIaZF5RRQ7p2y93
DJuaJtSlDZ1Bopl+4zMr3VHMMSzgU3MGQJvtIDjJYkuUdKKv+km4A8OGUzhmeczu
IbrQoxhAIQSg3YUwvZ3mYkHqC161rUn7plO7bzna/tk4zMswNrb2p9P0NmzVd1b+
TsfYJZJRtW7B4/8WjMDFJ3Z8wTzEKdU6pXnrnIADHP+IWfDzZgfaPUqBNXyhSNXs
XWEuiUzvAVZr745xzHU6oSJNKnesL34672KTgYmnQ95zDdSfiLVi+f3l0exj3XFc
grwl315/e1qo16p1PgEURujpQFkEGlG01vYTsFeRnh7L1TCJep4Gc5CVCg0pP4K0
IidUTCj6NI2Ys+UOQvnhQa1IuHWkTaE/FSN8YfZURbBHRG+k5s5z3NAmYVyiccjt
W1ltveRDA7d1E/YHfoIFB/GZiqjO2o6x/3IfslxVcRWoV74m4zkkCIA52+yyIYF6
DCLa0ulkmkxtYBiketbEdfJjK/DelgI4WZfWuVPU7sA7vNfC5qt7i8DIcg7wdqcT
DpJf1SDhE74gMlJ4ktVkv0b+QclPnSLM+Ql8Wur4pGQY6rml5tm9G9vtdeo0srfK
6nDNlV3sBA039S/oXL2VTGxN28tyy2srh0kD7k8aNE7OybgNbdwY+tZ0F6TFtZJg
vWy6Dr2cQWuTgUWVdANFr4X4agRswDSKBfjljOn0lgnJn30PAITwTuMQ+ZYTgiJS
iw88F7D3DX7Fhi+rq4ztM3UUJ/IZveFrGaNlpUV9tTfCfSK/h3eOP3IwGa6Pha8J
3u1Ijlxx4mzKgN27Fsiy15xEiovgwx/kk2f4yBgQyj91/fSq5Up5ttb2q3zR4YrI
dANS0fxCR1GfXbPzdzRAnUWHYFNX1yr94Chm3K4bQwSrTtoRbOeXLwgl+Er+mt11
TEFyBHHGDTjy6dOUZSoGELV/fWMPFZwXBEUcWhYsO+XuK7ZzeNzXcnp3M/CoSKI5
u0UnUyWnB6F3TDAJxFWBQMY0YBilp5dcFg76ZZ9DauOcatr96Oe3GZOXgqffnXxk
RORkGDSv2xdMDvLLsDYZnBzvCuW4G6u2/goO+/5qjqPBlcEzPfcMavqOc+0/lUQ0
3+FOwfrGxcQV+H49hB4fDQxmYxWd53qhcVSxLmlkDNvt88C963T4NQyDpF7i/AJh
G6QHoTur8rXScde6TNoj/pFJVKQi0uh7LFpXYwef4nko/MQljkuJUiKHv0p8bmyu
EcbItsdXYLvduiiEcqu/5zu6KAYL5Ec9/GK4I7Yd4PNoBCWOBUEJx32PFqZCfdHw
6BDdS7MY9UM/WtGD+eNSA0Bmy+8YXzgEjElo8RpMM/mah1F7kVEWi14THu2CI9kq
e9I+khfQ56a6XA+o26MqItZtVU8a8PRQ9fb5JB3AIiX6C5IyejJCXYrL+NuWuBhC
uZCDYtewpr4WBVcSFGin6FNcf3RNnASejgquoZo8FOzKLGZ1mHdVSvhlq0KNCCW6
8GMDVq6A+FeuaULbvyo4sVX8ycbnBhLvsUq4/IJ5TEPwtQokaM6dVlvXYJf4m/zd
KMm6dTMRvarZPeGS8jYQhYXX0Qx9DXg5jwOZGIpBEiYbkAY7EKlnyq7Twh8HTVje
D7BB2i5ffOVTthgbJrctMLJjJmvfn7z8apQtSqlIV5mu9+aiJ8YAZyhTI09QE2gI
uy1QNPSFuqmHajajN127i9uuTMSO8b2sqyxaMGhtL8qMCQphFXhBCtr2CgED50ph
pSLeedBHjcm6ipeTqnwORCEqILotRwK49hgA0AOQwBUU1eVkLobFaPgjFmohr8Mu
Vz+4NMBJWdg9YMJ6bnOEX8cJbyaEjiEuvN5Tr2+TwCHaNg6lchdS8BdQ2TLgER9a
g+iziTWWP95dC+Awfo39rditVEviTT5W0wRIUHpaXkV9smnCMMN/HTIHBeprXT+a
gEjf2l2O1G+on95zJNRx8WhgTQ4ncsqOV0MX2g2T+Hqa+6yRoGqobVedGh8mUFNO
P4ADFAGHGzv33AnThmhGXV23I3Cm0h/FJJ+csiHMieGML8m6esxo95Xx2vBaiH2s
eDg7LiTjS6YXGaLnWUifDlRedUo9NLLyI61cgvg7qB0ThXm5mVEhvaeHMsoSVcn6
NT6xs2qiqzt5ym4VyR4scOSTuAglZ76/cnEi2lo44u/JGZSu0SbNA0lhJ8XOJxHq
M+NiaeEpXqsNiHXnz6hi4KCxq2WgNaEUAacrNV4a+Uij9nxy0vGVE/9K8+Bb9yUh
RrkJWz4v0Mc8FkBCJU8BTYoEeXxQX5gmBJGwSfBMUh8ljbJg2jupbycrx1IeDnzu
8LUbe3qKnHnblr2Qyazv4rz83VfT5u4kHup1mGFwgsBnsFW1LZLgBjEMOaIZm2TJ
H1Dju15bfUYzUzHx0MARTNZyZDgLAHOmkMXN4f1GZZd25jABIMv0chReNdqwFO5Q
EKzSlVAPtU0r5Ky2D7ApU9/AbjOMAb8ekznoFNLPlweCPW4bSEfgQ1fM3Nl5lzr2
sIP7P/uwuNcefACjxFSocv/IewQ+xrTS/no7Ti0+tIyMaHL7YU3aA4DruhuB71yG
EH/F23NV/lZ+KnWF/hJSNCXdwA42O3RO2+8yfw7Y1JlkCp5PnhlRxQ9g4APyBjYZ
CnB/xm1M87hQIjdWQetUMvgRTA21NoZtfzYgapacB6o9ohORdmAEs/Hp1gv3L+qF
SutFo0PZeJ94TdLEMANOqZQ5lODIWV750Z1NgPX28KQOGaxM6FIPZPuPOI0KeeWM
eHRTLVcd1xbX/0FnbnmWNjeQaIdbHgaituCzoheQBJ4vXzDlB5XpNP6P7+mEJzFX
uF9wHl8x8PVSOepyet6mfTAL+JBin7F1g3tuh1jfd4BW9C50YEzbyjvsxUJiSl54
6macRKODsbLzou//oUMz/5YeuoXLUYmmnih0WprKO3JXuOfLKIJtybuHev5CaLEY
BT7Mj/uPPzNmGUmQ291hrFc7SQ5ONacfJ3rmm+/1V8MUAXcv72rikQs3MbXRscjd
qV1tBNLfTeiNtXxETP3yCPNkIOPWf1WRKds1WC9rfoRTPVP860YV38PoqkzJwrrC
nKXAi+gGAar9Q01Ko4a3fXw/5tt8RMv4iB5dvhYnDaKkU7zLtrRQS0IvS+o5G0VO
fxT5Gg069zgf2ZAVE+EXOZx23MlPRln7lNygX4DLM2YO8uk8yWTifibDwP9wqMPb
6x3TbxpQn31catnnKl4gkTQ7Fi7ss8tkKinRXxG0n6amWJx2pglFNYbP+Cy3iixy
wtootQO0lFFIAvuYwf42gf2RQvlCq6/1AfYj0mkWKYnEgLHySE2FmWBEKImE0DkV
n2+SCORizDa+LRebS+kKWX0dizCG605wRdpI2T5/xWN+Vb3ivR5ovWeNIJSKcpfk
T1YBErNMawmj0CiFBWncU9HduV4p7GQljt43dQ/G8++GXZnuoDeYaRJiA3qqsVdV
DDQX3ycHgDDm4CqByHGTew/S0m9kOfl7+OulYF+rspTHv368De1DuS/as2IrEzgg
j8FRd+vxkYSDZxv7OBGeCdIdLArC0IZZ/JXZOd26svwbjmnMTMs/FHWALjGptrV2
B/G2yWorXM7e1qYYWcYqUXGmvEfTE0DSUeAmnGh0Jswij9foS7DLj8cUOU9CQHmI
hI89g9bro94ee901wARuI6uySCKK+CKDYQM+bDdPK432LVQLuy2c1uB7yJg3+M1m
R88GZuokpjiZ/BYJjyovONxh28QFa/e+ycMNxRuXn9PIrgsesthdjtFDT2gVtdrN
4S+3m5n64iKK7nPBQjut8txQSon4PTxUB303Xk/sj1H3qekOEgmScFsTmPJK8Dlu
b6ktQ29kImgUV/PDGZwEgp/SUq3E0q03fYxKNgDIhCVAWjTeN8s1bXba5fuhrA2i
InSQJn9Gpmn5cIVT9I19ku1+H5XWJVeMe7qsGXWac7+PQhOgItchtbWGKTvq7SXo
/hxg/LuX658ZkxdYn5HxwOXwg7YhZq/PZyNH2r+/kY+/f+k/PY58jcpIploBYOVu
uf7U2UQKENLIx3nhwTfC5osoHjm+/QXuYFDW51UzoD3Hi4ULMt2F2lRkf2mMRSHS
K8rxPj3bqB3UrAqdwwhy8vjqTuL90+oJCGPSsixicPx4D0Xwd4nxXPnzy1000bQH
iF2+BYiDmixuhlrjYFCW1Kz1QPKO9yYIH5OqPmR5xC/72C4+lufgBV0hQGBlaCIH
g5Zg0RujzO6wApdyPoxpvibHUhmQpPH0NRqurjxIIfkbVoOZEe5X2w6515j8Zvyx
MfYwz8oCfEkXghx8+5eO000uci6rw0wp9K6ncVz6S1m1fKKvX66P/78lbYzSKKCl
cqJobqoIDmEkZCO3dDP8q1l/VzqoOOGSok1AvPhuDyQx29AYmRsMm482sMn9snmc
+ESbu4a8ITh880yhOJh+ypsX0gfiUfoJ45f9BtZ9fYSvOrN6AyNF9D8pru/lxFSk
ricZROz9q1H+TvuYvEyWAteb9mEs9Ehuo8Z1sJJlmh9DqX3I5ssjVZGXwhu9Zp5U
9h4LUh2lTC+GNFCZ9ZBxQayPIRyvZnFl/W57bB1iKPM6chkjIz/GENDc3LtE/zYM
nqFUBMrAZ63Ly4NW2gveCAs/PZSTKT+qp/np0a7EPIRq4YFsrRbqoxCKFWzh2QD5
05o7QY9A+oiqYrGEf0f8CJZEJlEMNbkN0RiVrfPQCcx/l0Se9x+F/ho6G3Wg1j5t
Rt1YSi98nR7xkCO7qp7yRQL9pYkjIJC0TchV3YN/yZcm7UO1G4Y1xNOW1WEz1+5g
exyr+xs5tMHvEMGL3+uqw1Sacb1O+zjAVwqBpxoz9w5I5i15HboobPlkjOAlrKZu
fK8mUbCCMEKhyRcjPJOM/KvBvMvTXyzMPDoKgaIyAl1tLgDwmBmOWudJct96Ll0o
U6MI2ZpW60EYA1JzIEhT51pUJgdL1AeknSzxbdUKAR3ILA3oKKJXePSz7Da3iDNg
qlwiEcAHdR6bszjYvl0/O9RK7GNJm1WqNaPExk7pef5hV673Wi4iPgeENgnjaclM
7NskQAsgXyiRQ5rgd2ANTfGI98QVbz7KiGfFFkIqWNRKkUtvqCUdQZE272SMQlq8
bNG/q5m4bQU01dYgD85rUeU4QqsWvfzM2Q44XYMgcC7A/PR91YXcMrwmIS7UqpuS
dePZooeUraC17DEaqFeNTIZlOV2a6AghpAUBHVf0iMb9VXQ8WVTB8COLQwbGyirJ
Um8hQwG49M8Av6Vv16ZJbd9dzGclZdCJO4NDugYcatkpQH7cOxd7aR05nX+9KdWo
XN82YXeilI/nM9sWgQWE/TZlpf6W/4cvsDbZ7VMf+53WYrWljkjTE+WB7G6Lw3ei
9kg57EpcCQGE3bfJqrujcdM7E2y0tEPM0iSyRHAaIs5NjxariSYii9tGCYoBP9+B
qi4CANJfxp3l+TKlL1stTJP9+rocM5CwzNh9Ki9Z8pGPyJtLare507JUTPCTc1gp
QByIOeRoj5XkJ9AedDWBvsK7aXqP01Yl4Jt4PdbAYUUV3JXkqz07z8sYlUs8aU5M
F+tGMkc6lC2m2UBIaODEtCViu/AeQGvX54rzYTKAahCXIXdDwT/POG7+jZu5YxFi
x102g0SThgh6E5zB3d6BFhm+wYAwazILkodlYX0FewHaD4jbtMgv7gf/q3QXfiZ5
poSsRKsAmrcQXDtpK5j/EFREceYfTDNGX6uzOFGrs7tdK63g4HnovMofWeGPZzQ0
PqIaDKm3FBeaAEhnmP8B5fEzwPcrddKjvNvI9xPdauw2v1Xo4bMFVSpNpqWjOZYY
UMpdBnH2k0usfFdNDikVnMc8x3c55c3OjCrffK4nDc1GXUjX5YGYKglI6yT5rBSC
JMMmi181bug1TcNVPSA09HN6pglyxXR5V+1Csm4YsOkPRTJhafOF1zEW39R+5QoW
Xwb9XSv/ScDc0kLV2S84oNcYgK2E9p8f+rrWdYgKtk0c8BD23twk6rJoIbAaLze3
EAeuqJwx+hJ0D1Tvph8XsqGhkW7iB5MIve/kzQ5S3bpdlcnZODc71EZj1dW3irtv
PDbaY0MND/fRKp/MLZKxmhE9Hl/1f2mf6t2lDMFpU/92e1rEJ4u1owv3sMuuz/+M
sNJgJguhPfDARAwo4m3mYe4it0/fScHNSilKL+Ll2qDdrKPcf0FRBj0qaEesUCwx
4suxsp7wxWoSECNhJPj+RN8xQ/ErbIZ/X4r+lk/XJMZPR+Vj9ZBHaDRpJP+F9yao
+skIdY65NnAnr8hrTNdLml80gVxK+HqVGLQkSLvONllH4VJ8hJo772zl5cD5Gzjp
1zxwBK9VPz7C12u9rZQs32vCjk0+Mkei33fOjDl5wnzqJisKrGgVw1U/7vfUhyUn
hpHCd3LHgRzVZka1LBZ01cQLyaBtoRts4KCimq93aV6UzFpEnwOyv5YFmK9SPxSH
izWOogo8ne2/DL5EzRrE78zHMVqeiVmg4U6nA/TZZP3ijcLgtCxHCb7sQUr46DCw
0AUJDCeqyc49keMpJ/7QW4SQ8M+j9ySFsnbGE2IKfk4VAp0CIjkymR9tzzV4gfKQ
BrPmMA0dOGyjQt6E2HZlBDBFMu2UgNHxFKw/X5FHb7SF1zp9wsw6HFcvf1sjq9xV
Yz6e3wYqkhIboXxN2rySfNYuZWpEDJKKc4G8/9pOujNSyxVegTlg2MqNqI0nBvLl
ChpGWz2CY5ug5OYr8fRDnzbrbI+Sj6yquDiA6VwHM7QJqWbN+71qFnNp+82Cq6Hn
b0DUmhjQzfTQQHWIrPskwUr4i5FmX2yerfaJAioH9NOUOsPFwQfNdUha6pV2eUx/
VgS3ADjocHqAgrQbn0U1PgtQf626W7rgw170D2eIh4veV092K30uRYT5e0WpdxWZ
vSr6jPt6u26QcmFpxg9Acg5X139xZ3w/yxYIYPHPM+jbOHXPr2XOyVt1wolAnKqm
XrWASVvTJ0bzU/RezQgKrlj6GoDpMk0oZvby0nK7meRUKcl8RcCkMJ2cix416Ccm
/qJydMmgooo1biEzzdlQ0xZ/grz+siISxxtdpjtbOGheEndiQQndCPQUCKNpRKQG
3pI1qcKge7Mn6/D29Ighg2rJNHZX2hAoARvan9csrrlLDq8Sowm8QuFYAxYzTqSW
YLQxOdyrvYt4jGUdrj8xxtO+RNGl+ar35+Swi3oga27+6XaQuL4uFxtRscbAhtou
WdUYo6oeXHmzXQzjc70kEXjIlrTUWD+r3mKA6glq77EqMyDA4bIwrgjYfnLu0DnV
qxRvXShNkDE1LizaH94+zipBRkharU1VdXmEYMjcoOwUkEIBRg9b/6mPUiHok5yP
jbcjqxBsXJ6yS51F3nXXhrAbRsGDdYf4H79pvpRTmc46btQ+l+Gi4Z5o1BX20FGn
xD2ydI+1RErMq5LN0o0PN+/UcGzzTqarFUg+JoWLdq7pOJEev77UraF5BGc0r+Uz
CGn7p11W2BH5qwx5bcRbWZBpDaDlHXMsXm4laMU0jCkv7+qCgaiVeC8WO50OORhW
sJvLJsPKbP7Ch3TfDnSwWMWrLurBRVO3+B6FWST7+nAjEbTf8loNqMqySp571jt4
wWKwuR8PCFvjJCutEiweYwGhmfYYKbJ60KNUuellmuM6Me0uW2nmGd83pZX1QxKq
BdHUSGTq76f0SqrR8E+ikNPfA1skx3a9pJgk5nql5pcsVF4E8Q8SVBXUTo07bdaZ
FYpIHz1bXTnb6qQaQ5+0s/45PIegpB7J1riWItg5X5m33xjGSlvto2E3qv97kWht
6QPDR1cs2d2pJDZSdDWesD6ZVJ6c5F2ZOYf8qYbrj/Lerx5ER14An+NXq4JDjt/D
x7xoDBn76tmsIeYqMCHzbyn+Dc7EAchL5Q7qCLAKT8rKw/6p22RC9aQ6u+hbI23Z
pKe+dUq9EpjnIkE8jbRv7Qnl3OrPwowzKBkYRy9he0OiMpVIxwkLJk6RxeYLdHt/
CyE9gh7D6YORsvtZZ121Yvf3JOEanq7AtSpT6W5oW2hr4Q7YAuV7KXzap4X7ND/M
XmEGyv0e62CyrtjZ+bePKdb6L7AQbbyX65/Xa4ErnbdEefnDRdgghYe8cr3Yj/hY
zWJEk8V8eszhyyl5Mpn0/yG8BB4ItX93XJIdnyWHQO44x7ychx91ofp46FUT/m2k
fmTBrkvRqKbAvWm+iHks35psO4K7lnne7k88YlBgHztsSyJgTi028Sc2xbQ9x7j5
DCafYVT0zSTVutD73QRma25umZDgZo0DyMeoVcizsfVNrkNT5yaHEVMr6j/LxD7p
eLVVahDInMrGyM9sULyXkDmQ7KZoxX1crgumqivao7JSNUjOeBGpCK73l2kQUkT0
Z7AHnIMbvgTeeubMfGBLKMTfH07BEkD0cX0/peJBOYlx1zw0XVxmXpzARoDp9SQk
tiXLljxoxpXK8KZ+0KQ5Nl+Q120M7v92w8kZSlSnqPjdyybCtA3NC2Atxi4lGTt6
/lGsCVjEjCo/ULYv0EpiDTlLCIQQ+4upcyHtcM2z0I/1TgoMYb5npK9Encn22edg
GeKxQyRLey9mD63vqMBkWJjFRKExzn/15PIDIGK5rWKu86T+B7lORm0m48+g22O7
/oxZprg5A84wNjJUfVkRFMpPoajNvqppo8iMdlZZEfX4mJ1sQ6etWNx//Pm749Uh
LeD563P7Inn8zREGooCW+FXM0RkiUT0S6xN1pZNxEnwcVqWh923c/i+dbjpexqo3
n2SAVRZroXY7QuFRvygAc8BXrMGiOFaGuYGP88jI72y7IEIdcXBPxRQhfN33k2NY
JCQhe9VBN95CLYlBhaKwwT0yDyuTrMoILZRyJl+XDsFUek7ckXM318XQ/tuF6z7n
pcN04g5IaUodemceRUP802dPleuaAsuE7QodVj1O2n4j+ZK3LizpRiTzUxeZocIm
v4vJyCAdnwVSoNzMdyzV7Q72hlkP0VpQT87rDTW2yJHpOkDQ+UbEWGblbHMmid5l
X4zbYLoNauxLpBOzfDHznDsFYxd0z2TWZFmez4wRtsOe9jxGsDlnuPZ7jvtPw2Ur
xP0cWWcn14CfRQMPpaMbiIL8AsRfJjZHHytLa7ixGgW6pwHMqs4c+E2rahZoJNtC
VJQZTP/LiFAQt+xg946cMA7cOF2ypXj1KdrA1iMxUFU2cbcLIoOeYv2sYRkKCmBu
TTZ+0MIsZSWOv/hN4kpBkO5wqDvwVqQ39eYxwtUWjiAEoW//yE8O1yKn8pN27G31
OIa6ylFYqKjhIjRPJbjF61deAQ5OzmXcY8YHpTSau218frIEKmNUyZ4McF8uDzbk
2L2B6Hgoy++v4a14Zng3zIGYOIktQfH1NafHyJE+0LuPBmF10kTdE8hLeqRnZxLs
3wNVqxHYSeRAiz2IJ4vPlVYeBSCg46E8vFDmiHXkAC7NtZIUdq81FSc3XorikFAp
BZvQ6DouLSJpIkW5YnpsCM6498YOjRjVbbv216MGjDk/49am/s8EcB60stYS8DI9
9XMREAgLmMi+MwGTOI/QJBW0/+HWAFaL3EJjImVvCx1RXnmdYfizfeLWb+hLJYMq
UKeCZXUHWtu6whr2eB5eHtUPsmeiX16ClD20jJ3xjdzbF+0TMXz1218F1AfkZDAw
iqpTaSYW+tKaf6gVCACkOZfH/iTIHaF/WdGmAO+0w6hGyEkKtDTE4tB7yE7l+f6n
rcqYaXzvxh2dNd1AZAi5XqzpHAJGJvXxVZMMkTeoJ/lPjx3kmXbmOJpZpxRwRUu3
LLtkFj85C+OhSQE8DkDhDfOt05ECQhVyhBCxjTeNd48kE/RZu8iEyXNBtWsv/P0H
ofQqrSXWNNJi83rAObzRzLBH7gD8q0lsZd7EJB+4KFYTJSfJT3yCB7w0XPU1xxhI
M2C1KxbmpZ/7zlqSOf/qNF2AaHl2eFDhLHgVMofyYlw4mvWtUMw5Srw0TqPQuXUW
u9FpJT+S3GiBiOwIAWpErKnRvsTQtWcMik7FwR1oahXy3WVDpOAyBDu0QnMK7EyF
p63bvL76IMaJSXjrp4dv0O3zKCmkNjcmQYwmFNjCozmpa+xVG8wNfhz9E9Pk8uMM
W0xG4nlLdcJP9B+tvWMk277ozgjs8q7Qn02QfpHLvZesBhI1J5Kt5QaXYFJUOzRX
kYXQa1MUor511AzQInJ3ZPNMVXPgwrtQTNATBc/3jMWVCVMFQwyumVgbVg/z3hzV
iVLIz6WuSFtxrkErZX4+n7UkS45q4/IJaLFIshhbhHRF2no1SyA/LTbA05UMHCrv
9FWokq9iWgIqXWoll65cBvdWoeajsEygrFoDxiVU5IGnL4+yae49aREwJtxDT8Mz
FvYYqKh6qCV1PYMbI9R/RyS3GvCY2RQS3Gy9jhfp5nV9Ik0Z0bVOJLwIUEie3c2o
VFsU5eghJhYJ0obQo0404hrv2iUFzGsto4XuR4hNILHucF/1tBWXbzxel5h/w6Ok
VZ5iuzf5FyYrKVBX6jNqsvdegRSQ4ooh+GYzbHDwmIhQrfJYikbn2e2rYeq2YDCy
FsBbA/uBLIVg8XpzQNr9UlqOpJSTwTmDNU97+udGKuY7BLIVx/eIG/42l8Q4XMJH
NqE9kag6ScQutRyW4BhYlblv8i8VXbWqpNk1AndyNgK/7/B9r3pUWSbt6bX6rwS9
bLvScUuhRqcF+aHu7rOCRytp97AnqOFqQinFenRXXf1cpDSa30qHE2db1W8eAZHg
ZfMfZyLMbdVuKZRc6ZE1RXQB4F6lPtbeFF68Fwg9nNRiHGsFcqH0KzHkfL90U0xS
SNWfNrmI6t1xRvxiTpI1cYjh/vIlDM7XAgxO6PTpJs666phTZOvg7EUfVccXatXL
0/kUGI45UmW3ttPqWaoRQNci8L8gXK4MLu0JwseY8qq9Ui4CQI4Pg5DRWO+gac+7
HiZSV/i3jVn5IM+HR74yEPDvee5LkG69ScOViCn3o4dWGBSpdB0bi+gssYXxzVUe
bz6cCab1IoxIGSpIKnrl53Mmj3tc78TAJ5UosK3g5lCsq50GsNcSUqWAZpAC+Xcx
0L5BkUVfZ8gOBEG1I/YyxjOq7i4nxKZMorzVUoPVFuq9ltQSTRGTwEPC8qs6QPdS
rtESQPYfi7xvYAMpddsvao3x3GxD+bnZOsqmLrkdySOzLaQtM25LgksnHhtIrdWn
FhDD564YgS+LkMUJ1GnPVFweV8o0/ZmXYIToa+VzFq/6J9mpA7YhmDFbBtpddIK/
xgGjY8odCRQU+XF9RuUIuiMpRtHlPuu4uANPjESbnDiTKaFJYNYyIeDtU5IecAyZ
BgC5S5kuSUlvZXOUOif+tLhAYVIRGLEJ/ihPOXImlzKD+D2n9PluEGxI5LSNhNYV
XBshUvIvy50nRiSaL1wWRN9AoQgNEEgV24vf/GC4AKNaBsXcodOeSo48A2E9tl29
V1wlpnlZjPRFq2GR6WZ5i8+8G6BoRBUVIg9bkWwzZa/BawhX9+59tRoweHL7mOLy
48fjrUnt0ZNvVMeNtHYbD7XcZJOAfwj6MFUSIBTvf+HCIUwWoRKYmBkRC30we4Eq
aUTH6sD1H242X40HninqhznNtXG7DTxht9lm4e2/kb9ZvxkQGaIl8/UqDyGF1Eho
cTwgTdJyetdKTMa92+0CpeCFWUXOpfJ4BqHH2YvoHtaF2IhXrAUoCHe2bYpXt8LZ
+/MLPyaTgAXgrx+5kHLYPEpifl2qcgFG0ENzRKiA+DWr0CB3IT85WiB2ntDG/ZzO
eMsPVUY0/CVQltKl28ChSejWRosKydSjay5ROKad7qVyvROuGpU9t5+yYwblAuQ0
BopX9oyvZVbUleKyN31jT/J4mbQQCsTQseNfAMl3gDr0THncqUZVJKjU9sqP80n2
DbTWpkzS3m73WBMySbQWO66N7UqK4vWu4EZnWhqj5AiU/F36XkcAj0iq3LSEZ2Cv
IdXSrCOF3JzexWNuRrpZCvAR9VZ55YFOfURzt9kuEVez7pyaNPRcJlviTonriBxN
r6LL+H0iibAxRuzfxrxfz08pNtd7KhBP4tT/TuESzmj98hgXGD+Y2mka1NB/Ncs2
klQCfe4TKqE6KuqWRYm+eJ+vfsPW/KjhrLGCyjdxLyEgL6j9DQmZKfBwfskJ/Oj7
9FsTE4bi/CUGgieAB9mK6zPGdV4N5SZdsVLnxsxUSimCHZQezfg13SRmuPnxT3jF
Nh55WHvfH3IyVWO4/jOOncZL/u94nkjIsAVshfUwZFHwxiywXaNoMfoRyn6WywtW
k1Oa5nspH9hpo1Whv5Y4en+PkYvk34gip5djYBLowuscIF8XeVV26rqWtN8B6/jS
3NBS68oVvmulE9Fzy5uUVdtDQQcvumFEHnmncYV0VlIehyQg1Nk/u4Wjun3zaCht
l0bBLdELXCU4JmnoQ0DzrmE2nXK6uCs0+imYbtcAOxQyuLhX1o9Tq5VmuEnGMvPh
FXtqzJOzD0QO2b9VNJMDU6Mpu/uzd+9ZPk6Fyx1WR3Ov1+RZtZojCxEhUH8ys0is
20AHT/6QPVfEfmHgOQTIZhcStpHszKE+0iMG8B5Jvub0bwnOA3IuxLHhHWAgYZpk
r6MfHqYtgidC+1/hJgoZBPijxgsk1/rzbJhxRVPUoDufnuozH2RLNFIR56IjJqMV
ZMWEftBypW2ecmJtvtdEqlhZNAiDVgUkzfiymnqWOI1ZASDtK7YZnB6dfJjBfhlY
HOuzmHVYQw+l+YTn4P5ijllLmLFk/nvnn8fx4Xwyj4n1a05Ybi1WrhhavVslRqSa
1mIbD9o5hO7a5x94gxTK4QZqW/8ONrnqSgQg0EUy9y0DqOM5ZwT7lMjV5dPugIcK
afAxM5Xp1a44xb0OpQ2tS4Vy4GYXnSicx1wYtIpipHIDxPFehcvRlk27+9loNIXf
mP3uTRERlgjhDF95zpt/aY2O2LUZR+6MtEV6teFwuPfzIcwVq8UHW7XAZ3sjJLH9
OOh1ekGrAFrxGuH/Fs2XbOqO7LuMGVk4cb4FUQufOpii8cK2bW1Ow80+6rp6RcrX
NJ3jge3VXZdlQWApgCApe5TQk8yiXJYcrDKTQ1TIGUGgEWe/encxWXP4lI/w+2/r
mhC9Gdn+Qs3hcyB3TNwdQAdyanTvWWMHwsYysw3qdgZZxi3DWVx/c4Ew2wJGL2vK
A2vhSD4wyeCaV3thBkFhSEnzubS0HaK7s11cN694q0Ez3DU68SItOomzgcUgay93
iPoZC/eMlOFzoor4p/mAjDYunOlsWcaU55psIQWsSxp5HI0Envr7A1+SZVy+oZOz
q8q5t/oD+BeUDsZFwJezXJX6PlH9fwXHylINDZ62FRvG2DXeY/Evpr1FC5GdSJpR
2NqzF6hQqMNNUdmIVMaUG6HvaQRDPspNXrh9Cr2APd0fIHV6D9x5AvFwqoF0942X
DHeDxzpHsev3K2QxH1cEozWwYiRchiHxSXjunZTafr4VGQtDDcrwQagEfeX7d0TD
6xtacmGfWbtOfa5Q8AYdOqtH/bZSNkKzGfrfeW9qGyS2o7xIaf9FjPxRo/fg53MO
3b/IhMlxNsmuiwik/n48FtAGf/hsM7fvranNYPKxFxHHZDjUN+yqTky8/vO3+MeD
Su5V2zoH3MPqMsZCbL5iM39cMwLQpLUJVbpVd1iIJ5DYDHU0tD+y4WzvD19IJTid
jCNnQ0s9ZYelQ48MU7ia1kd6XB2eJBCliW1JhgubYsCmHB8bt7VgDwx+WSwBl892
HccotBNx1vSbp9SrPC7dyABNcWJFW4xtdES6qmt7A/SrTuPfh+51U/FY+lI8Eejw
yR1Yd2Mrb4g26A27gm9zn7I3jSdGcYD4KZ3KG0yO9gywWo1quNR41Dur5HDg9uKP
FRV5NiBeaPXWCDJdDkqCT7E4IZA7BDr0eAF3LupzzNcm3jLmX+wzBWjLAA7T5ONy
Ngdu/V9nKs+MIsEB0oZAPN9b6RTj/yM1aLG/vzd7U0cMwmzP+9PrixNdsugq4IhG
x10LGRIzyvN9+PENsVyfqJwYLq05+lna19n1IC3RVOMTdYrybTUisk2OdPFbDuiQ
vXIlyVrWsSxLh50ImY2kqHlisFA5whz84Ps3viqYLQ1/ZDZqkdwAhHvRJvHs2HEZ
pID6jOuA6xByPLdGpJRL2mU+uCq+zkcOqcifx03DrDN1JLeDJxOH2KFGqcQk6J+j
t7PTamCmPAZ0A9H6QFnqxGDjMHaFeHOdVoR6grX7tjjGcMVag6zErt5x/jBSERfD
Y7lkWcfdSd1ny5qadLDAXlLJH4cbAOv1Y70Xm0UndkUxQvouFy/KoqKdcQ3fXkn4
8RfCvN5RwnuCQdzsvq+Uu2EHLXgvEoaXl9Q+Y1K39h9SKf7et/0RahQRfBPv18Tw
2koJ5SNo7um1CJmVw7UBwgUCl59lggSVpsEoolMyYs5qgC/mEuvmN1jZzuHymxOg
MVSPoQbikdAehDQ1EMAcBIXHwWuVIPE7xRO2xf5lKucpnTtiKlTvPzLrHuaBttLs
c3KHPtJl9faRC/LwBB4Kze3yBXKDIAglgRzWjqry+7odroKmkX3N6Q7Kg/xG453M
VUMo0vanZzGh08j/GqLhscE5dWBCF9TFMoWeVzQbjWRtkZ80uxk9TWJc32/gcRxj
KC7vyG2/fhM4+W890iQZHegPKRrk3+f9w5XKRA63Kh9hQd7L8Rq9apHsLIBXajMR
kqKep4wNVAo3ZJDgDsWGzyJ6YKn3nF6WpAp/dBj3OA8fMZU47TguOtMj/ft0Mzrm
+JKQsxIGvXYE00SRY08UR1LgSvB0dhb/iYCbM3vXe0HH5fVYmk6UydCwQ3hbUTb6
33/WNm9UDMemCnL0S/NbMLdmEKhj55kKdBoBCsDctQO206uUEgueM70XmTH95Mza
SeMV+8/2Sv9GWFvhkow0uYuLgxCOcFn2CzqPNF5KknJxdlK7K7WO3gNd170FNLzz
APPne4jBLgTGj0TRiLtxH6GhNDEki6lKM2h6ruhqwOPegcIsxbZU6EMiiA+2PYAp
Odyo0EGl54MgkLRGnueGxWe6jUrupvvRjvD64sd1SYQCjDrzZEAFQKWmEUxLVVtt
uYuQ9/xfWoWY76lAV18tG5tqTh0qOEoxL2mJUAi7Z/OqHlXruEXeLP7SLUcSRSMj
hW3FJcSuhWf99lAXPKHenE+v0toBIXSzNEdEWC2aL1Al11dD26QIHWQgvpH/v7XB
DSOwAAPmKzOq/b9Nanm75L3sUxns1omTix5Xcs/QFrAFUwksXyjd1eP23IRNZCGS
neC1uoKzw7xcP6gFQiCb+5ijHu9t6HyYxr1If74CTSClyiwCxWcewJfR1bU0q2WW
uSMGAJBugHaHnHPZS7Q9YXU+Zdg9+k/2jybJ7/jgm5x3FtmzEKnWWIzvyjbc5ca/
zckgbJRssIxOKwiaBvBaf99eLKPBF0Cu/mPrQzmxq6jglVHnZRQvL4pgSh4ez44w
yM9zL6nHnkzqBJDyVeWS3kYW5jG6Fabi4VAqeqldiVeaIZKTUqsWFwnkiicSqIN3
DQqQ5h1fktDQi6Xt62ChZl8gX33Vc6dshEXXY8atphYWeoexxH1q19Q9/KMOxfTh
EbqQh6qlL+buLvHcayNZZd27d3h2Wnx5PeodKt+P6MrhiUGw/Xxu/xdqn9Bk3VRk
B/t66a2NH6QmNbFkpmA6tlw2g571YO6L1S9ue/Czx1fM+O6sM2FoQ9aGimHv2b9f
x+pmTc/azO/Pcun1tPk7YDJh80zb8z4q9m6iME9z1qq2T89VDd9Zm8B9jd7AERCj
wu9uJIP6jOuc5Kqv9e7EIEBRcwCMNR7OFqdlvK8OqC/6NdMHKMVxJ0s2DPBB32PG
/sveNY4Nch2dkUZpfo7FIon6GyQAJ527dNT9Y+ZfUsTbzjQWVBLJkalMghww4b3G
SZQX8D4lBquWDPRSP54QLAvETmNp02tpldpJEKYKwaQqj6OW6Z16qmkWhcwHEbV1
BSF5RdZ9oX4Zs7vYlwkjo4fsrLJf0tS1hag6nStM4rmPTpS5v/pFPiDi9IczFzCU
lDj97695a0KKZ5JCsKVfW2VFymJDMSUCDRgZy30dYVtsVxQoj6Wp+eJeCVr/8LgB
ITtqe7WwaZ0ZpnM1C2TMPzrLbFv7chBAD/eLskhP92rngSRWWAhngaCluZ+58YkC
TZlRp9Ro/AZjI0J9XWbPtYBKhXTZvB2Np8x0nJNsAjJaHK/OgS0Bx0oYh/c6HQ1T
U/PzsO3WsW2Ub6Fldh/hf5AOU0Gf/c5V55aWBrDDOa2G3t/4lSuvn4F/ZNyoLPzd
NAgwfy1Obwrm1swE5200j3zXEtQdQfd4Xnr8sL7eU4XoXwbSe+KmeD2FOhhdLwGn
UqHZ8gXJXyDvtx1T+r7x4tf/pjmYmxIvebrQUFMc5WjHy/tbtqYPuFERrbB0brcP
5x3cW8uIcsv64yPp9sTxrPBVoLLxYdQeskxqIWan+niKfVOTpu+/0/8jM7+NzwdW
uWGoOeLz2AVIKOB6HW0vj4QyJJ09rm7I+55Tu1MSApcf/f04jF0yUqcAj5KC+5NU
Wwih+WazeOExMH23pu7EfAV2j+9gzFW5CDlnNGVDUiFjaxv0/4KgaFPIXdkmo+Ww
q7uxJOD7slXASWnGNxkdeDcEfwlRuT4U3KiUixjny6QMNRgxZMvnYpAHkt78G/Np
08YkdSogLqKcsbefu8isdGcuGIFTWs38Uv+ykGmk6vznmdpGzF1F4Q7pEbOG7lWo
Nk9iNn6wsIHPB8N5j5s/CguKSfO4eZFAHwmc4QsjYIexqj7+3XIB96+c+rTYI2uz
xcy38C6KyNdP7okNgYKCkf+UJq7R+ODipshY0CfdUqcnTg9ut+x8KBnd9YkkdEiS
RNskAjdiG0uybM6KfI4Y1Ht9wmmT8zeb9I5hNMm32YZA0Rm/c4qXpFmk8s3p7WRj
8NKvi4ys/jADzMa7DtinOoBTPqYvsWyeHjA7eH+Y4iIrkdgMpSBVRNC976YITqTb
NusA1CIHA3/UF+oIIileREDJPSiNQEf+i9qYnVkjI77ZGpsU4qb79AZDMZCmDCsB
uQNKSQLIKGChXnd3Zx33knW3zB8fH5FjzDZE1z7NwZtRtdalhXEq4GosJHFp6jJm
RpyZ8YxCGEIXBa2azOfw2YA/0A8PfrbAHFjpD5WmWqJzidOeailqsbHDVY0c3PXv
02gut4LIZwZW2VxqeVOdfxEoPQAouoTfjZXmMmKvIR71dSPwWlt95K0Nn+k4hI4Y
VvCnsXjRxoLoL0FIanvHKSVj/UC7186hqj84V0D5+quzeUD4S0iIx/seztc9fHYl
44QO4hE+K+mzBrTTFrvLevvIQbGuU/cVRkrEgRMONye8VEGhVNEHT24IC7fL1OZq
Z2L6c2BnxtHSs3N3sB8L/HzaHQ3CSX028mIMbVBHrZWzACTp7dp2baaQEswmgrP/
2Uv0xSE4QSAGa3KdFgxMFGYyZtXNQMAApqibG7hkk1FDFaUPINlNqFK9u2om62wF
P1825mkHqlWZTFj3HJDvUQ/zB0Ix8I2D+wCLjJiWQe2dpdfsbe87oc6EmMMOMwwd
56c8o95VjdRA2FnfGI3aK5keNeiZS+jL2+4QmcJ87PhqconlXn8RJq9HemYnkDWE
fwIK2rJmFTSmfiE04qoJuUvHJkofrMwvVzLMEDyvj/VWoZ3IRCDg+RN7utgI3e9y
+tzICcldoPdCf4eJMdjUBwmRdAUGm0obBVtaU5eOJTdCyiam3mVL1biwSJPMpTEq
OUyjoAeLzS5Q9DygYkYHb8MBvCMq1WBplqi9qW1ZO/GDGFcO84eMdyPehToIIGZN
c2o5piwZOj7H+/kOz800dWBA0S6XdRChjxciOwHjJS/h1U0XgJ66CQWnxyBMLqg6
rOSOqHC8wuhpAyaQd9rY6gH7nK9JNnndytCtM6yXSYy0415O4JVcjmXTJaktYE0G
j1Es9EY7/IZmvXu2WP9s88/mWvHbGVFHoYVfWsTzfroZHEweYRurCtRguD0Ve3Sw
SCF88VLP8z1pRfBNk1Itq0KSQ5oWoL7VEs9XAdLTuHjfQpeN3A4O41aZaslPtBT5
hp0Ky6MlkSlnLk1qUaERN61DglJle1KOJKghjBAT2c2PbvaL3aGwB2DUttPMLbOk
NcTZSXnE5S8rhh8oUrDdGPzD3CrRhCE4sC9kdrfSJHUEKvBSfQggfkdSc9l+IKmu
r8DhQMN1Y7WYHbnvIT8RsmN7FU8UQFhYN0UgGdLIDwewp9h+0dFORicVtwySldqg
tt27Nd8JyxEhwWPtfSrr575pnoVkkbWc825vaR2evXYhGzvH5v4l8Qai/CrfBPmx
eWbrJXsbOTUjUMHIm5Fae/vxOsIdmbyFso0CoHfVoPHjNGCPHakXappcms94VhVT
DFV7v44ICbxBf4+5GA7cLv1mljagcTtIwPs/XuQqnDBygFil8Jz3/fm1IERvDadK
yqddjbKBduyPC8MXMjyV8jxmwvKzG5LUtz8jcedFKcAXEMdnE7QpfkdC5yMPKQEB
f8ThajVg/2dq03tqxun3j0M7wwhUuHHFQYuEOksUXCGZSSOUqiz8XNnYqJw/h08/
yawxLr8oTAXW58I45D0u8umteJA9JHYuoLzGJrawuOsudMACseEyPAPM641pYeIS
FUWauy6NjD/YWc0zgLMfXpH0EAhUVNVN36apPSt5LhTRYPbZPS/D9UvycIkBM4i1
CKmERrxOQ+TzJlZU8b/qM330paUjnU+GZRtc95RoC7Z+gz/j/zEPxYpK1i5Ln1TS
dRtRncwHc1tvq8P657kjOV7k/YizR5dAywRQJYmVM0URiGyKCbUZNlZ9ue8NRjdp
R3dD/v8n0F+hDtsuoqCjA3fvHurBvJ07F7qwEXdICKA1XAedKKBAj/L5dL0y9oe6
EQle0YcUncR01xSVTsL/WTwi2XFDwwBLYSIsD9xBISdIeFvFBAS/BpsSyxuqsD8Q
nw7j/9H37VQyB6ZkGnenX/N/sEoqU68xAHHebGIcvLszu2adnO4QZOGz9nt7+qr+
alsdBZFX3U9gpTgQMFPF2kIgSjS8W02Mzg/DZF4e3smE10+97oSvC6reQA6toElQ
O6MyEe0h09g9g+IXRtXgohA8FjFpJQo3fz3SCEEQG5YqyXAnIkoNrmCVgLjFUh8X
3LNm4hf93Cz5qQ2FomuZoCuhZhjNTDogRarhJ5yQ4xtSUN/YBzFqO7SoIIkHWzV6
9gYF5nkpJ+il6zZdkOSLPgnk+l7a5si0JmnSaelxbtQc92BrE97944GQ/3uxhWiv
Bs8aCAP03ZZsfe88cMrxl1xmElmUwQ7GSEjQ4XgrqzkpesJ6IV3eLz2vrf/q8vb1
ajiV5wsx9NyYhyTTspUGexyvstRF9we8saQ5o9Qo/rE8wMBtnEfVc0oOlTutW8Fn
D2FzuIxadG8rYQqqTg9MXbdKpiCiIXwVq8WdZ7t4p6hySUtYng4e5AgfLFF/lqM+
TKsFoVgILxfgc9hz5wx2OKgdl7jPHO1hUXfjfJAwCFlkLTEBlC04dUgFxzGma/1M
RF4feEUR6phTlFuAdZVU+g0kDE8Y5kbaFRuGoE+7X3KX8qTub2iaKUWfPQz+dyBm
GeK7DzIEdlKzA/PnLZZeed9/VX7w71Q3S1DtaJ+3eP0Wo+kWvH09nAyDZY/aOogQ
j9tTN7EmBYk4J1OFoQePHxZUKXUA/15LLuS1wMR3QyK+55kzEg8nhqW8DbFlQ8tQ
TdV8P6n5ULdNtm+pVQAjGBOKrNujdpn6T3FpsyytGeqBsYAFL7m9PxVGDE/NkWtq
A8+KU6Q7N8E+ozACwLrruKDZhq81dxLwp+2gYtB4MA79mAfdvIJ15Cun1pPD+8R5
NSNki4+lgJIw/eXe8YzDIoOJXVPkT8Lp6XSZPiRhZhx9x0nOx2iImY5Giu8gPlez
wO7zgmW7twWhgLznsklqyPfm14fvOdy3sZ90q2oiizGB7egmH41i7qO2FeydI6Lb
4F7ku+S9BsZ1IfdOz/koWu0wJFHXm3J5Q177sRoeMJw9LtbTZkAYhK3y304SwfD5
dznRDdQG9WxIBKB64nmcwheMliZcLj9IMiUZWgKV2fWDvh3smKmxCA78L/Uye/ED
4YEg4f5rsW8TOrkyXNWIQhD7TckkNvTFXr89ak9yZvB43itO8lJYMsUErWWE/3pf
GzSTEqK5sQON4Z/1TVXg38MyChnFNKW4PWaPvYcWqX0PiHMjgJdhQ91cAflojtWA
TOBkNsG2QijqwEpozAMubAWXGyvT9SbRmPAwytI4bgo5Pr+f1mAz8ZjYyL3A0EXc
HwHgpqv4bftAwM77ZILy4lOinO4/ohDSKUrsqzRLYo+cdCKQLsd5JTW+YiFP91Mm
fV97EJUV4+3Ui7k3HCU56JQ+wCU94+NNEKy/fBR26kVKFfUzj1C0sakN5dvU1k3M
lAk9juGhNv2tUWWRdnxSEO9p9yAjph9NDSfLs6LTaWMAnsyoJvaGgzVSDlRBCPBW
eJYakQOHFlHtnU55HLWVF8SqLlCU/0VGA1PwH3FiwV3Bv2Y1FjVSZc0yWeKpCPIP
h2xj7UuYT33ljQlrP+BJyn6thWL42WtTprnHuoPpRGzRUVNDRphmzTfzCTGDCt/b
zgf0Sx6hcCxu5+G4I9QQjetbgMOBfOAJtqIiGeb1A90WYuI4NxJqskxx54PBE8FL
BgvI1WF6RJeZ5/4Ktj/hGStRyjnIBKaE6HHaDAn8UfkY22fK/7JyyyNGiX65qknP
rbh/GwrJiN+eu6pcMa1G21N0CoFnjx6VIoxnrTTbBDuQTVqotHfzdJ+zv4brEmqI
OZjTqGE8Kkiimo55l3AMHnyhRwWJP83/pa5e78D1EEZ+Qd/vxmFFM1ef0mFx8Y34
3c2NLXDRPVGJP+zXxGt3LiTeU/b9lkdqw0GBQdLvlB7ogkkgJU/xir77FGcUhvV2
wfGqKBmlNMdfu0bT20ezxGD9zrRPwmRkrfQN7r8Ml/3mJ4VsjsOTbh1PRfuNsIzc
IYApg38SBdVtPNh3QnItw6uX3FtZa8XMzNEljigMDiumoBKn4hqH0drZIAC04Oii
ODCRWcQgqgoe6x8NUyNktX4Vh+ChAAy/1/VwO1vSPjBTIs70pwiYXDP6nRquyFzG
hcCmtOBNfcT3iqnr+dDlQwGbdEZ7uFs++izmPbArgjm02mLIQ/pXSbZLRfcSOf7d
brbqjU7z1jFuyC27YXm5h7LMA96kRaCVndZKvqzLeKNcqt5y/R4YcXh/Az4MY6nZ
eYnV7JUhujerf7r8YW7Dt1he92tis4ndTzmuXgzAGswz+0RKR5B3oBZJu+FKdlic
JrGuDXPVCZUZx0EV94Q6GPdQXrnZD54K5SvwCoosKb+nqeZ0wCJ+5uPXN9KXYdzO
ARudyf6/d1awtbgFDYcq3Od34Rv98xfsc9GHMuKVuzpkLPgJZpu/CXcsH2UuCxAD
34YddcyReun7G99c8nGStR+mpcXxt208iPiNfARddStDwd+3tGWxpqfD7huUpMTp
3w+UxZc2AVxoqFD2D3hOG2cNQMNCyBNJA0seYoVZqDZBvbuxBW71d8J91Zz2BHJ0
ATGz1jGfDUAZtZI+y38TvC9ntQemgIMJesnrkOPigSnizBQv6Gf5lR4w7XGhRwQy
kxIGgXIgzpXy7L//Vzv1defd33Ss5mi218/mi+GJ59lJ9k4Lg+PcbeDGGe7ChQki
fanApd8ylp48OuD8DsE+j4PhySd3KGp8LV8upBVFhaxs/d+Pv/KQhC/lf+/Mtxvz
G5xuK5chXvGaFsWQS7w61DHG11gUtUtdyYbGu2ClFkHcjtg3GGtJj/Jcd4HMQgaa
55BnlFRFTo1sRfqgLTHWFRnZX6TMGKlIYIvrITfYBvIis/AIlo36iYc464RAcXN4
ESL+0hz7Hz7cyw/Rbw8QzcQAuJXM6gtC9HoHjjxgNI4Sh509oUfKiplAk7FaPNPj
jfBysCHgVEZ9sLb0Ku8CieeQyADL9m1ypY50HMWa4hA/WFs6+aPoPqJBuacvB3dt
hD5Dazj2HSwXzkIJJHelYJ7++cy8SQCTMeY/DtBWYyRz8qkfr159JWo96XUhkyCp
2zbIt7CTGc5dMMkI4Dj+fu0sGwKZGr71Cix5ET9sT/EtP1AnOMjJV1l/087LqbfE
xnxewCi+UNGz/sd9cKnFgUF6aI7Nk7tbAsg93X6Zt6595Zss6Z6ooC2Zli6ZPWr3
sSiXuovkk1K8hVU8J/KOMTgvrCB8+oScq/7OzIRqGGMAlOdmgCQ7XheQ8DwtaOxg
Hptra8J9GQh4f0RNqljM2yEeuVGMSnaI6RhRIQwqMIaiN5bXvkxDRB1kVj4Safch
tOc3260jA5Lj+iUOqm5a4F3DXTd2W+ivs5fEnipmAa7NBcEJo4b41ojUWhrsTbk1
EC35MBEiI+e0wQemuL6LG9CbEIOUgHTU+XxKa/j19HhRLcCGXDHYW/vKBqzCJScm
HnSt1aBqCOeVct9m8dttLqRkv4D1snD0teurONqj3gjw2SA0pC4o6u5gE7uSr8ng
0E0ETlwUKFrrpasfYVptHYyRWGBAl9XuED4nNCaIZe9nb9rJlwV5EcNdfYGm4RWv
ZuonutVIkXDsmdWfPR2vWa3sLcRoCESWKr50Gnb9OdX6WybO+Vjz0g/V4sQEQn/Y
UwVfieH422DEbfJy4DQAh4MlA2wUBz88lOsUP2WdHeZOhWkP1/l8BrtAfMDhRwlz
kAHU/inMC0cmT1Qaz6YvtXabUQh0BxOssWfMmtpuse1LBLPJBd/FXnN9M0yYFfcC
fLCOXypMFGn7+Ef1tbopZ7RWDo/5y54UWeCx+KbNZwykozl0UyWVyhItY1X22PyZ
SIN9TD83X5BgORU2P+U7u6lUeBdJRBjzGNRCMPNTSPtYpZlUgB/71ivNzVveeDHO
1SVY1SDyYXbJnFqu7q14pnLQOs3pas68d/CYhuDeJ7+PNpg93xF7QQb8+b208n7G
iykaM8Q3z6ipa622/RU3l+ZSe1kt4K+9K2QBKMdWih6+qdZ0bzuu5S33MAXGpTy+
E2de/fve76tFFbXN4yw79hbrKuMUubE4f3qVZl7nzFwLNC75PDOnRR0bbl1eaS5b
HJqOM3OJuRIlIemRQYHh/9HCDmVGd0VDvqQ1DtIv3zmQcFPQOGvL4p0tUotZKIN4
sAIp6JjsuJ87rofQiw0LrUD7DWLR+sbKQQXZ97kotvz+06kKSrYGMIGje8RHBAjA
/LrqLtveXzQtN9oXETu7uCaPstuHhMUHluGb2cpfAFyCdAwh7oFxtyZqt0OaYK8i
km0hiOOWrytNcrrshm+7YOSiRedgnDZsOmlloR2s0Zht5rMiHuPFHKHxOpU0B1QW
5LXjpdE/sXL8Z3boGGlFVOcTcW/hc3uW92OZXvWyc7vk/e63I7FPNB1KJSEQ9Q5C
MSLfGmdyw7caQaXOZyCrHb7+2MrY/hZ4VL3H1Ld2Xqhnx2hmIbxukRhgcfgMUdnJ
Yx7vVMB/JyUrcSzsquZknzCESzbTBy9jILV1fooq1BPC772xhoP5pv6l/gl/WPWY
nmGv/cOuBl0cbU2ql6NtydCdaIMkzX/K5nBBUOwDeJWJOI4F0IHgLHGcutRnjxkZ
/XnOhyqe0DLcFsplYKYNUsMEmJaINVC/KZMkS1Ww/M+rlP0eo31M0JPdO7piYa9y
AtOGmBY9jENo/GgS+K6/lO9Yxa0aO17zk6RA8vAGXDuTcKe52SZ+ULESXFBx8BNi
jidGQIxMKiSJeIjtDjFzfcRJB/CoDoSxyD0d9U2fD/IyfyOHtKsKA3uchIMn5U+L
VCzau9TB90KHAokMMRb8HmdnApn8PGbRqH65BPHpgUgzXgLriAcsW7YCALB+Pm2o
Y6IXWTOdke1GMX3iPUL928MF+59NNwQ3VgdSVeEBWsPaIBPCOBQOvIhWj/+BvOxw
dEX4lobhQIHoiQ3Fj5e8NzNDsOdT/cjWIaAHV9wnHWHSguW+n7wD9Il+I6NMqODK
OYPYIlgfR75LVaCTGS2xJdfRrWqlHFCMNp730Xh220k61Nvnm3k2kN8Rr4Y5QEGs
bnDB9mLm/Jr8kqGPsuIZmnD62CGjxjrteAqmp3qQXzd2mzxxxUnb/v1MPZBIhS31
a8Zj8Nr9DWLf9iMOhAr0SqtsZ8EFUlWXJDzn9kGVwS7ZmF9QnmNcDlcPvXQj7XrC
d8FqYLPdoAB6q7ySMrE2KMYwhcCynAf5Ln9isQ9tRwRzKlJxhv5wMz2qLT2aPtFd
do8OlZM0K6+XJ9fhrWpX6uEv9CN9pr8GJlhOhVyo/SyMGxPvO58bCyq/GcEZwH/H
9j3N+3So+4hMQ1ld6viGp9Qokzl689w2dvR9ir+uZ7D0yhGJ0Pfa0h1L9pCRr/Xs
nPDdCJKmm19U6WBRyr4sdxoH82hNDhKRVcw16Um3lQ//CBMLMKmzVBOkxU4uCxEu
y3ET5mYHVn2XPAT+yS0Y9wtBZpvt15wJ0I1ilrV2Cr/K63FBAbvpAWNsaOAPojQN
JGAecoId8w80VL0QgYLVejD7T0FmGbC3df0X3UvYSd96eBWLhgg1t84bTOHyFd1M
DxrGlepOWtxW5GYn2qfZN8u2nvTObpdnt1T4rOLoiIT9uSvGbvsgjWBzhFQBk2Y8
GcAiDyGTuJPvpLN69D24ILsmJhnJt4n766I/33oHC82MIs/dj6yl0VZ+4cqlOeGi
MchNAp/g0TEscjTHQUoXMSwq/2O6BBuN0Du0l3OD4tlZ3E4eeTCLjVm08Hr3hJzA
mQmDeNi1Uu8VnTQDkpQ2E3ID5wEvLaqhICj6B3T9Vufd+mxbCeApglb0NJfn5K0N
R0Nn2Fykct8xyJxwGJxBj0ZchDizCU3aut4xwSnbLl3P3W1/lLBlbhJpDX9AyQS4
iwl4iP276UjaLYQuf1bEy/m3h5TNL69u5lf959++2lnSFKnRYppJQqZsvQseMnEs
plSDPEPxesN9bsfCS9iXFVC7DV9yONeZa3lDToK1KRN5TkwW9V7iiB/NKNiOlJRu
sr5izo+AXg3XmSsPsFIoxSahesqKjpyJa3InmmA786fnkNEiPoAVtuf4PBTgdGSP
JzU4pHSv0UHE858Z3rEKbNKeMBa5yVmT5jsBNtaKMVY5C6krA+dThZVtKoEIXOQE
8VQfseh6LM3WLrIyXlALSa6BQHEhwcJPb3CFPFRIk0o9FvT6cKue7cGGHH0PFh7o
iRafU00ata1+Saub7fTslK43L0gykrdOKjV1pVOjOtJ7Wctk1mr+mpVuLgpKDCQ0
PckztTRHZ2SuIaahoT7z7DktANW9s3dLTlWU4KS3DZsI2eA1TCDe/4CgFITVdqBw
ik50q6QapkrgnLDQhpfaHIVZWahwDpg5qaf4OJsgC8yz1tvEp8ajE1FXSmxgpTgM
BtRDzBvt43BRcr4i8PUcxpdjGfuedOmqnoF1bolAi/orMTJl83bmzBbCs+RLptql
EkUztHHDzRqcufKKc+4Mkmsvxp75sLB1qE2Eyb7SO1lwW0zKGAXQ2++3ecbEDY0Q
pudoPrN8hX0hnSaNVTL8XwWPsSrnIy6CUf4vaN58PUgxUf3nZikY9hFBqFAJ3MKW
9Ai+o9f7fsN+xPKDj/trIFm8zB/YkKh/LuoZjz28Lakir6kYdppGpUGFCwlXkWbC
cmTboME4P2A3I+GZHlC5vJgIpCjC9nw9LZ53WuTfXeVFfJhnPi1Ll2ns3hQ8AKvH
6t9sdyGJhfcKbX6kP3UsQ6/WZzeM2bOq0kcd3Bl6LJwlcOmgoq3XgJAg2JHpNQf+
ysdhB2J+wNJuctEBp0qJ1aXuYzwbNBjIwMmG4aRGSaZJjCNihq7wL2v8PRUAPxvY
GnlmHrjapSvl0fVgvgswdu9refsTgi5wnbgIiEIG42vx20yxQd589KhQnxEtKLt4
8+Gb1xIT3VP6h2zWdjNaFAvlXQJzCL2I8XA7WUNFu/DynN3LiuwZze8L8zRPKOW4
RzmreYey0VJggNpCRRmr8bX07l/RHwrm8xjHdmrfxkYSw/8T5VugXX/UscXrjnOZ
OPmXaiImy/fRU/Jz0mlNpTSKOhiDJdMPrzRU0UWmhV24Bw4nKEdRG5PgmROKycW5
zt8k9pO2ANmei4IR9aHtWnKhgkcgeiGTCEeT1jYLam2MEpt9svhzDdyEapHYevFk
gn1vtWA5ZOSXEhGPp694nxa9k1maermZK5A+t7v0rQWX8g2O4r85YEaud85odoaU
XdPM9x2eVPOczd9bkCl0YUcUXNjDVHE4B59uK3Ndn+GfifRfwMtUCcnqCJRepUtx
/ytgT8qX8P9jgKADgck2StY50bQWE9Y9awAPJpsfKW/RZU2YabnQCb44DlyopFTF
WlTOrlRkyEbna3bIWW3ZWaU6wuqtTvyXrVRFfk5SBYDKb58HNiDUdZDf7fOnJsvK
rqQ9Oaxa672fqtaXOAr/RUUV/uhQochLvFSk3EHrCbyDhnPBFaDODIX1FlktFdsl
abwLsTgO/JM4oAjooy8zvtdAzSpvyQ9ViLYLvyz2UpxeldX3bcXfenvMJvtL1S9u
xI+OJnLbbq0oodGMZcqcJmOdPwjw7DYzfoLfgeVpZjls8au1Gk4ZNoWPV3CqAL/e
OXkVi9ra19aMvx1q57g9E6W/19PS5aib+FBbegbS8gn+eQbV6v+ETHaoY6lueOsH
PwMjqU4eFtJcPlGoNzr/GpVLo3cyOcx60vP5/Cq0UNDju7lM4iUl9KuSFJjFNkAK
SgajzPaTYoCqVXd1ulfejkVjoi1nzoCle/iWO+r7Xawq4FsJCoQ+rADkFXHRbGM2
yMamAtmRKc7CFrrLYP4M0V2bgeajTGejwfDrzGa6yDcDsFihHR03A8T2t8LDGxyQ
U/FiLIb+JCfmddqqq8D21eo7FgkwD+vpCeWaTCgB23kV7AED6/5PrCYxxrHrnMAr
106D1RAJX36QfQD5XnRSjVjKnckHRzxGGlPV1VKIGat4Rw9zQVuqn06khk3Y3czF
+MlX2paCl+nlM6SLhQuDsHQ3rrebWbiya3oh9UExOegldDEeLOSgGRPjlLsQiY7M
0Sn9UGECVmS1t8XdEggxeDldnYWUu2APWeiErYFZzk6e9uYJeyWxSBwd622gYscm
ohS0/Ys7DGD0GoesSdQYjLCv7dYY34DlXYku1VYOHO7nHGNObaqzVJnUhOE+ToVw
k4mGm0R1smCqtIlhNpDuuLfFFup+ag4Nm0g/F3x2+aUYWiEunmupo5hgqcH4/xkI
moVLZcoFuJhJhXxdNguV9CXEUZfF9AyBL1h0tPuL8+gpVMr3ppiDBrg8syl0mZxG
P80jAcKpbepFNeyHgbeRzmbIx+p7EmvzFGGfJnV0/90iM6tXgPwDyKX6RWjSeenW
rZ4ow2u//uUftd7GVCfe4lZV8vQtH+jpB+EsAGLvw5IBxpbKRp5H5Q/INBvIXxvI
IsYo0LAyzNF5hcBn1t/Qf6lWKPyqGXrJmUOOuRNKRf4fLI5y3o47e+uSTiEwNTe6
jrcDiKkQ1vQWGHo6jw9+l4AIGPh92aZW0tfr4cL2EXgDjo1tCemQwobsLrvvYNlI
7BF+z8SRADoW5KgTmIQEbO1wHphzp2nkXlt0TjyCFz8pASSIYofMhnqJ7rijZ9o3
hLlMK7wTITCVPFLWSLfTcEfa1E6Gh2T1oJ68cPB0SP69pcUsJGqVSt4wl2D92lS2
iW6u4KdGpDPEc4tGa0PSYZYOPkaJhrFr3Ve2FWsEaXw6Nvj+ptrjZdqEWS2Mgf1U
SN7KGpqpLDqSEdwqH+4uy7mi+xEDYvKr1k/Bpg1N2JLm5Jp6HFUB01ALHpyJCobd
lHXfwmva/6PyCKCsqWGCi63vwJmNqfBhpP4t7cQvCunO+guv2ltUYyoQ/teyo/KE
BrriXNHfY9pTEKXLMHwmDcU/SOmiaj7kbF7OZ2c11GTMLq21BUvuky5bEdYjw/95
1m3FBKs5rPVUgSuRc6sCWt+4nWLXFHpsQ7jPFrd79EBN3SsMCtGEgDcPJAggrkXR
m2yo1FtjntpyxOV81RlLeYDO/nyUjfk6xzLvmYbAsTUq5YO1nMbui1aPnUXTfkus
GKibD/i8OqBpfEbsWI6HQoOWTv/dpVoERXyDFyCIYdQepHMdoccVO5Hs7F6V05rV
O494UewyxO0UAMDQ5qm5PBXWq+LfTbwrR+MXSzvIRSY4yHMn5J2rLOMh2UXbwje8
s46iBFfXUzoO2chZbnjik8QA9muDJVcB3AfT7lNMWhhn1pqIRfqs2orQ8+ke4o5G
qvNhFaB1NBmMN5Gy8TqWGrsYoufaoLsTAmGitXe5RnFbSPImjQjBIZLKTmtOh56c
oaTHFrHFpvGuyB7ok6EU60Tm4rM5uuxpRoTFbmNCIW86AK7o7HrS+Ta9sN52mHF/
p5pHQOgSmenBzmfttP8Gt3/LR9tO8b6yIkZZYRFI1IvreHfm9oHAzWrElSFvTcMl
oVCuVOEhTYsWN/6BmMxpL3dSAxl+LVQ4XrGwD9jcx9jFk/9l6awghEicuDhj+RI8
orG3vAx3egwBlU0byYrFhrAEkWiolOTSJ7P0LF68hpujcZLNpYZYD9m0VjaFqY79
7l5IAlb3qdEnJdqMR3fksUrcqK5/qPhuGILGjHFS0TY663uZNWDJmgmT9oUiTDxu
5fzxSMB6MI5sOWDR4gRS7RWRSwU0z2L7QIiW6e2p3biAyb9nht4GsAxs18BUbHSU
/cA8grilHXiak2w4KZlfVjaEz8UxceVFoXT66ZJ6fh9+6Xy/XTsxhoUws+s5H/r5
6n0+u3Q1OJBR7HezQ1EKsj1VRxnO+gfcU3y812ZB1fXoZtE3auiKANPvSdqbozIj
brxMaT8bJWDoM6gjuicm7FCvZwYjUUKe/2e5eqkx1jXkqTsvWHnb4UsuZdxgN+Wq
oTRb/HSD2vIJnedaglQ6OB6O2tRJCh04T9RF+OFm0sUnvpp907fCDZr7Il2Yy9n5
sbJJz4IUVSiHmossc/bZ/PUaSHXDwu+XlFLwf1duum7Sjw+mAlAlejU5nFgjvW7F
4DR8goIPeY4OgRKehxyApj2GK/wJ7QoWYSWvjEMbvXq1jQ16GNYLIDCMq+648aZT
JLPa95uwOLn+1jHucRYyf2gWUWsazDrzebAgejicVZokgJKE75F5aqUWH0UOKlCL
KvMrkcXL6dD/nyykJRVFX29+RbTEn1z0rGaCXCHPYs1UpVCYpUNC3ldqoTBWkgqy
SCIXbmw2WuDANcGXQVkaymi4LDb/9k9o/7VN9tYc9kctDTjnLCsSW4Zbyh1/EIIg
i+woeecnamGL0JhqYdJR95aZaG97ZKhpl6cFnP/sjoacosC4H0z4GZSiqXbGqyty
dfzP7pU9LwJA9m6VaMQ0Oy0H2QyBZdNUSR4iSBgDHe9Lh44TPB3+2dBmoHh+dkRe
fIAlG//4T2Lnprvz5JR4tFFrFurI7YOiCZuu7Exv7yBm2uKs78yfAJpW6xEyUAvs
LXxOzVgiwMntiki4uyMeNWIoCOMd36OwaiEDkqKFMq6S4JEm9XjIz14hj8Ri83x8
HUr0uLdtbl3ojteC/DXhCNKivrjbgOTTX3oPmaokvZMmmVV6M8Ch5zNoRqebBGnW
Ej8m4jMDshPkejisnuASTST5AkEhqW95W3OW2ltzKqH1edASkEOdQUVXKveL9iEa
tjphaD1NLDQYqqVFx6ehLGbjeQovk64gJWI7mCQI0aLEp3DwWl9sFcU3w5q3Qwh4
0jDcKKyG9zQw1IWpIWGVlVwzznM8oDLmP6vikAu1MzWHD5kUCUVTgu100Wm/F+fc
Zw03b4ALI9z4idQ+3i7VdtmGa1p7tMGZYZ57/aHH9S/uhumBe6ZcgWDQ9wTggqPq
km5y4CSssBJArnrO0dOfZDxw1mKCALLhCTRGmP21gMwiCNTp9Fbi9QKmFvncVoHG
j+mZhmxFgcteuY6Fom78LPfV4zrvtOcqNF9lZCPvxtwSTIJGKQy3djOokw9oLRJZ
gTdaS0FCvNaxzog1cZOankwCqlmtSgO0aO/XXpsDsbfVZPSm3TO+hsgD8dwUcdp4
QBuEsQCPE3u1cbP4Vc9b/NB14IiloXAtwtM/dOnwjqCEkmIZakY4mz2b1TX+sDki
4TlWFJTb94MCdSPCGH608bep42zeZzyjYLDWWM+vL8PvDQR/PB9Rb3tX0q/XLxEt
uud1lMMumFEGdAgqQIVnZ2rRRmfYAFiQnxWUL95514LYccVPvSzFx15fGL+NySrM
O3qLK03jLCoUQJay9rJKPjtly0bfDDuiyU5iCoG3JqvWFupow2MaHwHMXJSAVZIx
h8TggtPMEMSUMhiCbv4p6KqmY6dlaPtW3OO4YibNGzPU09ssWcEzycxTtf8zRUe5
94Ijg44gj9N7so8LJLIEp8Wh2BLsADAbcGV3mpW4RkrHcwZAxtVyRzLUeCtlynZt
wFyLiVileTKl2rUIqCtsVL4SGdEYbAWFGvn3a5ob8TWvANqg1jcdNguhh+r1hgfc
qe3dn/nLFMql9AEREz5HT8fM9KvVWkob8705oR8GpO77ZxIgdbQjFqniDTpanZFx
ew2WhffyckNA2tox+NeyDev2HpkDEQvsvmJ4T3kbGUImrRof4Ts/gFs8TIkkIa2e
rvxalEn1qzq255GOSHqS7hkUPfiEPimHNab5gRrc5VvYJXoOUZ9cnnHC5mUT8z3m
02BZ87zGQvfKiybF5VI2TbmzQNbIrIW48c65wQi6vzGnoRWI2snM+UJ9ojG8AlAR
G3XzfebIJgOWbpdG5YX7ZATE/aAMy3ssslTSeN7fXYzBWJw0dOXjk0BmrDNLIec0
sq0PA3UJoPBsU9QLe0wQSiyxz4/wrU4eGCQbYe0NGo6yIXco/O9KYW7d8mMvqTYZ
Un1qf86oa+Ysyg0jlNjqkYQ4iLHpuSMQqlWef+OCXEFQDYgofTWdqLTX74KghJpL
HbjCG2+ySJfaPPcJSRQ+lODWVk8pakrCRk0I7Ledu3RnGERZdGrvxKbQia6ImDNB
5UJoAC5vS6qH8hFb/Q5t6wpzWPwYWq0gPNBL9yFgqTxjmNDMZyXLyY7OI6dxjRES
oZDrfiutxt4vhpgupakvgEuvQRPz/ngAgjMOgLb/RWdltHNliWBqDnjVVIMflK3R
k/UA2/Id2EkZM2axziV5JdXV/3zavnhjxxBuSRinIsLvtIKOsXqSuIeOeeJVmui/
uZmwAq++LUkpbb5QZDhKFExEm55NnkQXXzNR9Z/X1TMRH+RHEeptykCdRSVeZiK9
X9z3i6qWzdrxlp8B3L15XyLEPphvp7c/nWY6I1L2GKYU+r8XXcboAJ7ZX/UOowUj
7r+RKaPuP5yfitpQNv478DZqvTQPV8xsZ1rIyJcrXuYwLJ/otsEe0Rrx5qel0d3p
FSSh79LC4fUWA/Y1nhWw5WlsOeRmRTjA1IiqScMbhmzmEy8FVPfyl6uwgoAGsB1y
rGlw3hp8wbPE9ftsX0zaRdirGTlxXZBOd7uayOnb5V+9k4Y783uzVfHN3U9x5Ugj
7iPsw0TU8qXhSrIlOxitRw96XIZwwV1QgKREeHCAJ41dflW/LJtlj5e6mB4K1qHb
QKPJCOCPcNlvWxr05++kfgGMVBSrSCNXFi1ThxZ2ElIlby43tS55c/ywNzO+xNed
kZUf4IKdWB80sYVW8BClqq88rLCC1mEIorMcIyJuTCw1sTiIMiEgbDvo6PkuHMV/
igaXSApMJ6jd1gOZMqXiPubhpeZ1P7FMHruWo9ZFKDX9iGiU3sCu6bRB3/YAbip3
yTg0P13aDHd+5+2wHolKhC4m6dji/nVlpCrL8U0yCO6Advsplht9rMWmkhiCJeub
jukT7+z6mKgtg8UdSMD0JVsHdIyMNa1bj2YTaUrg21toQarnLLXRirqwUfAMZYL+
1SIKS0taAwb4XVRBhMexea+qgqW/uBYUl4sZ8OdRTwQAYqxqRGZWXDlEssX8PInD
cYGwkunLZttJ17ojg1YlQ8PP8HiADITsZKUpgXxR6zvnSpj5SahQKtk445J3YPDE
PQAeBZ03p1yZ55pXbVrOxPKpV1bipnoB9WCByHkp8RG3mEZ0vm1FCU+SKyjv6hsZ
cDfKjukH1YNa2q7KB50WFy1KqLIQtE/vymn9C+I6vLL1k4nrErffKQZxYGAqN9vI
WEzv5g2NRjRgznzoyXve9gwyGZZYkv5+RqPaAz0T7So/bseh65Cqw1jcl/0fBcZY
S9IVdhJK6bh1qpRv0A4/e9NJWRlH0huyPKql9QMc2LYvM9YNJE8+/73QOQZ6mRPw
HoM8zVUtY97JVZhzHXVhyrXuLjB3tqzFdVx2rqxmvKk9j4Fy/jUkfljtqjVvo1k0
sc21A3RBaRpHNPMWD8amvPLQiJhGbjjSPmiLsAoG5rrCajpK/Sz8vtQk2cAftZMl
XfgNFnG/g3ikq7oSz02QCr6mfvPAKUXtJrvhHn9k79Xkhag0gJwjIy6dXW643jQ8
akJV1kIaHpHxDu6uiKmI3xEqm9lhw0DzjlELc0EVheupiw0rL8zDKqakpWPMEhAa
GJghNefBsk9xY77Rea4LuNkM6aigR/RQhC+unAycPhOiXKCOR7AjYT91Epp3ZFgO
yTMQWQXaqc/mgNu7fI2yepcOLmB6TznSciby1MSj24KIULgJvNn+Fx4+TQFoH/Lb
pwcJvTMIf9aGzc1bLhoMUDUP1q27kKmnRLTjNGMXqt7gZuPb98tG9Nhn8f5pAEQV
zQRGedN5j0TeZgfSnvmHRrc+mKyhTBR1sFyYjMOqEvxoiK7vJZss/FjN8OEEseM7
EeatWjuBTLiW24U6VYGzh8Y5n5VdCsKD3PsWl7aTCM0dTUqu/rjMGviOi9iUMym5
NwCGHUmO0ZAiiyL3WmMhPp/whcKkjoUNC2s/kJWXbKNVpNEaBmzzJNdDyGCELS3R
2YHH7VQmeUUcF3ckb8trgKJi7xUmbEIBd7nmgBfnjirc23GcPsq7VZbRWhgFOn2f
bh1mIjUbVmmwcjJ063JWgs5GS85ZpkJYsPOeWMAwosywkLxre8OQyGa7QDsIcqyU
376rvc5driH3R8vrJ8vBsXUeY2buJI4PFwe+cJ5vOmyK0jzUvG6H5GbVBlosMRg0
pCN2qdtD2kcKm/apZfVahIICNJNMCzqpay6G8Kob1iHTAuuwPUPHsL0S+L+CkHJd
Zyf5pAZPNLlBySlVXqDrjLe0oIvnE918txocepCup5kwOwfADtT46xM/Zm0hnP5B
fccHmMMA3jWFjtaNZ9Cvn5hWgIZn2EaHUGzMEGsUPUAQSGdg2FBPMIZ4wxQ5WPGh
ZpEPhEI3PvfNVDIElSieJt8nq8F+DFvsgObxU5D90f7vB2/D0chyNE1G2+cyDov7
e4IZCHtG+EVI4VnE8TeAzhc8o+l5KB4hj5bPFWf4SXxbtU2dme7JVnx3N3aqc/5o
jmCn2G3CVerLVhnWhHcgSgOvldeYkQ1SnDQYdtxFLD+nhxhnuRAtRggtgtoWWwTc
ZelVP0NL1fF/rFKG3rM9lWUETDfLYQgUD1SNyYugf8jEsD/lgfuOGAMu26+LqUE/
g1uBd3hioZlC6uhS9e++/rsP4uduj4MRP0BfY+B8eH0=
`pragma protect end_protected
