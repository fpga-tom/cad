// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XB9wMG2v81r8eCSSMg9+7WlNK5wCP+wpvMoi3HjyOGIAt9FrBm6dnPu2przLCiB8
yUlwYPs7JopwY0oZzpw75l/KSViLAXbxhcfniqXhDhhPYhKaSp7M/eJDqXpaZqo+
jU8gMNJB2wI1X7FXJ0/OfYDNLRPXFZRlHJZYDg/CHmk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32976)
XWbAPOAb925/9259Kjop9c8dAdpLZ5BZQWJ0/AdZeYhuG2OUf5p6G8WYwhrawQfy
s3Ypz9JRQCB42rRgNPIoxIde3+9Ztv/4wAOAT20UrxCGsWZldE2IrWxhZXSGS4jC
RwacICgDOGXU6BgyspvzZI2hAU7/RxYlMhzN16gk6R7JDd8wzsSFrQ9v2FR5LeYc
m3mBo4Yy9Yt53o437HeOpNUwmtBX7FQqclFY8B5Npc4EpjAd9ou07bIQlKugEZvc
+ilJfaDT9AcTD5yRmaCbaiiHWQqVPbIbgLSerOWecGwuaNuU/g0U0tkYUMfnMmFp
/9pd8LJwwygPoxxB/JfJZrlgBu+xd+b2DoWDNLE4h8FOWQp4a1GG7+caCmGaDQ1I
juMsuM7mlcDZqu/K283KKPhMukyYQzgREPICJwaEHDRhRgvOIZkBu7kWcxS6hUFk
d1g7buoZHpung3qE7pzab7VzSX3g40WRyDvKKg/vmRFaIgy3gyRC9RbB7aCRWX2F
+39AhMDj/VdFIsplb343OC5zZVznTp/v6tCpb3QCFyZZFegYc3FHJBF3xwicSmdR
oPBwp25QHPDc/HA4dr9Px1SP3RPkxcNBfYZDxDZfdQmCoN3ooPReGlJOpPeWrECn
QPFc4VcKTCLWdrc712VOMoUN21utpH2uGtiqWyo6i/zrFiczg0IR6uPvpIl0tytw
Hr1R+T3Ohr9a1BU+Ia19Xa9Gth2nj5KAA5cqqBKYEVseweizxbbeh0I+kY0aeAO3
DczaqgR2gEXswZb0l4Zf0xIa2ZQgKhCwwPLFNcyc/mQKKDWnaerEgRndJqaZKYrQ
/Xpzptt2CXNZlj+/A6LW3UdYPdNWiNChBJINDFvg4YuB3DSKTEZeR1AjEizReuCL
q6OxTgZvd+aHNf+CjhiwwBuoqEfCr6EdTScNmarfP92pxKqWFulSBcMwBEzW3EW8
lJ5mraMRxEUFAnFMoFsAF2eNLvesAjqcK5+LlZJpIJZsEWnWziRuYE5PJhmU319R
FHaEOb6HZ23J4y82VYFYEhGUppP8B03mWsQYattyMcaDbQ15AzosFkaYvFzoshKh
2ZW7M54PqpNCTmTbf4H4bvv6H2NWVK1WI0CYO1ybmElkz0jnQ9mqrKLpRg4JeHgd
hcFKq+Ifcx73AVpF6qBCoIxGqlKTlaUCtQHpVQYTueOi5CfmPHJtucZchyMB8q0f
x0ETcvlIZUrqYGAfBOmaz8b0qt/WX0thPneGB8FoaVoDlGhjocN+5YorDyYXESQp
z2lP2DpXyEr2bH6NchrBOj3Ox2alVajh8J7iN/7UxjmpqOunW50c2LTsO+HGbtZk
9esQjpVOYdexM47CYBrhDVnUStA4FLK+If4sCgVfhCzT3odFdouf/LFQGjLZz9VL
ldyUcdiq6AqBbNlHyKrPoPk1IJ+Vurvgzol7UDvLwzdlt7cckDItLBw+ODNn9+vU
FxjW3KZWuXglGfC4477onpmAt7LE+BK9ML5PZDsvp43Srhgu6WzmOl8bPVDJbJ9R
K9h6z3Dccmv8/eoCHPB78IV3OhSnQqFS70v9oWD36Kdtru9P2kJBcQL8za8KIDfE
ZwTQnGcSaNsFAhpervYubbdzbPm2cssIdDQv1UywOCmvFWv5EBkFhtdgK47gciMf
YPmDQsCRyRkZNcZeVV9/5ztCW0mRwOKy3MyteEmDFJD4okvhoBCkfoqfW3CYkPOt
A4cViO8/ZAxPw31qADQ48VsVQoU51Rsoft/4u/hVezYmzzj9aSgU4hv9TStpWO6p
iYaTUEiIxUfIMlMHobLQetehHX30/Uff4QGqmY2Y9FWU0iolOcXEz9PXcJHmDUZB
Nop3smYkSUbDEj1NYrQ7mqh67yEge6Mig//BmzZGm3AGkGv4tkpRkzAOt+9Aq/6T
NJUMC1mnmTB5RydFbGZYnnsHK0+Yc3uPzBK0q++tXLuCU02aJmeSu1MKPCJtU2Bx
DWPlf/EufoEGSeFkMr/in5D4TR4UVnk6SQKEqgNE22Dc+WV7wEkDWwiCFQ9SJqK6
+wITWoSd1kvqTHC23yYSOU7j2SZqqZ1sTwIHwpwqpfxeNC69QbdIShGf93uqad1o
77/oJek0Sh0Q0h5IlJyxNBPPa7kX1kTJN0z9T5x+knVym6x85JmJZWFocRMaY0dn
+UzIidIwUlwFwV4PPxZXcaAp8G37OenfKjLBNZxPsWtoB+Y/dXJrawxvpfFeJsFt
dqDn1Z5C49dDpFSwDEfmkcSv53Vy+nCQHkCCVYAnXWLuG5oynKWscMqOso8V1k7W
8Fwx23NE6Gi35RbEE/nHbWiMd+wKf9wEFA0ivsxVZwDMk9ts187Bm62HlflbiG+k
vhmVmTfeZRfcU9nJj8HPhHDDaeCIhhaQILXGgqw+oiL6X+ayMnNnmriRim9e8mTT
l8RrVb+5R7LeiLbyo39PsydNcKXARVx9J2v9SGpbhwvL+UUqpNXh6mheN9t5yyoi
vx0ti1iF4OTd7JyvN95kO0L0SzXMlMzWa0OTUcry8CWr/xs7bH6PnETDLlRVPXDE
M+sHBtIxnCgPrN833jefLAqUF02rU8ocTr1CGZ7oCmJhQViGJsQunPVGPv+xFyhJ
KCHfm8dr9qmDGqtdwwY3R9LdBFsLo7bTh++tIXvkn/BSGzO04XC68MOxLW2ajaFl
Lt55lRfQNdQhhi1mFzKXhuxxgIfrFSu4eqkiapyZjc22kO8W/dqi9b9wTNtWL+tb
Qxk6IobQzri5/R7tKicpgWEeG36B2a2bwKSH6TYlJHjJJF49iWfgw0u7Z2x4hEH+
U+vuMAJLkH34c2RiSooJmY2oEojzAV64hm7d0baPLs0Drb1C5ERctymUkAuiFi6D
PLM/1s3WSJUBJStumv7M5/KJi/PQHU8V4EsyskIHkeSiqpBOtu2/OzdLFAPHCiqD
xnY4Ya1bX6ak6OL6DKzEbxkruCC97qc1A+6LEkxL8oWunYF3dJ2F/fNCi5W5vf3Z
9jO7LmIOitz2QcksBm+TyLBPd92lMe45ea0BobEgPPNJlmXqM2LmO/6NOprkV3YK
FwV3tq6D3oBzddV0n6kr1syt+ne/ENy9lf9/nl+Bhh17kW7YCuP0bkdBBcCNLYHR
Yy5TuVUDHCWJjTeQ2YkM6AZAXRfxnqXNA+Atryidr0F5FFwHfHgE7Fj/WLkenhYs
hT9MA6pqsar3/UF/lxReNHSvQ+17ZeIKwYK92WNcf7PGYxHg4f+tJYnvS4U0Zgpg
o16vh5KAkWGH0yokU0LgjYcbg/fB+W/huXTnRZ1LyBybkHsLl7Zm5hBUXCQybc2E
v7Yd30x2Vu/pTunESw+bvYUIHXduOINHYyRKbYcUV+ejvpd9jncP6kvhLB/yppPu
7EN2byq0hiJJ1myhdTacrVw67/gafbb04mTUKnjEuorUffnIcJYGhLN1lvNSdBV0
IsEmCX4OZH7ehgTpNLkeSn/lhctlSkp4KNt3tjn+DR4wU7fgmIo3ydmmhDhRnEp/
He/reglYlzoiuyMK53sJJEYOjL/QQp3zMFFNE++/1XYfBHLh1xZjt+shav0NieUF
p+86kKWV3xQvOIBqeyYqTAlkaCEwz41CtC4aCzP4ICUx73Dyu6/jT6qCNNQKMLvS
3P2x/1rSPFL2r3B6busL72zC/8Qhw4Omh6eDOpJofa2hBg0X72i/lqJ/uyuj3UL4
x0CMZZIYU7rP9hwL2Y2Me8lsnnYOSLkbCCgsOnEoQF0ovwYbkCQbIRXgkIH3dRmz
xjVlJipGKjMVYBUN6mVVii0WAecDlvHhIbWNAjTjDniXy1n3FZfjnF8p2Q4YB/8W
zm5XEbUznt6IpWxo3NeQSoU9NJK0tfSjrXQH2SdpPZLQW0iu5kVabQmT6mp9AnJC
X4+KvwqtcE3WPZ8W+zN1DEt0ol2dFTqn4V0RzGysipdPShHIM+I4R8XOFEYGaV9b
pAo8Vr79p2rdlvLz4re4K1DDu11rQXzAKcDuEZKDoPCLjlupLadF2/8BRE2K9b/4
D1YA4+tAUwdudgmicmcKkupj6LmK/BzbddhpEcW9qhMkh+Vz5eWvOh6fyHKVhRs0
6ITpeHSse/zc9z3YAEnH0qXXBpN2N9/6fJiC3/nsxqJ8bdCNS9fv+atRW1aWZIjO
Px4NPZUEBKurs4Fq3VJfZuIjJCPA5OS93h/b44YHpfgbha7nd9u4/gmJsfh/eK6u
skjOtIseU41b6+pBfszPp1J4NI5GEWPPuexvN3+3DnQNmbJDZGrFnTQoN2nHPFkG
YSPm53Kwe12C/nYeO5EgjBeciUA59xKiDm6FikbFSlUGcpNkVnTiz2+ZSoU2FP3K
PqhCm3J7wjDEaQm7YlrTsyQeOj6VNlTSHPc5yaVlQwMGvF/y2vgut0t9asB9lqVI
tkVh8VgLqq9R86JvLZHk1LiciJ7K3qLgjSV39YGobQ4D6hcX9h6wlVqa3V47YRor
WrEqAjIHjKo0SooNTHkeqMT1+ViHkPhQAmI1HEs94gxwirHCNwUjgnD3JDrPNlMo
ARTvoQKulM2uqXx3BQ4Ew+UmxpDuX5qur61Zq1x8k+t/EpYhvEEOxNw9uYH1D6TT
u/vXmB1USEHr+QsOBAHto7kWHxvagjVq9Os1Wk/msiJILhlQ5f5K+hZ32kj74uLW
259TWm1ipk+rKfumMrYA3b8uw1wBN7RdFkySZ8BRBiCKhactArju4UoxTCeeVPsa
3U+9OVkHJGMMBRjmWXFFc36tryIH2T8cOMrqqViPvtwCtQy1cCy1Fu5Hl543tY97
uMWtka/m0wOIejTUkL6JRH7RbO/C9yoianztUxSVxMHeVWIGFEVSDSJT7EAhX7Cs
FXLOpO4E7o91+Di8ldbhlV3vqXfpL2IKhWm4av+wnj5AoPzMmviAz60Mr0aKkp/5
Iu4XuzzhxiX/MNdLJGd3Q+SacyR5muNuvjJSVShryiKPSeY+2t7mpb53ZWWV84Km
xB4AUPlkkH7qgCWDZgwj+PhNPXkCiFTQwe3N1En/YJyn6+5pE5iVEiuhBo4L5T1t
MmxWkfXaZjlt1g0o0ES0AkHUcBOxu6XkuDl4RzI51s9JDH9ml/TzKhQ/uFLleuek
w6J2gCMRPKwuY7opFynyCvr5mIE326dw51fGkKrT6UXUJxascF9J9katnu1PtwSp
z2Jrd3JOAAx/KM2oc+0UCYSxRSsq3uuMBqMYwIGPS4XsaASTpzogLx9mcbJWzlKC
IC2ilxhXXwUspQ32JThg5M7navMm3Uk/0xHO/JKmjxDZEG+RV2xGK+S9xRNUXymX
+NCYMlJKniiY6yY7xtuQDfoDBYyxfs2AVWH2jUEz5d9AnC72adW6u1lVVmoJMUpH
5Cbk+yguKeoqkU0K+KBGRls8jJTrNiYeaWBSZuhdLqovQXzsDOn7xPN/QoUHEwfE
1xpzr/41AoRv2oUdZdxYm0ydP/Ra3Y47vf+xyXH7aK9CI0iEQ99TPCRKHB0O3Ugp
QRTUqb1nRlRJvpXyOqpoadXIJlWwvoYREfwWYrqU+XciTncMEx4BWV/7PiHH+Cex
QMYVDCIQEL8y+YDzar2K5Urnmx3ZdgVChsO/4lsC9xT1QVJlV3Kp6TBCBgtvqsOE
We9SRZoPwHEamuUPNrjjW0zRCPTm8crEorF64nu4YbT893SSZzNqUzG28kzHiJWT
QB4sxppqB/OxYAMLLF33Ggbs/P6JfxeebIBWq7p+lopLD4KcZkIvnIgnuHkL1awY
t30v9bVHO8/RbuZgJciDULUoorkBrKaL+5hC+vQYTxrw4NtRjb3s0OhncZTNf4D1
UN6aOdg1zQu5o4LwwGwX71kDumw9NND2L+gsf6SYoJ+LjaEm0hV3IonkE1gE2onT
O7oj496jFi2/v6q2GTBixJTs5SBjwZGg31YF5y1idn5RlFmenl3b7rU7hF1GQDRb
9NfC9CMfsCuYTh/9M1CzfCRo663w1TpySi8ZDLNBwsoz+GISvNa1t/sfoEjUecVL
kL4Uvoz0xbgR6hXp52sEpyv8gRoTa3LFA1dsyedXN+L2pWtzwrKv6ay0VUC4MvXD
xhnoR+W0MWGS/0MiaNNrE7f5TCvcldbAnR8Jm+9GNSfVumvCSlYfrJoz6qiRZt0j
NLhmYf7Qk0utWtqojjy0QcZw/g1zWXry+BS85F4PNl+ROPLFb4jpme0s/xOnBjCx
Sxz6dMXdRMOMEaJ459Mjb7ON4ANKwhzHoJFR3i96I9lWBjMJcA3IAax1lvyqX+Pu
7gW3OBvV+KQ3/BW7YeF8JPAgrimMgoBt7800XinEXKK7mvqUHhcUlZUAGJFJdVKp
G3Qc/AmQzd7wTmZTTCmukUYmN3bbQ5eKXn/mTWj8PpWmjXTFzT/BkOiEui7o8WLL
SVkmL9KgLCCNYzxSD499xud3We+4g9admq3RY6AwCpLbf4T0Cmg2oAj+YApYl0s4
GucjdLlRQdShdBhKIAeRNWvsIhNtr0iBDnoPJTn8qqz70/wXqtyW+9AIGw6kyUWA
PRcWQLDGLVCRgKBlaI2Lv+eCdJJuTCSS/zjZ12PgkXuMEBPHh4A5oTUUfjO4jEvH
4HiWdHO3ZV6UmeIPGOdolDvNGCe+2XKp9GyQmEZ4Qz1kwYEpYQTbCidfU4UdFICY
l9KiwnJKhHtvyLWgzf0SzTx1h546N3ZP4Q7pix24JyVQctFCcZXO01MAF2Dyg48J
B5HWC13avWGhexIqa6RIChywUeQmGUjTg5DNsQPRgZVfibqXYLEGjQXQjzdw10TE
bkVvbxFgDPNJsp9c/shXUp9yJqpCF91OmS3DuA81Iz8bQ18bqiL88FxX2xqsdgiq
X8G2bF9AR30kSK9a3CodqUXCX6gdCa1nN+BkkQwE6rwNH54hvuio4l7F3uLRORjP
wfB5aa446hSR30AY4OhU3hfCWy5vH7bh8L9j/OI10cyCUouDr7ywWzXRcPZdZ+Cb
k9SNL5r4bR7WoT16Z6SjRQRY2dG1cs458IC4hd6Uipoq4iVWXQW8Ngzi7Z/oLw04
39/FVxHi6QfCBpbxJKMW1lo8n1L742YESiU0lxEsISyMCBGit5pf7+sh9OSpfKrr
BILMmRRQ+oFekEHpBq8I578AdJPsNDa5BLWaRqy4ntc/3poQ4mYRNUoGygMq7meW
Q0ArbAOgwHIJxysj1nq/SSUm/pdmKTgB+apdQjjEn8rf9n9P96R0b/kDVMxW2Qfy
sPi+JM2DWGIGF3rthido77xGFJfuMQNGma8GbEnusvZpSV4IAo68mGF1PaT8gm51
HKT0NnIXneAGJsuaPVpCOGTiS18jwXKIeumpFNhn16naspYZJ8RTPnjIRQmmJ3oy
H+S32M4QnfsBbHbTFADU5BA3c3uOoUckTNgRoHDxBzjIdqdXBGI/pYNRxqVVkioI
uL6vpeKsYxOtVSPKVRjXJVSPjpdR1li81iDENpk87zq1ezkYL043EPsVY3YLtsXZ
X8oRLds+/DzgIYdMDn/ZKTGaVS636MijQfFK8CNytAwCkjyQmZRy7cOAtiWIDQ71
AqTkaN2uzgzif0ySyAUk7FFCF14k7KS+2H5ZGVsVSsiFEt8/AfggKgn8EH0p38bx
1ZieKX9ztq/odFXk0ena58/d52OXT0j4ZyuEdHW0vQpnn5RKthNl2/AFB/TXUiqR
3WM8SdQL0p8xVmyFseUUSoQ5PaCbARZzwPmRbQz5jSa8nd6jMT7PM7C+GcJ9afwi
2hlAe21ykNRp6ODu1a3JZwjR13Ha3KwBwFBpNwHmWzNGSoJFDkkvFSy9MdkUpvAE
NTMkMk3fL5sKeh1ki12BQCKbpMh7VrW34aXkwLAyRm6PJeFm8bmKDJXbv3MwUdg3
T0utSH4MqKoKHYGDsm88ZP/oJhYEJgbrKwG3NJVLTWoqTNl5AbnOb/DPZAUvzD1K
1DC9JFn5fDiLFJXVuSXedb9vZT1cHENwpNzh7Vs95QmPdM8IO22Rx3oEZHRc4Z3R
Af8U5/oFlZgmlQ97tFqFYh8QXtmDgydkP5r0/Q+KUyV+tzZriwYwRMqvPRqveKp0
1Z0swi7n/4HxBvDlIxCme9OzjxmnElh1/QZ67xZ0pLaxD4G+fDwbD46o2sKfoipj
iZse5P4yanwqNqNyQs+72V4wEHGxm3k+RbDFyqTSrrX/h27gJ0qysMl6n37+YtM9
mRSVX+E3UZ47rwYNdVnEwDhkRWBq87HsIiwb1NgyX7DTK8VDqz9ft2VnWmtOCNXs
ulaUg9zAIWamXTGnzGyUNvhrVpHTFfqZBjiENmP9WdOC30rr9scCpibzIHybKJB/
EOb2z2E3aW30+9DsW+r78X1k4eK/WkYjmlBpfRBCDoNHopn6BXqXvszye9Yok5df
nXsTXFhKQdKn16+zaNBeggLpMjodfdTZ8i6h8jmBkTspslFR/KS7Kfc8T+uNlMQp
fuZfANYPAoDKjekbJ3+nTT/Sg7bs+uhIXqH9bwRb/BK2vECg/p91HjtaXjnR8jDz
1k8q1htaaeua2eetOfqRacxZfjJ+szBeJUZbuadMKV2CBa3fNH2qtTBGIiZQQwa6
dS9h5lepg9rS0TbIT/mQzaqbT+gR5nOizjDTOrtTjKM5LNmAjDQWW0szHxx4YD3h
oxsyLzicQha2WwS6qF5wZxGdS3sbRNPOUiEaTrC9tfBh1WUt/GZQQ06MzzfkAYil
3+VgLr4726tib0HgMUySFdpypTDX+7oi/Tin3Hu1SBoXoYPCxZ5oNtz+1qaBb7Gr
vdnqld5RHJ424pK1WdiuRZhW+rC62xi7QVJSdtTsnRgwIwu1bfnWpYZhWZVQZLev
oLKXgscQAXHLdbadmt/jQjpF//hj862QdISJEPN3RwB8o70M9psEkSdWCMbyMYms
pOmt+vf+d1jTp0bu+uRou22uKOh8rxtBoXnXUaY6l9XiWxgm4aT0gRCkAzWLAMUI
ZRlb/6eDIXQ3N69YTafKtoF+reaZ22m28wD+QhrWxSVPzSwRlqXmljDR/w5wshE7
8y2m8iprDwfWT5qdDNaQP8PuPcclnjVrN1CtDR8cg7LUY37R4ZCXy/f3WyrD/Q4u
V1yeSoDarrZEFiiydjk0Pmy8p52eUfiXMVh1LtH2gsD3XobjuGNmbjuuP5YS1Vhv
rS2B6LAOGVvg2fztlLQ7wfzizfTQIcMlBsn+HXb4AixSfwWwm2E+HClZRxOjXlyh
MuFgQ7SpW3oWaq7FAk0XSvaok+1f52NfUUK+uqX8N3Vec4ogs/PMHv/6Ur4jnDFb
YNuLQXgVCXYFuMJWvYS2Gt4DfNFrI47h4QhCzahOVGMIdKr5APsQVhFvZU/9IgED
RdGlDGbmXBnNC6eWgpbj85kesyF+EmwfvA0xfjcAKNT/Ga4WvF3yu+/++InUUNAX
kSPaeblWBIQs7twwoojnJ5JrsfBD4NBrAyih917wOwycR3icxxni+MXjw527X9Ff
+lEhmLuc4lw/ax1w/vNqJQyPk74JAk7pCg+LyeJ7BAwV7LUeKHkj66hEPelDjrVw
iU1d56VQm88qQyoG0lhbQQbwBLRqIfNoFl7991j3oXnBNlraIPbtl/gzIn73pPpv
AGibqS+RcCkMyvdf6ztAFauE5KtfoiFPJBi+yLJ1u4jFzUKiIYM6uxgycTs90EfP
c3Z+hsvLTBEsIVwcImL5S1XV3ycLSIyUc8gJGDSjNjGrUMf26mTWUQnhr3bu30GA
s00era9VfEI/7Dg+eknbfVd31V+1gXjO0+BU96DKiRJ/MZ2ZdCACrlWJ7wMofNG8
AzI/ZspDJL/OnvmtpnxhIfTddtw1pN5L95TAXklsngh1QH25hECmU4fFZZIlWN+m
QOQbMfb6E8yjYp5kW7REaHme5ww8DleRs3hFJmiCrgMB0MkaBQMtj6C2GrRf2y7N
rcxPGRYGi6hVCpKGJEor1JYbJJ19s9NhQurkeRPRDXPxLITat/H+HmcmY9ImS58T
2ty4WVGlxSD0LtWVwP4mfaP2qqYiS2/sUgT5qTfTDmwKYirHPGDopg2d5Q418Hrq
sP+0QaUpggGrZh8RuzE0Bf2DrxGlggVfLuT4DunmXRUfHLnKOpJY4ss2CGM+w/oW
1dzW8ma082aYX0cyPapkMs+HKVHYCdKTJWoRN1vZWNW29PFVoAY6EB6Vyk6V6tXt
bx4hlj3Pyl7kctQWJpjAUX2OQu7xAt1OC+L9pwGaYMZIa6HL/R/52DAUjaNPRYZZ
IOtSRs5VVQcNWI+GM4TGOTMrU0/puLDPaO0uYZEyTST/IGRym6CUN1FN5ZqTCUgt
yYyTnE6oMrwn8L7d9HsJyttNJV1Pp1CqQKMAQ9nXms7DpuERIWzKceR2movSXX6g
l7nqgOm/iqopUsp9zvazY+nwh2Vj87K3uFZnsgX9i7ip0EC0taBpwrN0U3cM8kjf
wiEnnwpAWJWQ32f8u0s2+yAEFjTEEknVnpYUwQPeYGM9w9Eey5KxR+2lWy+t3ZTs
egJXbkSOAGtcNnArarQg+rfDIWy2AiiYi2kyOVwrDrKU+MC/YLvk1MC7aP9KqK6D
ATUTVsOiVHa6hEaaTJ1O+mc6AxbTfGRyXXsCrsdozS9aTBy9t66zrjI0h+e2iEGL
jbDitL4m+Xv11MIsD9a51MkZ164I/jPy8iatTMPSON/LQfsi8uB/chgMqih2k/sS
i0BwWbcr+GETNrk3LbelAJJjclxHwFRlGGDHgaLFV9aTop5jALd5Cgv2EyBbQ9d4
zqSsyZLkIv6J61oJCCyn93sydtaan5rHEv2+1kExfA30/Qu/N/U6wgDAe7+WU0ZI
/olcz2T+k69wCI8YS2gfu6vKj8op37i74Crs8/T1Nfg4av4Bo9XKtTSkPc6oI1ZU
7IBkRY8bXGsttUjq+5O5AhgBtw4+gC2bgHc6FAE6glZdw0slgJ52OEuauAXJuvsy
8n5kW8WMR4M0fadvDx87ZNjI+I2cxasSoY9nlZtb98zqJ38n41eFGzuX4V29goxV
7+8CH2skKGO0f9q1DU+o9vPNccBA5UAEhyulDvk34Zh7V9kr3Jvy591mjxwxCAvH
VACCwA02QPj5LCC17F9ojx5D19NNQ1Fli5ccS8QwS2m0KBt+XR1gN1MVEOVnt5F6
g10I1HkWw2UagksLWoPGpSFXHiAgQBDX35xirvlI9dr+MuUDKYKAYPbNpBQI2pqp
VnyyL98wl9Ao653hERjW5aYilq+pklHfbM8tgfECKx7bCkPvrljB4oxSYaJofN//
WNHgOS1DXJoTFy/TgBDUCLShiDNg9bmE7YvNYwuUzuLZe9u/lefzU8+88RGKOZjE
RAxq5JQte4YJLd7UuWrUr9VH7o3Uud9qv9oz+FQt7p9kU4gFSThzKz6iWw3WJcgI
bPZCoea8FOjmtL+VMkk0SEtkv+LOQAVI5CSDZ5yEhpBNhNeSroKHPuKhnwncQaKF
gq1T6pcMGBi4LkxNFWBV3C1HP1D1NMgArYIOR6ASNd0ZGUeZwtPYMBbNRqlYvfLS
MWrEzyfn18Vy0bRLoKazL2knOuXyz2BjuHZmuLQ+uWqKMHWeZcb3Kz7zYfhKQuM5
9i0D1PlpzgP54tVo81XIhADUCkkVop9+XvpqrPWfl+ofRKyEV+w1uniaYrgKdUwW
aRHlo/9hT9mpbCSLu1H4XXrVauEfKBllsNsyJXEjnElaoIEc7qjkQeTsmD7PVgXx
WuK7TjapqZTmuA/9ygCJ4RfFieJHqtU5rdG9iyjY9240CrrJR9ePDZ2OU4wetfRw
JCRt9Clxrl7WRiHJqonQ6Cl7QsKHG/YDlTRSMZg35NRLfznYA/JCRnWX/iFmhXwK
BJ+EA1dsFsp7H7m/RvfF7v1Zq+4D0fEelFkHm7527AsJahmXNMlHDCk5UlZBqzZH
TQ3r2r7AJdvWoVce7m/967dAct+AwzI+Efu5LFiNf7VT4ItmJEol7D/2gc0pqTUP
zGnjjiCbVLF9ztG073x7SmS5FL3KQFlH0/R0SWce+0JlsICSMZWAaK+DnPWiOjzH
8Q5ujWcKufoMh+gAKHbBBKKg6x0oD9+TfR1IbAuR5oYKY2Cy6i1VV6y2iwpD/kM0
3dsb+UgiIRBLAWR8l/QqgfUkkWA3NcEJU1xb+aLCYXBBX/XjKe9XRfzJfH/CM2rd
uuTsBcxXaMlIrDHe7o8cfn2HFYKJD+kGBMyXkEg+y4snmSFJCJD2fOqNS0TaoW9U
9TAko70wCncMIWM2zlqAMlbOWb5kvOpJF/yrb7Z1uSudmtfjB59YLhxUDVuFCKPP
fZke0//jovJ49ZYeBsSaEjVwrBaWhmNbEit9QzfuaLWV9JtAw9FjC7kMXLoNejgz
pRVxbACuAYggOMKbfzJ/ZEOvD579QzV89Y/2i9+IMXyN8rzpxyAcWY7l6z4YlavP
MZjvUN/Hm2gZrsWdDoeQd2WfleVeGpab03lPTObGMTq7UPGs1O8r1IZtzxXIOVV0
qMe5nl4MYSrOz0Ai1vMZM2jD4TLzKOzn3+3NKS12OnwfSgTn0ff2aynY/y3APzYR
kSPEND3DkabHARTkRZgoLEVFNcVesx/PjvAhzxbuV4qw5JtdS/SRKdJC3lO/p6+w
Ufl2tKtXF2vfucjJyNdM+Wy1ets7BCODaZj5kGU8zjr5hNQqzigMRu1FZ9cu9Xm4
bujTrv53ZnQUwrhl0e8wQXP56ruvtK9upw13hNrgqnB4QCttHE9imXqkJUgQvvJC
2DpVVf3txAMwfyDp9C0wcK6yCBAEJ3fmvxGIFHxE5SWcX/O+HC+INZe7gnIV8TaH
arRTshL5dzGxAhQNeG1rCzpx92J7/lp3GPJM0a+6muRqBYFMgN9c14cwZqZUxXOf
qvgjY7kTWixq0aAyMNYYsry1kpTetdOad7l6gno7l5PMqdlZMLLMtX+RV+XgsQTt
cRiF9C7Av3idXA6ul15Y1reDnmkB5DDZoF6+YOZMSfMhBQZZ+ZYmhD/6qXndgC9O
tkX21fwqysRvATxXTGO4JGQkPV9VnwVyd+xTV/RTQ+pGo68siybHGnS4osnsdznM
7C6o53aEBExUL3TUa9DXS9K214crkzzHSHkmxa7WnA0acTokHxkxjXLFXKmRFR7o
WLxjJCx+bM66iFrSTSeuojTaOoD5kWuOqzRm3iMsStVuw8QChrGMXGzI66lHsC5i
eEL43Q0n9pZ4ngGb9QuI6fB8mpsFkC+BJ1MnLjA6ZsSCV0J0IiTpo30cs10zeyTA
Hs/+7aQTKZoOduXGYwlkas/uh9Ee2ZPdIvjzzElPH9Xe/dWsPHvMF13HRIe/J6SY
7Pk3rg8WTquA/nkFriQZAqlisHhCi3wSPdoJHQvm06XJZF85KOLDHIRYRHyaXSdx
K/4f87r5xAb/+R40bIx4Zbo06rJIkh8BtnpNx7ezyomlFEITkZHfbNR26EurEUsj
G5oBwxHVBHLQoCNuIJmdiAuXS/sWrNFIVOren0kVU6cRuvsBx+fXfvlfl4iJ4lqR
O8YsBypUBEhQF6pbprx+aKNKfcZY7eu6nclhD0uAGrccObjv6ZYBZAAw3f6s1Qh0
cX3wVBzsAXnNe7fs0lTHMFUqLod+L77SiMnZ9M6DRndDmFTeMu0ocxKEU3dq95r0
7F2PktRZ5WEZks1yJWZJ/lrIHcyY2Hm+seAU4bBM0vVVweprz2BFhTsNNpAwVaXF
XKBbRbv8p3o1n9YVGq8NbGVa0YJIFTfeoHm8MuaONElkbMgq6/JKpkwQDCfj0Q+U
m+31xrZOg+5WUB3BRHoZ+/EoGupbSde93H7f3VYoEmPg1A5eoGbThTVww1l38jMx
PCo1yic75riP6B0nFsI18BsYjXU3JInofE+OBUSRZ+8jp204fc7QHJanBVbbIcNW
rN8ui0S70nA/SLlLbwcWUBJRwtMHDXjl+4luvt8K3XwvVGHqkAN2iNsu4/KxViZZ
yIzrlG9BlKQfRKxA1Ea8SCPf8pGqLk7O4bNJKeGBkJK34JZqY2ydwJgbRbCqqy0B
M8bZmJAUN99/k/2rmBE5VhtteAPYb22rl3a/G0hWi2GrgmZ16cyWmgGLWKEV8rDd
zBnKXqC2KXaSyKJ2ZV1IdhXDP5Nly7gQDgwRlpa//EBzuMY7aj8Nb+CZQbC+d/DP
BOuwpM5GxKDA6wfDV2dDdb0hcewKPbBrJlFxBB32wGZMnuWLpEBGaDt0LP5x9sw7
SN3+5kbwl9N6SyLbFZctMUmBl4wdrfwOHbsvLLc6UMbMbrmakLXTD8p1mWP5hx+X
l9+2ZAgB2bUtdJWe2QYwZgb/Vicjl2dpR2rTp7QsgACRKmOFm1sI5FiVT16UBx/9
fOmOyTXA3nG6y06eXiYz6X+rYlEwU72azCNWIpTwATgLcXSLjw13iVXLQ6MQhswj
AXYB2hXmupPrBnGPnMzGrliUy86pD4rGYVWOCf7hDLGbnHsIdVzOOKunR50EtLKS
LHMNG5e+qv9fzAzFG/XwOjzqSmoiQsyn7fqTI44vmQv4nAApS4iJ7NNPzi/5NZLo
cYFkEG8KXwCQ1NGtH5LtsqyxkghbrGjLgfDeFbRmX4dr6WrB5KBhHlDYVnd/qlHW
1qqJS17+1GmZggH4qlGQ0gnw8TwD+j65twZjoGYC4Q86l8JYAlaZj3W12ki9tKhi
WH7nzYpwOrFXFaOg4LOhCPRMOfGvLheNpx9IzgzfU/wX5VlTeZSG+gf3t1mEEnmh
DSHLiJ1Pl7tFtMFVK0GH5p6LdQny7RhyYG3I09j75wGKf0T4Aeier4hAuv40gb9c
av5e5Zpv61v5H0y0A2IeL4qKS695/cJjoAnLuH3cjNX7kezMaX6KwBKkwoK6VFRf
Cr7ZZHD+UHMfx4Y0TJqDXrpxAqJYJ0MTPrCGyXndq0rogVVPMPAgspb4nZphmu2c
tm2tqFgGSQYww6FsL0BeUZVnNZh+s5Sls1Kng75LZaYfJ3SSf+FdGgoSQZPPevUN
Nj47BYO7RrSMEu19QTXqDQiFHoAC2U8GpPn7P/9bzhgw8iwDA590E3zRrfbRjMhL
+dhefugnT5QpfPgsFKZu8D237ZuJa2AaebM+/GDkLoAvhIs5zB9MbK3Nt1lQjFO8
a+dy3LII4lzWrSs3Wywh/06ER3PCoHSlPI2mLqrb2JLiIhPEbvIqxuUjJRPvmEKe
OGStQuHZhG4fgpzijOtni0Ub9LmSSMo/229bq1d/RZdKa/L1veRyLKDRII6Xr8jk
kae5Fu7KY9JEhqjOG/g3XZlaKbJ8+n9jQc+RnDUatZhV33ms0bwta5O3mcI5FzMy
tDs+qBKafZn0z8ejqPBQByh2Q32iq737TsMEKYqr2c31J4fSHPVaZk90EgG9QoVa
FLkQNiqXHp39Pe7B1qgPSSIqeCTdqF19rN/3NaMPPS1BCaO50vo8/2L7JZJ7rrDG
9eDqP7m7QbbsX8j2B0dovlAtqp5jAzv5+6QLpVQfZdGvqbx2M6n7udehlr0isy3O
GvCpQeTp+Ve3D+fBKDgB8EiIkb9a4Vhi3Ha8/FhTs3Tq3vKIPJKmApUZWBIv7F5H
UsH5pWYMBkggfIul4JqzzeranpWgYQozTcPL1yTIjU38VZHQBBVb7vRgF80D8VSU
noh8r0+DJETzmOiK1uKf9OHNMeJptm5el+MWwZIvZF3kAuukfaQGqkhiuB0Hd6YP
vONjmaI+2tz9GlvB17sNPZ7UaQDMLhXep2/crVELRDOdLR41aRIYPGbAb9J2bjcu
ucovtNFQyUBrpisL7UajFJwtaLvFIaOuJErGx36cRbCtY63/ojOTGEuRRJJdTfBa
GWxyLOppdxh1/zOK7QtcGrVvmRmhNSA2qlQNhVhhf+s88963rwcSWsNzCkzMRHVm
BNllwBe6BxW8/Rou3DnT4DRaA0ovmX7G/udXmr8kJYuBrXz9AktZVpwDlxJUKqii
Z5hp4aUXpndnf5w5dByxvA3v0XZ9+p+QnwTiIIAWLOx7AMHaRvIe+Rj7Lt2JFGqr
2v4f/KKpyYcwGsafg3ceJxrMAbEajBwmnX4Bvgux3ApPAiFLylOZEmZp1+MpFBIS
Hr6ool0QuvZvkdAwRq4Z3um5QxquWrMxKzvvFPfgtTe8kzAG2WhvZF4lISpoyUUS
CVGbSZ3wp8btPSMXG3vqytR86mcE3xES8OkefCRmDzBWYgQrXqliXgs3XxVVkbHJ
Sb8LSXr2U1s14ZSF5+hRQ+BRQJXtkKSRYOcL+9mO5DVwZl0UdtangJ7BfaJDPuWl
vb6VBbikSynZAD3bUp37YCKLPkkZBxpo+fjxq6gJDMadqHr3ef5Sxa0GVQmAk3Rn
+dVaDQBcYcYrONu94CfcoBKS+ksSiXRY0WcB6+JxNAHFarChQ+SLu1Sb59yn+rh7
RZ79Id2A2E48tYHGlxYD1pqv9uqVfJs5hm4k1GFlg+2NwzlNc6i7E76KzbTGt/TD
dz03aqT7Amu4cJu5LWKp7TPTczPy3Lj2CWEv8CTGjUkJS649v2RkMqf9cVZQqV9y
VNIcuilo7SgguTZMs/DU9iCMSzcMCryLawrOPmBHnZDVFkGAMZVAbMvRAyPSh1Sa
9HTJHV9q2gX1L0m/w9bkAa+vVkgJ4HuvHGnko8UYiTT83MoUYBmSB59yHdDOZwug
CSSp6sfywzK7lV9olHFeWAGwQnwpFh7nI3saUzYV+P5ma74kMJmh7O7aJTSxLhXT
gsl9Wt3uFdVy4BWD6QSOovBb3lxJdriauiGrDhGcb8evhtmOUegjfo6cihHjdIxi
LIvBLmG9Dn3lq+KoJAPJJ6ECFKg5oawL5UbLNKpVjXZqGkne2A0OywNlKHk2JKP/
6zOuqKyVIBN8mSkBW3yVq+oqNfVJNVYzkwDbnqrWqOc+4jIBvPWj/9HV+9GQUnfs
bpo+NKErYDyRTke74mT/8e6GYtK+NCbxkeGEjkTP2QknQopQ9BqKhb5etwuNBJns
LmOsmodsFo7hYf4kF60xX1BOd9Muq2Tyl3T+Aix0hgzP9RytCmi0aecWCTNZyp4P
R3lM5S/h9plSHWFZ0pwW+q3POQvlsLEcbx/aNX6UTXtXzhUlr4Vr7twoD1mJV6iY
lyQ5sPfAT48tZeE8FMnhBq19f03b1E1WN2Edj6sTs++sjz4ymL7Z68RpfWW+or/m
Td6tIR2aESP/vEbRg4qFv1hDx71rk+f32BGBr8KGC9clQxGhkxpcHrkrWOTA6BW6
RWcjGb6/GdnbalizK/SbCnitIiSxvR8iaogH/Ojrip/aP8wJutLoOmruWrHmS7Rs
89XmJvznL9GeAZ1hqZZtjxZSHkbECUTIKgpfCphC54RCxurgMPoQO+z5HJDM+5TP
N0yZZytQILaZv5Mh4ML8by8EJ7b/PWtoEaedi9CzhD4b2+splKMxg268LZQHaRua
5KGcLskdYFPHcrqQrM0cntIZpnyR5I+12x/WmJQf+Q+EMhnIb4ZVVvpF7anbUvxC
hpi8Iyrhi3eBM6K/CEWc3DlIRsqOu3JpSS1rsg6QT8TNcEfz6s4tb6LExc+CVyEC
jvaKcnBZrlPdLXVSrnDSTy3g23sN6cvGZAUIcE9e/N0a2BI1U4Snsnjno3iFRMzO
tCWHAZusRPKtU67YnSiVZO3eDql12qRFAjv7QCHW3/f9vcbHKybm45i90FHG218g
MqbHmbYMuBmJmmmRCXXowmUOHol3owBaGLgTsWPQfdlMQ7s9o29EoWxpQ7V2khcL
LxUeVt27ruZXcX/57LqBu5EVveZqJPuHSSfSiDrwrm+9bqFwS4yWq1vglyuF4mIF
lGbrmM8uXQGwL4449Vbqfx507eklEB7AZNm6dB1/uG5UypfwCWUOQNu4jVwoRCJ3
ZyX/dwRy0XnPx9ryxxd4oqoj5JSoRDqj85m3aE6QI32/9mpnjwKmCiJvUX5hBIlz
QVSEAeChnE/Rd/x5Js/kHN6S/4r/ED4hDeUIzRjwOPYX1vPkf037k1f8rgGKK8QN
ucSzUAc6ogNzKU+HLdNqodEwE9yjJ+Mp8l4/kNXGouo1MHtNYJZiv9atu4/CTpkv
FebWnB/FcYXJEB7HkLOAcwoq+ezHOk2gqXIPhVPCg4cJ50nRZaF7ZpVQMthz3VFS
PChvGHvgJJm3MWa84nKeFsjA+ZbwuiaPTW7EU7pMPY9iLhWiCuB7KxVeoTqLF7wt
E7NiYIToZ0v0JkLhdGnkf6r0zWq6aNSR1WBB0YqUOVZy0QfuiH3LcqRs+ydGU674
fxs+98OKM/AQclm4E0/ng1HPo10j4NU61hfJa9AqF3lEwZZj2z607RJo93bIOLpa
XFnmtBxwTTwcuD2OOouFFKDC5QjOpRlogG76WMKgoI8UHTY6MxmaQlLaPjVNersG
WCq48EFm3OZRpzoaleEHLRoWmszKus/GKw1aXLu89cMZxyrdB8g+lx6zYYMpXNnE
74uoeIM1eiyNGIMOViqVDCQ9m6+2PCghoEG/OKk5fRqLlxUwGMUYbkoyRnX9bmaY
ZmpqU2VsrkbVk71QPSZK6QUxJNTx1oDRtDTnHU2ku5IxjjG2ISC2kTjJ+PEoi873
z6/yOTKMQA3KexiPXhQfTOJvYgsp2F1GzC0KptiZY6qI5u5Z39x2YFXSPwDxopKL
Cl+3sxTnAuXdyIlWdTQ4hA4oobJd1YPa52EfpdwnSNmXRVnMBcBtrfEyPCv7tGkm
7z/BCgrcPy3d+j5gt/R3g9OCLN3MfzOuc2MFxn79QGZhE62xL0VrZrwYj/z+C9QE
In5QltX/4cOLcHT967I7ScCriyaVhfIaVqHAKI5PGGphr1AX8lV8mEUvlAKbZFw1
SYgTDkkGZCjVJtmG76cpCKHwyZpXsceyvGvfWdWaYHNyZBgMHqo3JGJP5uPWS5QB
vvbPtvaN8BuY8b7t+nk1fo1xSRtIm1eNv1fX+HgtbHhdEPAThRpjrWW03pkOPpOi
4zOl3OTivBTQo5KEah7w8w+b5I3cltBtwwHi+cncEmSN+RdFNmZ6sb0UQwhyYcRM
UTWD4jMPDJIbcg6rs3EUc67hr9IbBG2LopDTeUetz28+kkUj+DvoPMbjNsVf4X9b
AnSRcXjXwPoLwJ34/PJbEPEtIudF/f9oQW9fLvng2xuJJLawi23ojMagRn8ltc8J
YFuZ32P4PyLTflQjHO9dNFF1D/C9xSd43AYKqjJ6qSs+SwnsLkEjCEPfvf9Cqkqd
pXURQTjBlN3M6jlshxVGFYev4yau1+nwMPiKA8OnLjl8+xhuNI48HA5UIYgBIVR3
fK08Yus8IOcKlryGV7HkIYxmt7clTshuqOgiG6MLpjOtp4gSsRlXot7MbgDWsFBm
gaRrS/Rd6s7HvQgEt558/wMtaWvPM+NbNdhLrLBbQ5sqYbB//kMmTeG0JRuM+rro
yjR5zcDzoJfYiIpe3goa6/kY1QnT0mMOxq1zDRrOdqp2yeiLM7SlF9JeXKe77Q9f
sZkotIfEMJTqGXlOP9vA/nrU/EbbiIKfYAvUxam//y+tfROHIszUzJvo01wrxrAn
Hj+ficVfSB4JuEZTkx1cm5KoqQTdoBpFuFklvDQJFwVpwsQAa0hPFoXbYPWa4LDg
K0HV0MutC0j4j++ygu1yjLYqG/gM2ztE1QGUDG/DHaDnEIr42XDl9mb7HkArPPIa
h/HsCpxGkh8ODPfijydCzlfC/2WfBl0Ow2fGXw3SC9PlkiI/yhkkVoVcuEu/xe/2
N0kniWohcDHFCIE6RITXNPqoZ7FIJbG0TkSSuMEmvUJXI40ePHeYaBLJ7urkQXPq
QzhV3i85u/OVwqNYjc6Rr5kXDX2F3qxGWKu1Z373DiB8hWYGS69HanptUARdh2+b
PJu+cQo3ZphxtRG2EhjZRZPHsMtUFZBZUCQApu3pvc3jo4e5HABBYxThNUZhfXWX
2EolROWIS4kBqXFYON0+Pldd+4BIreZsggiQwRLpFrPafc/G29pUZU2r2GbGIMDb
GpsM1bW2wY2R0TuRs41IjNJdzW5DuNLqk3TYvv2ilOgVmgD4gfUfozsaWSZatwun
lZW2jvhwbQ+3zcuJP5nc5cf777IGRjT3uMs9JPg9hkTWtxSNTiFNsZsJubYRU7Dl
XARDtpXfd0EV2o2GdxHVyA3xVLrHICozQ1iMq14o7qHC4p4gnmjypSdS4BfgsaHB
14MEXx/Iwp5iAvkkW+z8SH9FZrGbwemyQ7188KP0zejf+uUi9xOH9OPr3PpL2VzX
VYUJ6Ilg6Z4Cs+yRgxTJDFmDBty10DQ5ubICZuWPuc2sV5wSREIji4iufHbIoetQ
MNTJ4II5nS8PXHf442W+pf6cL42wzAmT8UTA0NBrxMPyDp5oJnj8iRNmYg4e0DCe
oAtcvkqK2mjAAtyQB5Y/tujdU3BJ+ulD3ZilOkuDq/j2TBcQDbbuJKvb6PP26+ju
UfOePzKR+zwQgmHeIHYOS3sw4hT2KogFAjkFSVI7RPHyuqhR8134ybYXcpNetTU2
YWYO2D78Im5Tzh9igG5dz4LhrO37dHCVFUBcqHS3y6E9Q2rPQHIwUH6YAQkaMzJX
qOESOnIBaWLe41YJNAy9gMf2reoO6/y5AIG4sybdc9kWFpiPwwUVC2EWWT2BFVXv
Xz5dDfnBdtXB1LyG9B/7I/9JKkTS45nhLjwQ0/MPSr9k/7dYhuJzIrkilY5+ES9w
4rLIbuup2GLHBJ34pnOpCLpMWcWY6/lZMvZRm34Sx9CGvk5qsCNjKtTK+BsTY4H9
L6PL92zGTnh3FwBfckeaG/dZzxIXFc3vyKknD5HcbHidscEgAhQyZo6THdQ+7oN+
tjdKrs/89kxwCOvBstA/E0RFrjUts6db82mMTISW2FFdeY3UbGbGVapAE5FrD0q8
0uTCBLfA54ICmTdaQmdmBhVBzf2NmeOggRrHAaGZDa98XZyVynyCq+/oiEBYQj47
yr6Gd/nFIB0BIS5Ed9YJ4R5fZDDNjkwO5/yLOGf3N0vwpngq5KvN+eslji0nJ5BQ
LNxIRR7RLLnhtrY1OkaOzrszpoqj2iOlH7mEwUaeplc5lotYwFR6r7HXOVlTHDO4
eWVLtfw9rGrG04cjoUHNQWxleFFe7cq8buB6SpekYFPozCAYBpOk+f8Kyu8DNtRw
dTI+usl4sWKcEsbmbmktbknFqOP8apJ5uZBeKMpm6BGaZgQtiZIbaT7IzGIf1fyH
Zm4Sa4T3xL1QPWoTE1z5ge6p8hg1ZGf72R8wm0UJFCHgqSFUd4eE6vk9L4UrQqHA
oyQTOxRxf4b97Zu5c8akmypE/xfdV/wWNMi5JKgwF3VQ65wqwHsGHyWLXEyWRwwv
0ALkEIz79SXQPaEopLTS9Pyu+pDNaWfYfsj0i4NdKwLwpCBbgoMR+ZWDC5Hfs8A/
uexr+HE5zxOVzJlVXDyRevSuZDL3tHb9UqD+S58vLpHfXCVvLa2OnIVDlR0siFyx
F67xdTWCiH1LHxBBSqrLALctJMnoKv5fZjivv8FWNI+cpCB6Q4J3E75fVI+usHZR
qsTFKkG0g4dkmr01Ar8Ad/hf3GSU6dQ10XI2g26g2jA3PI1SbOLi46+lQ6hMdZmi
FLmzQ3hO8BDIBHs9waQecW+hWT0u8DoVuodBbBhy8zIBVcUwQvJ0udG638I5LQEY
P1glzWRuJ2W9GRHHSfrqqA1/Xlam9zBgYSDIVqoLYKXVjThhVKi4B2tsihu1O79w
EJpnbCWAtD45/1ajR5eNWm97/PkXR13Kj0CWTzO/3i5Q6QYhrbAywSykZAMlFJ4q
BRgVQxJDN3Ms8GteJd+QQt+uLfpaK/6MOJkdf26aPgYy5E4Ppbd6AtECS366wd3V
lQI34juZJ1n1oSWtUumxx4fuYH2YK5HbP6mqzgEKKmO6bFump25wbn7wy6ERXIoW
cNZEmeObUHWipLS2v7av8tJz4N4iHdF356epP3A9EleMDEfcSdy2pMGlnxcf8Uop
JgWxUCZT8xcBgbiWVdOHqA2PoABysnquI4B6DC/iEDhca0uvm0KjEOCauml3AhjY
GdA8s8eidCdGuDCQCmzimuycyi4u/b/RytmZjBMJlNh4N1CxqC8eLc8Vi7iSSDAF
7JpyuBoUlCk7EzEldEORQJMa9Q/IfJej75ufuiCctqph/EcX40R30jM912xpM/vm
ZGhmnWDG7kyP6YCqjh9pj4/58wf0JZCgr5h94tZEBtkFDDjBkCQ2dOGJQlwGinqP
vx12mH5tA02DNkRPaNWN0dGaf/kiO41MRX7/9GK687J+EXy0kjOXYQbYb+tysRws
2CiEy1qZnHbi1Ym8eOAd/0boeQ8qvTuQ+mRWEb8MPYD/5hCDEZAS9pRr8VcQ6T/A
RMJUbcgZ8lu+w6xed+FRKUb2iVysDGUZ8MqK3uH1c+rp0g3xTRQp1wBZUkJAeQSW
NCJS42hgr6OH74RDvz2v+PgZREHcmX4DV1UYA0BLdcG2BH8I4vr8TJVWCfFKdYhi
GGg2A8sxGrH+Fp+Z9JKojZsRUJhw4hqQt+GA8VuwY2aSvGZ4KCk156L4gq85HdjR
Sz/q6wtg/Yo/iQUq6KFYtMUtklrB34Yxeu29a0X2kcFrhW58zxB5jnW66Q2l+iWe
GPQnhvCT3CLzQ/a2eo8okEs/AbAcyT7HLBRNuVtCMbKAGG2bFJUkbDH0uKKOCfhs
WbLUQdSnd7iC1LwnnXTuWsIzmRAr/mb5W31saZeFpMw22whdHbWnvPPPZHIfmafZ
Zb46c/TxxvlQneTKIhwhl5jsaskEulY0o3l+RM85mvhRiBu49hC63WuXpvVOWHWm
xa5vzgOX6ep9LsJ7YV37CUbm8frRQS0fvSQ//nIPfr/U3ktvVwqom2DZZHp+yJd4
aTtts3xUyRcYw/R/T1G+weeXO8hcCdA4weeCcWjRpQeGhRFIuLOnAg2+BdAZixqh
xEttDlowt8/igqbkASfGPIoxhDz0aBKRv3bU/JcY4Qr3Bjm64zI3FVM3AMvwsvOX
C3DZFPZQVaWqn6TyGmRvvCsvBEVqx77peKTymX5UpPCgJfLFUxiOY41OS+F4v0Dm
smwKUL6cbmunMMFAwpVu3jAiU92UZ7nA+WHgT3Tpus7f5wMKGJVMJ+80W7e4yC5U
xRZvLRor97Z7oqNUiFbD6FXwjpOSYYi4h/2hUnOdYjXAE40s2swpMww9Fohq8EWH
B0FrnhBQgMXGG94EjpxWzPenBzJeu8zoJ7fBG4mo/wbrfvfQ5ShYChQ7FI5Y0Yb9
wWBgzwKVRFownrLcHctTksMqVGUiYtcQ2IcEHxIH5QIaAM9ny+GlFZkaNCYpJ0YN
7C50hnDEK1hYhG4Inv30cLWj1chVD2SywUXVtWimig0l2WeCu02Tc5+qJJgscq3d
6TVBrD4VeBpYC4+Rl2h5VJXzJ6LYuqMcx2g4UwefY4whN96OGfJ96y0Cjfi0Oo0l
nQIqFSOSofsLw2eshmYz/axJ7CRoFzB2HzcqjcoH3KXsVPNcpbKoTFf76Wlgc+ma
TUcREufzYiPXQZQ3ER/tU3J0zMnquJDTXr4LL4q3YLryctO+87c8hXptKnPzJioj
YpJODLWMYJA4SrX83xMDf3SlTpHdxyt5Zt/BZKEVkgfLfee8yPDp7p1duWqdhKj9
JCIC2wKKPLudNi6IiEpRQJz+71/vRsJijP0YnOch2nXTDgxGAqwN4oHnqV6m0K6z
T+iFWNEtss2ztUO2JgX9am7h6t8VL3bSSbIDE2PFhN+Dj7iPKDoCGxfjGEDB0qUK
ZXFiQBz9aFhfpOAMC0pzxF1ltNkEWEVR+nXXhegGOPVCKHeX9STqCi6+O6I7RWWm
Rn0MmMscMbt4okAC9fK7XhebDnjlmlM4W1l3mCDtwDx4TOJoOX063jKb+VUqho8i
CUwPmdUfwKFeRXAVrlOEw8o41wAW9k/6uGDWfVfBwIc2BxeQMyShPjiHyVCM/Je/
F8ISR/HFkC5bg4WYxI0xYakLydJgGH2i9lVVU9vSSdNm8+mb5UaM2EOAMAogZl+I
/n86qhkUfBJfsCP24iPcn/jFMCoDoSiTD8xLJvOSZSr5Kwo19oZJ9Yrt0RArrZdH
ynxBxWQOJfHjE+4OkX+LxlRFlqkrRKQmzMqi/nXgrxWXjONzYFKKO5wEHmLE0zI8
nSAkSVRvyAb5EWKsikcuB68z0fYr+T+9c8Qv8Lzpf9b3T8zkGGD+CaVMpyreJDTJ
Sc4IBlKqBe8WdpWX3v04IunXp6+pwbbM8KtUA+eDVynt+swKJ0l1Wq0S17ycR6Zp
N+eUsLT5g2XGtg8dKgmHIaWN1pLujcMe6AHOK+9z8S3h4szHwtSuOQIUAZpobtGt
mFQYZSEVmnW9UvrLyF8En9194IYHjdYDFOSJeWXANxAqEk1WXAeaoF+t/aSpZYH+
PypGUGA/LqcsZdDeC8LLRTKuZtNSjiKZ6REDgMyQN+qI8+/cUucvdUEU7ipk74cH
B0EH+yCtJozls430uBFd0kJOnMWdaGggGRkvYkmJthNxMeuu79sw5oH/Ph6LioVQ
aoMY6hB2i/c45rHKRW3JXRBm7vYneb+sP5XcELhlFN6hEzFT05bzE+l8fKLC+2r5
42cp+Uiwfu988q96jtcVibrgtJj3dQN2kst1/WOiNgYvSgIbjb5VLiSt/2Aeat74
VA9N1dEO/5iRlN5t88ZBsmrSmpDpibZW8Ndh6QlbZTrdeeuNEl1nWnzfPcdjB7Oo
duOVFVIaTAIQUrjch/aZjtbx+NiXi+I5T90vouJwFkNGI8hrfv9NoGRmYuCMf43D
rACwEKrbYeu0RGxGkO6+rWIRSmKNy6hBMB1Xud1zcg5LKQw1YkgBuAVp0cdtuejy
TPRfceoW/+wbI5T1zJZu4m+F7De7HlJPkTMSp2j/ve2k6V3UXXTkxEzIE4FPOad7
aOMuS2UehjyAKB7WF/OAWLZYJ8SNma0osYMu/uwlKC6MAycVWlY1/LVyvMjc3mFu
TJkG8u+QVbSrrGqHW0j2HMQ6FzPcnDzUwp7G1UnSl3PP+AiGptw/KFRTjR3ELZoB
R6p+E6OGoPWiFsYWLrzdxC+Y/Mf+i0nKvsHwYUwwOtj6Ho4D2PsIl4Tcc1GE700W
7RlE+TMAIYXwGWUG63eMn9ZwF/YE9NzRUVcdQThQRwCS7NAJLOpD96xznuIK6K5v
nweiobgDAAoCf6/q+eavqmGubei6wkrQbOM1h0RqXN4EblKbWWqlqWYAdqoJfqhA
kitqUTK6UaZBySzJeAurUopQk3Q9nV4x1RuKJ9VCnwnHgNFec9sBXk3nu3WbstI7
Qlz4dOxw26rqUi8maL88XN4Cg8bHqOZmqpPNrN7GcRbPS/QB2QxBrEt+P5HuVGmy
iY/y8SaEz629AC6bQLpfn2qhwodXgM0Fx3+2hwItdU4JGAHlPndd5DR4q/mv1Ifo
Ok2+LkWtE3KQORDa1tdQvizePxZ3z7TjaeRIf3jotQy1kPbQQ1I4rJUKIUwh4lbW
7jyopt4i83rNTbwT0q87kO6kLwFrhimmjIIxCt/QLhZ4bUXycsJMTPg2JmcK0pcc
WaFf/KZ3QT7eh58aYN07ZDJAr45G3Pkbt2Quv02RjfNqWYXWDlFce3Ljp4vjwmGI
0DETbM2VEOpK7h5XWaUBSXCSPA2mYk9ysIyvIgmIyNiHD4p1xAlARuGPl6qPx0m0
ydafEwn16RoUFR5y2bD9hF0d13FnvCA+HSPoQ7Obuw/N6ll9UW6ybzFMboI7C56s
mL11yAt0p0QMjvlmIcjoDkzwVA++VK94rUE63jLEWSQR7jQNwVkMYU1cGct5QfWL
1+C5HuXx34VnM+psfcratRZdorbcxT4ySbPnnV41033eOoDPYng8GFSFjnu+hh5S
hkzRrlsbHR8d+M7/otAQtDc6ougoMRzJdfjnDl9qn9AgNyZMo8CfQp7xMngora0t
o8DpQOnfs5ZrvufnQZPRWqWREgElWzfFd6D8NlR341dkkPIJMUgZBSIYOU1QKOIz
38ZyJ0oqa//mhNPYkaPrCWsy4SAPXyV2jnWmgFU87bRAzfVsqEdJFFl7wLdDqyya
arU3TZyIhH3nLu5LnQW/Bdw5E7OARBtMTuEokSttynMnbjtgPMMt6222GBM0pUwd
iJYSEFaVAGX7kVmc9oeBYypj/9SwSGllFblAn3uM/ejtRXXNWezxg4B+CZZ2+Htd
/7dK09bAa5rUeAjf0++t1cSEI86vykCL4b46xpPVh2Ut3w1/coHuAihyutbJnHcv
InV8CUkYQ2n06ny/A1l6XsLnykmJCdwK4+7zFY+X41SzyL1SpDcz2DQt0anvATj/
oMpOe1jPmElX3aZtx/bfcl6BQtRw30B4Z+kfFAZ1sPp1xBmBW7BtStU+85Dy9N6s
hv0wKPOs1SzQUhDH2t8qmrzXpoM0PtFm/EeQ2rt6U59EtCoWwdhaeiKTpVYRTRA5
kDTrywV+5FEQrDu4YdHJV/iRxolOu6GH8eD+UBhofWuKXpapOwMD5+n0ukCiMvf5
b1o0uCu3QfQAGZmZ2TI87I4RB3ecFA+vWDq3CmLfZWpzY89Dwl7KwyeNkdZb3Aj2
g/3PjWKLY0GiXVUZ9imOr6a72OLwttipStfMVwJ5Ma7DgLYYmpx0zBIcBGZydAlz
VlrrqmcBEFZ64/N7j4xJnRkmpBwLDlnJfQDsAJVSf7rPU/qGwrjE+gO2n5KWzcj+
v76Z4vLIpdQkeW+VLNfYIEhvHcdsjjmVrcvP+Miwnf4btcmuidMtGFucR5IA01s6
+caGBQC32DHsMGkHzfWaF9fhMv0XVyrjuwm4a6XiVzKvO7689D1BOihY+ry58d6d
8cUltgEepGhBUBjv5qrgP5GbtkhnAygAzvc6M7OE6qhw3GHy3VyGv43ZF5+Mv1zw
4tvV65fuzZLZiTlhlEW+PqyI1s/dffbX0h50gpyZzRKhA5GSDhne0e/R36KUD0Q2
6li9YzHNVYpEvFyZ/k+cF780/YfVb4QAjlawWyUTEMbkdvCivxaWR/Lgi0+LK+zb
F7XxEbkXAnq+Q0jEEPqDPvaeJCjIvPD7t/AFktKhsGN4Pc9kfXbA354M3v0ARw3m
SxNHCr3h54Nxiudm7M0ZlAq2/mb5+66LMBSM06YJgX3pyryquArdZxUYeeKWvkkK
H2xhz9pjGRLGnn9xHpHpsftzVmu73nohBub3+Ca73RtjUpK06aJ7TWLk9b2E0q5f
aSSKacHH5Ci+GqeYm1HDcj8m1C7fQpSDYl6M2SOw8/jlzguLMMfAwfpcEkWmNV+D
AK+QtFsnK3auLOrd0AZ+8nPbcF4hI4nNi/JOXxdHt1pZsx0cDSn7Tqk6Vo+Cl0zp
bBLhRUH+Xds9l8r5IB2OetSvruARmKVZ673e1+JcFQ+zuxScZW3GVT20qljwlMdZ
pMxxg/OMwJB/5F/2/bPy2l7N/zI0MYbIo8z60avqocc9NxqyY4+Zdx3lNze0HWFA
72Iyx7tg0fVXItlettDXTnplyOsQjncygnOY+HgGqvnfcrkGaR1dBu7r8RN8BNba
gMuVkAJ2/OIWPz+QuEE6z23LvmlQsKgzotWpT3JtkUHOxnsRMl3ppseV4nIERCAZ
zxO+MK+94de1IpTDytcb5yfoCbI2s74rspJJqJ+wej1y0uK7o2vqBslYXn/0KrVO
nasqyi3LgE3AgWGTEn1AR3pomMqVVEqWv8SdrBzwtEolyYdQGVQAyNLHfw7Ep8h3
TNKUkqW7JSttE4YB4O+h/9yMUnu1J3EO/pMiIx3CC/C/HHrnjTayI1hVMv03RJtF
pq48YvUvSsi1V0V+5KdVDB7SyohHxACj3njGPgeN0HUFBSSFjbZ8xi28zA2/ZCYW
AnIkHoAHHaE4JUP3noChvePoDg0zZcKt/p+UEtVuXdmyucB86XAdFUC6GCSjREAg
m0HH0i9hdCNIWxUXbIuk9djsON8ymrZUBp+BBWCbun9ODXpJJMTyeF9QLp9RJCeP
l/jO2Vh/1YAwxK2nqEx7LxUU8lRDzAezMVmHjmvqDsOFypNMt5nZMKs1zNYCIYIP
jUQ8D+EOBLBPQv61Nx/kBq0+Fupzxqj2QhWDAUgz/JP2HQAz4KnTGenETRsl/Zg4
FbnpHHRCsEjg2Am1L+Rmb+HrrwnjhQAQgwToHYAzKi7OtbY/kT3PgYsOgOxam/te
RWfawhJ77DLQmC6gEwuM1lPgfUfTY2sGKGrLH5t/Mws8V5k+I1LcNhHSgPhEFWeI
trDvr3Wqeoguwq0sQ9b5B8+Cij05v+Ri+pVPEo7GGdCeceZCPZ/A6Znah3nRtv1Y
Wqt5H1cvSOAF3T7kloxvLoLU7BjXAUq5JJ+OWxKOvmCskDYOFWSaGOhALrl+4X9K
FouHkNRZf6WAJxaU2GBbY8AVT0P5OEQiQmWvz2RjPsBIgDfUeGLqEurY0hhtvM0J
OaNB/V8hZ8cOmcDalCtUDRCTZFvPIpjFHCyinSHED3tOX5LC3Ddp6+htM2vLknBl
Ivl480f0G/JTrHbQtguoLgtoj4uQma5kzTTMT4d8Hdx/KmP6t5PZhgkj5XOertGP
86GBrrUjGXOd6B68Wb9naPnAfzQDKlY3DBIO8ZIfCtqnM9QU37jPBSoUSyuqf+z+
FUYjLfDiPtMS7WPOpUIh6yPVSP0EkK1ssNSh3Y32WaceOGg+yHX53ki2VON0nwE0
gAfH0t5Q4tbMjbGCjLGR0LmQz7Yy0DiPI8ofmxKdRoW1Y4PvBPormhdyi1ir6xx3
BqieJwH6qv2dG+iPFqos+RW3yWZm0U5gHQW6Fb3E3Q+gZKDOD4aXRbjdQgrOud5O
RFBFJvBWjsZCvfiuXbOc9cu6xNcNlHZpPwK01nEyytrcHnFv8P2nVPVjSQKuOuWA
KozF1zQlMcmLA27weD3rPHhHYrKyh9Tr/RnUx4+1lpW0NGAAHJss9zQ+5oSy/Mkn
65p1ZsVLrML6z/b447tyXa6eCT1Go05xb3so/sfzG2oXksEGy3dqharL/Pgrgs1H
9UMQ0fPkw6LpNIBHnOMDHWuB1tS5/RwBC5awCyFsSuYjIlx1IMCXrq7345YPrwPq
i90Q57hzcY0Ff0aMUSVJDdruo2FyLY4dnAWB2gGo6CFnF+fimXZIURDBDhQdh8Vs
QbZIYz/vsWUNO9Az1MqVC7sRw7wARWFrS3e+A+lt05aRo5xqXqaTVNratX8/gxLo
wIAheZwOFFQ1Ll3vyTkx3wmACICsRsEm1qWHDeq9WVR9t7aSgcahFusFnWVtKRQ3
zZq3411pUf6wdeEdD9Sh49XbWSoFstmwf3qHWitMP1Q78QtkJP3s/La13fDJt3RJ
Mv1qFM+bKVWJhN+eIvpm/+Zz7lOSn3lDt5LxmkciFikLmxbuLLYMEZ5rfb0Zn/2b
bxbwJOXLQigtBle5RpPGmBp0HcyEfcJYlA4JeycCE4ZT9aJffym05+kF1fLZpdp1
kf1ZGQDoTnhxHg2LkfyZN8QHbsOmwI1MdeYfK4/vV7O0uz4epJNMuxqdZraJ37VA
ADFpFNY0XxWPk3M2VJ1+1HeiQ5LsS/8Rcz2TCKwN6/U+qnW42V6y8Xz36JV9Rxc9
gZt/GWBcw3RSIfU3VdpPMdjOTbFP6Gejzu5Ra0ZIlFEtmEiSa3Dn4f6nwC+gZXFY
azO85PU0DGr4e4C4uQCIjrrsRxZFVHqXK5ko7TIQyw67PSRfBIiHF8WVMwZp8kfC
DPnUJNxadpKctjObbyerEKRC6QSsl31FSbr2cQX6EZ9EXEAZsVysB554KrdGdbmz
Jo14qu70XhlC/ra+5BcALyD8rdJ0aPpXDTBqWbWb+yqQYoGadhs0zo+v9OTy0KyQ
/yOvcYHH2VublDaTxu/mQClU3taUSIyH+noGc8MtGN8pKcnveAPgMjvfXO1IQbc2
gBW3SRkLtprKp5f1J33LBhgyYnjkkb0ZGMXHvf0Wry8WnqEuIG47Z3qmK5EJypEV
wp0Yd/rM7awV7bm4p4/o29Y+A7QoeAN418LU9rzWgekevr2zALSMPDcBmYHfB6Ra
n4KXvc3RoWekPl84IUdI12bfjvE2uYqvt/fP4e9PvDnOH3DKz6+sxxwobCNw3DkN
jJ+nUexCfcFASF182Mws7k8uXyA9OemC7rQVLIZy3MGBkJm4zMTYeXUXWIGPCfGu
+DiLdZxS6wsHN7WY6fzIfwycXVE5GHSIhOzMhIVKnMoW7XemOzpgOktcFmawLInQ
WTXsvlLlnRqTI3yFT8NYN+xUYrhnqr8AIATKXn+p7UZLtoxWqUtlQ9Q6wQUAzO0W
leSLfnpI9h+RjbLr+D+Cu4h04EIO743I5LHy7KTTIP5Xi/vI5xK/UPfLDdSN4Bna
KQyfYMhbVtXlgmO1RH+tqcftURXHt/ybsvPrsWTl3qMfACTE84ZZ7wPTPqrzP8OG
/A23VhcorufWnVyNqJT9U6qWgBuXMP2DhyqPggiplmipHYBPlUWP/vZ7kXNWuPPl
PSDiLybtPR5mCTfc1k0T0iqd3fM/Wwr7J+1LfO4zVgy1Fu8OF+0AWfEkFCtNzUPt
9R8fwTfhsS2kVkrOundGyI8784kQZ7JOYgRYIPCQ0L1seqRbsE6VLrD7h6/Nmq4b
Xvp6Qbc7yOuE3qr/PWsV9H4Mha8JuZfeDpoyl8GOyib9fzbddyvqvNxNTYRH7eTs
/RRs7sZAJO4JSQ0WT6/Yth4vHCQRJmWNDy3mPV8HCSkLBVRwfmUaWvzjdGAfalkz
1n+IfTjaoy6OzPO5yp90yHOwWZmY+gl/Ab3ImJ3Xoit7XiKLQ0IfHeeiEdCiAkMB
DOJIhKWD6fwn8dt4uZjAp+NkC2a8Lj3p3pZnFhd1HoyPC7cxY057kKXjybZtoUC+
c8FSXPbZ+2zmBvcs1LU/afrR2NLK8x8oBDYVUC4cOR6llAi3avNk8zmxGWFSRsxg
HNNXWLWvqc+w+LM/8CQOkbQRK98YemfStyKnPbYmKRb1lYtW3WDHOBsU46qGyRSP
7qF9msk9Dz/NwQTq6ck3CY0AUw8J2fXJwdvEpG04RzhhIlpycTG576P2i5I8Z0ta
b2g49dOkgU8k33GDtaN+TGxlhzznGpjMVhFlL0MPnkYdvZJJz/CMZQ/zEjecxyWo
pCaU4XPEDNwwUBK6i/8Y6GnF5qyGcuCz0s6++SJGteqoTnWdE2kMLSgeSEcF0T7R
oy76JP0jRFIi4MsBU+F58Ir4f77UtVlGYWQm+3HuEIzz5naeR4KQ+uq2C0a+RN3S
2jDIwB9DMK+lHYL6LehK0gRmOZ3WW05Lt/W+hDUoJBvDh7OKy4YerU3MeGLcLWZ0
m+/x6yRmKGmbsH8fAHlg3xShF4LTl825BKimaKVQYLMN6PBMqRJUdkHAgjjOBH9Z
zZe5MdNpdRHgt2hUgN01lEHTe+zQPJ/yCJstn5ISnJMiaICV//rN0bP0v9iipTTj
nW1/j2GWcObTfu+FrxRX4DkJG4o2GUpxsu30ykkd+jpN4tqyfBYXqJQpgRYmDXCl
kGBuhOuizTnc5nYIF29ZD+aVVkYDIbQrxLyF6+xMMFlJaPvA7pLGKtRUsvDCkLCN
Cr6nWA3i7kVt7cw8VvuE0RdnlPbT6Uy5tWJ4I+hAaoAaWPCvkjH1H6FPfpgON+i6
ZZoG3E/qCz1Orb+fVbyP2U/5Uj65kX/6cIvGRw2wz/EGYGpVkAd8Y5yX9wwE/zEZ
8ysfpTV/TnkqeiDZ5Ww+T64B29KbJkg1xQXJXjq7CZsvR618aRdZLznskgYVZXA9
EWUI+T3HhhK2nwG00FPBKFf/eXtzCCNC+ht6doiBtlb4SUZxbHhjBLOGbStFeyD2
pUBg0hebyMRmjRrcyCcee+j1yys4u7L8B/7Eg+r17P7vmgByTxPZqznFHU8U0dGt
B9axPjBGAEZIyE6hUSPfdtrYyKBdTnhbJBo/iRnwVJsZHz1lOqG/4xT9Hi4JhI1E
waFa6J5S/obHmOSfsXFely4HLzefDUF7j4SxN+NKWWLIqOMBQ0RXmUHzmfsp52lk
wZ8EfxbHr+0nDOUBEP/Kab0DHZ+AwWL9aVfHglukih3aOwq/W9FhELWiIGchyCnP
RZ9zQr+9+JNpVjAT5FduqageXkU8u8QgYSnFxb8UQKGbxCI32q/rGsfKiongMcpR
FYu3rz2ELqp2n0bztrYIamROwkqypiRLmjtSDkThsLx0y3N6YShPIjdqubkEDIrD
/XsVFHFqIx9kS2jZ/z74XkOGwG0MHpTysa86O6efaC7qccezaVQKQqKcjue58daw
iSRWseslBqqNio+HM3Uncddm52uQqZwHOqWWDM7vUFjgtn/gDT3Z7exkVJLcSgMu
YN4aDksXnKu8bkVLfSmzEj3QDcTDAZZqpB07SaQYPqC+kxFPdHGddKhruKpmLUAG
d25ChWZ/YvVHEvmOCJqwHikx0dRtqVmDXn6rzNhtdDpIDnBmqUR4y8tcCw0BwUL4
eXg/zcfvW6ZpT6C0uV79k4YI4eGWG2CzMGWbzzOQQYVreVn2GholDmgL8efXzVi5
qhbNFjQsfFfm5cl4LcL1Z7bo9Tlp1W71p2zPp0dfw6rXQAbsf423VOPxYALEDIzI
4V6ArzhqtcxAg+mzyTluP6pSv2TF/QXZcdqJ22PICIfflV1xP/I3vtY7yHZxSJl0
jmUr24wj8TKiOmOYP1MUO7WcyCkeftGy5QAm8yz2TYQ01wM1+8QLdoH5bwFdaoGK
GIbrrHXTNZPkQfSjYgOF5FMh25lzs/QVfYX9AQAFHQ4cTu+LYH5fSn40apOn8dul
p5dtAws2khcBCOglAfvcypREyaxhuzoQEZVlRzfTbQVmYxgXH7Zkg2TSHzFocvvO
QTh9a/ySrjM/3Ill9FT9ypNMW+DNoqm3InXsrgHpxUHRy9EUTqlgf4ha+fSM9C57
uO+iiR2HeoARp7Dp4ueleHVhXIVU+iEVvTuvRVw9fAsKpgxJwE9hkwo+8S2ZXVWi
D0DW+M+zNvDCbpXaYxvGqtKK0jagqzpALgJcHvhlLrO+61Jlti11SWjQXJESnbip
lQq7Ti6yxy3x4os/OlywSQVG5yWNCk/UOIm93VNMbZEbXR94j11vRpTZ1BhBVVd2
hbQ+ZP4sJkv5wXfY9p3izEg3bZ6x+kgLa+T8p+gLzCDZitPsZdpezih71ZX1w4h+
Te+btHbKCzN1ffDgrrRaVLqxLA00yxSTWPcPUWl6D9PN5V1JP9Si8fnCYXZUiCwL
C9Bt53NIN/Rf9wnhkkXxWhf/+oYoNlxSXEghn+j82E9vDavgvR9cffKroh8tYSzG
kwgRS3wYlqfiTv1JhuMfrmFyj8aS8atdgL3D9nDXSjFOT/mblUpcUBbLaDWQad5z
PcTLT/WbXZrg/n34MN6FxO2nHUVZyDYjk0aMI03uPK36mqXyMkmFt2VnXlJTJDh0
DgmB/ksmgCT7BByhoOseIbTBOAYX4JiCOGJLbFZWV5nfUSSaewe7HQiWskEJJ/Zl
UX6+CUcZeYnveEkhgO2mXvKYlEZS9c1AO4WQf/yi/7WDyGWc0SjNpJ4WaYqjPtCQ
wU28oaRMdt565BUgV6yoXe4rseU8e6cPaZDj+H6zEjr+NdO16wS538+h+nd7hY8J
bF+WADdFk9T95dtWSHCbJ6a7KP6Igpbks2OdMmI2IrZEj/lQPT+m3fqKfAnBHriC
BPYpkUoX0c1wvGUvAhYfKuwMWtFIKf6gfyXmMhDrNY8pUW86wDLi0fcWIjr0/Rte
11KrlSXBP3Y/bgAidvhYqDHq0/EPCuhLF0JwfgDqB4wGd3cerhGToUC9I3h+mR5v
SKlu0VjY/puoKWV8e8rvinA+jy7cd04RnE+2YfVooUt7l73VBn5JFJk7giUlj5h9
sY+5kFimW6Fetuhel9/1NNrQeafD93+UjH5lUJA2Jccn/1WruXCQRHAl8Nw8SW3k
WKoWueii1Sjm78TJZ3HRku1Ha3DiiMSDi1qTRGkcJpfsJmO3knzNfo5WkuwZZNon
xthhDiX9gf4Vv75jWobXSOuinbfqKVkFJiJbV12dYz8U/pHttLOwVzCTQXEAkKl/
vp6Nu9sKGRB7XEUeKc6Wq2cfmNdKNH8lnfD8JAgr/01LVq4ZxWlfq4soQdUbJOdx
ggQ8MPm8lv+GSLPyVJjP8xDmSKoTfgxmYF2VuLrO6xQhAi5ioVQRsiWAIlCzuCm4
u8Lql8G7iJ2QGPimzvoUzD0iLVSMM2WvtOX/91T3WH/I1wFVEtTl3zNDW6KgYwFV
jVH4TtYzrw3cPJBAgPKuZ+t7PQtCp5mw8pyjmVZEXRe9RC0MvKbcwWlhUZvWE1Jm
hFt8pEAN7J4nIEDWiYyqZ+O1gVx6xxK6lKONVJE7K1RM8lOppjSNxMoBhiguPKS+
zv/SkapnXw9sQMqYXWHqorkDJALmNGwU25tz0kGm/E2rxCo3LJibLJYoM/qPMwji
K4HNUBu4CkSXh1OdYa1r/jJrXGKk4rRuFzpbwpEpoqbJ+jAjQttT48q7CAAR8ItS
mS7k0f0mJCs1N30ZTC43X5fQd5h20vj4X/QUc+e/p/W4nPEKweBb0u0amr3tFrfK
jJb7ODSnclyZj/LpsrInoW2jqnWl30h83e1/eosScEnFr8pAGWsLSGB/CNlruzj+
Cs82Z3vyR1LWYp2qPSj2rkcR5P9FXhdZTtrr2EiVOKSApepbYEgEHaO3062F6qVW
y5JWPviRxjxF6RJWaG1OdYtXiI2TxK/M1dWZ9pphhc2Mz+6j60T8Vs5TIgx9pxBG
zxyrCoE/5pl1kip9ItR5cij3Dcrpf6zfqkEDxrXfrArO0rzgReMnHYdgpUlAgyHJ
mrUeIQnLztpg4+R3o5/iNQ4m8Phm4O7c0RwMA8BbcE8CcWqWdwz6K9Pgj7PY4j9n
VhjpAY8+A9A6SkTjOa9s71aQrTnbIf5Q6xZssHOQhLZyKYuHacF0sgVfdgeK6oTs
U9x/HGdT6Td0atYPZEMby8dKmC/rK7PRaaV+aJD4l9vjV7nEJu1OLnqHofMX6gZ8
CaUeVuZhY7euQ+SODsTe27WMqGWXOheTHtxSZzSVZmRsbAvRcfSBgOEI70aNGKFu
jyckXSnAfpbwFoO7u/nuKabHb6OWuXr7OhG+AwqzCM4cBTdP/JWCw8NYxm3NhoXb
fW+gSUbfjWKHwgouqYcd5IsI8sqvPIfny+5Rkhc9b+y537eEsIMAUC4vFhI/32i/
iaD7WN2H1DvINlegHU3PF/7lw9aHFEXLiH01eAHBTm/LenSSC04SAt7znG91tW6X
6qYXWkASRYp8+3twzA09eqMhbp48q6a675pDAiElrcj1Uk0IlXCpBCn9GGgr/jgl
id63Dj1rC1KOXtLJKJgPkdsxCIeNvNREc3Fcfp4dj8J1l7yeKJ15Ylb4dbU+LR3e
lfvOXL8W69oICSsexJFG+0d0bxNb7a6M4YS9opaOWDBpjSl3Siv9cLV7rsOMJdKB
7dENiyAgUjA45rZP46YvHQL6xzrDH2ZQN/eNVILJZuSRP/NaLtTgg62lFYvjJIaX
9Pd8qTJWDBrGVIG13tQhdktmqbKXOXAmyDVncbpHfp3Qzz4w1BQdx3iMLJKe7DyP
1KgR1ecuhZxaaSQ8h2O6igQ0yyda1uLyIWNNBuIddBC1ghZ8Ew1kf++cOZHWIaO7
UC7et4boIgJvqlrbEmA6psJjz7y7UHqMgpXnPG9nXquABiF7lNcuVFU7/hfXVI54
q8J+uDeRA4bll+KlMT6IHHzaDsurgdB2ryC8JknNGjJ/q4qsqpxi+K6/ptQmPsb3
V0Noew88h2vu1W9Xbt/vWPG1/8vJAW67/VyPsLGI2nFyuVIUjogaS6gHetEelbWz
XoVuRiMCahwAehSGtnIPgUycUlQz/YOPfAMPGllmbN87a7dZnQ332ZpbTeCRIq8q
q2LaJOcnX8NWkhgF5Sxk747WgJaS1bLPhi0SwCFOrS6EueyTwd6h/AIyky6O5CEP
SUvOtEW3QVOlOXgKqIWX8mAn/99ea6u30mm23EYcRlxDCkQLLJBaD8PCbBJBFDWc
0KToPVpPR0vhqqbsctQ/mDGtSxKx9Y19r0HV/f9Zr+RpIilaceCwNhPMrBdjENtk
6sMevf7BX8JyhOGv/u9KAj3PeMksja1bm0I45UOx+BkFK17+0PnNJdtsT7QOO9rh
pfWV25B5Q9Lsn/xLbuxmcqvTENKLoWN2V4pBkScbMb6EY8IZdUoA1Sj58gKnjWBG
/LZIJxJ4ebny8ERKsgFOBUEdu55UojEvhjnj9mN1QjDGRuHVTrR4zGSeOx/yfYUj
1gWGAt4uyPb3wnChBDFs4lPUWxYb4xZXe0/9ISjRYW3vFcsuasxbW2ou119pz+Eb
qNghwDffqo6YC0s5on3qtE20nrnLeHuusPp0dantaQmeWm411ybr1d8hMvntlzxR
Wl6bN0CBioc+nf/p8h4opoQNYOCy6wFuyseo1AIdfDIHVEtrEcz0ZM/ekQgTlO1Z
mHvNwl2bDRgRQRCLq30k9Z+JPzT96AiWSVJt36kOB0SUV1FeKTWwMWpJhoVT7SAB
e5EXEFIhV1e743Zjf5UF4Lhz4keY2tHEx96dTDyxC9OAms6lU9z71R/WqCuIy+Jc
dYN6wfnBXmTYEwKWMZ9HcLArZqJVKldeEV+oaMLjOTOpZjhwiOwT06gzNDi63y/F
6MPPpfTDGGB8wYAptMeRXWQ1HyOM68G2lnS8dtcrmh2an53cPB/MRB11mKcDxgmp
XnlGm8dOfuuk8MHWxbRaukiqbpr2JwRJxhvKuHrU4ZKtPWybVDIf4w4RsfMwoUJs
PQGgU9ObVSbtXvl0PxURM3khGZ1NPBL6TWAW/VWR6imYsyqAZmsz/mv/fiQOV8ue
Yy4w4PgyNxIY6JItBtvJ5SnZC2ncywKOw+lQDsb95apkM6+JxTv0Pzb0zbkZ9+14
/GvGI0Bk1fc4d1t6fqlZXG3MOrG+vKSpigSiP93ALx2nf1zPOGvyccGPHKgxCiV0
u8OfSZnsf/TZqpY0DyhxHiSv2lbEgtHZT+rt7lXvVP1pnGiswROLodb/W0wVMiPB
eciGG1Awip62W3U2sna79PZYRZvItkblpcOoO9tjcpsX10fAabQAkcSc67l/L3Pw
zBSaEb0UxO5mctO3/u+Czovv9MDOjVONKHa6MKcXi6X7RytLTQ/Uh75mplNev/Lp
3WJBQKgmLnIXzQnC32xcXnmncLVzLe/Yz8zm4nwUtSVeo27l7E/UZjCuWlQtvYBF
I6HW81hDmxzMHrfjYrs2rRUJuwKbJhp8CDdorHq531cvvJj3osF+da22roF9qVys
FTDq4svoqoMNBx8KgwYqiBB5XB/rGnlMHqTdu8zY4t9eYU5SCjWWNDXWAB+ESy6m
g8/mK4pmKJo4QnUzhAmyax36oGLsoc3SZe6XJmc9WyVS4Wg9sSQ/yIiXausR3KTu
1KMODJxpiYoTtLrGsA/QkFJmV00ijZZWkRBYrnSt/r+fT5KOAkDmkZi1m1XQTrc7
BDedLa/0PoHyaCZIe+XhKfT+UnctrGcc9w8kXep6EbOZwD5C3YNPZ1PsBsHPtuMU
Iv0SHSs3EQws7V8v2YOR8j9i+J2QbKR+4lp95zSBzrDXQHV4/Bvzi/QcqDjkLCBX
17QYZhNwQV3wvUcRXGjFVQfylP8pgUpMvmbGSTw+N5VMfkXMsS+HFOhuulaVJ/Iq
Tdj0XbrOThe6bqOsVB9aFIUcXHQfTYt+uUvpq993vR+uyt5RZCI5sKD3aB0AVghm
6/NvRglaopKhVDufcl7newtsR7DKcpmtCQugl5H0KDWAfTvD2hcjOFZCATHxpuzP
uRg7w7JQMs+wPNN/mbiYmzOCYUWLEvQasbJeihAyeMfzL7/Vzt6mkREhTAnlnXnF
kjxcPnOPrJpukxRYfP0R+8w1nphKAlbKSmV9zPn+hqjIX21BdYoeSckXW3KC/tNv
MsMQY44XC5Hx21w/PFFoDuS7no8DtHMMKR3nDNNuq4/a6xh/jLIVfbM51GuARLtM
uX1M/GcCx0LwXwD3BzqyvfomM85l7mg2SimwcMRLScgkI3Ojt864PtMWkfDs/ZK+
hf5cfC8yZF3izQPx7XV7E5bt4Jae6ZCi9JqDr3BzRmNtL8AMT6UsGDp5+YpoEN2V
7WLb+wzvDejvlOCssoGZo5z1GDszMlcU7FcgF5H6uDDmn+pzpJtvVGbjQ+vsYoRN
waTVOe0UeRmh8GKMGoLlHhbALbr3tvMkiziAUIzHsBobuhhtYy2JzjIwpXdMSbvU
PO/dcqBhtPpvEVCU/q+3XrmZKE8MoAH7lVg8TG4s/r0JBcS4r8qYfLhxUZPPinsT
phSlXXYJfX9vLAlcXe+t9PRsuFdR396jgGcEFCSUy9pUH0kp00HfKhQs/Pe1KBi0
8nw6SObcy2Cg5S81vbo7IYJ9EtKxo37WlyYqhidyhUvfWLJeBPobu2ETlipSe3hK
pZxnCiZOIeGDpiBy8ORZEGzofSmOhxLL7anNrPN9B4FruqVSMfXaBpeJyy8CHlaj
7fNHv8pSI5kmFCY1K/cKSaylBMSMK8LaqqQq2J4boqyApJ0yTFWV7W0IdmmlCgj/
ZgT6LEWs/39VBdw4gY0F11ciRRJ7ZAfWi1Ss0vKkRaXmB77yDX5d0FcCS8rl483S
ZFvh/BDAGEu97uAvmsMF+lolULHnJ0QPhVFxOOYePEhCsEkdRpWEBYRzEfmmNjxN
7kky1Ey6QqpwBbOgiv60fExDLwfjZAZdv2T7lNI6mhLeV8lgV7YgH7Wi5qd9mOAN
IowzJja1W3qh0bBzwp6CEPzo/EaE9OdwVavU0OpEpnV5KOseIwK60kM7iKZNT5Rq
46Pankh+7lb0EXnMQgACqlJJJns+Vx5nyiWkThThnv642P8njX+8hTmnNmy9g23+
GijirOqlRJAiwtZX+Wuiz0Gv1cLKbiYkx/YYaMCFgb4vDTpcx+PPmK6AmPF1TUz7
Ft8d9Gv+DL0jW9wDWgdvK3UcvNRnbVrShGpOo4zEebsaJYXXHDXBz+vLalK8tMJT
q+ww6+qa1se6PvdBoOG+NesJK5/CqKUy7dHjaGWW+SGf4RtzYpDHepagU6v6kTGT
cw8OyaDy+wwjuuFZnoIpSbgQMIxFMB1KR7UOsyL2zqicHMzdYiDVbUe1rfi08Lic
Tm0czi9c+f9/Vb1/m94OXMai4bg51W1Sr6eftv3MvxHXnjC0d0+j0Qoi1PIJtFAX
lnCPfzZZe/cl4Ye0XBaiC5OZ620XcmR2e9eQlN0aTKZYCWKeu2u1LKz5GdYQ+N63
qvrhv0qN3yDR5L9ckwqdweVt75L0ULwWGZgt7RmR019uLpl4MK7Kwr8gODcyXaWi
OhpbDVSOWZ3v8GhdK1E7gHYStSNFzs6pbVISj6OIqHhtC6oJMTCPA05La8SkrBoZ
qFqr9MMjMjA/almhUDnybT/vRMrC50SFjH+IAhg4VN6flszBZ6qvxVMzRVO/CviJ
A9mUTXiCX47uuOLnQH3PrKc/iqRK4LbMhX4LIX677uB0e8rsCmom+rT/A6tzqlo+
HPqoPeXd/sa2l9Uc3EV/EiM64u5KvSnHDV/f6TU5rpxbw9RRrqPkR6fB8BA1KyiS
NHBnTKo3/TmeV9D4ONxRKJPI56q1Af5yg0r1r+XWiduusX6nuw1T71fbfpRQweg5
33oihvHzKoIyoGi2A8OYSflI4wnvGNhZiWJDJsBNwTpyRPa8ZzvNiOq0y0f4P5r1
NCqnsfvb0+sq14T7Qt5/zHxGf/pGL4kSEg71IJPIinK4bJ0K4MP58maZrYC6PiqW
PRADLgcZABa9gl2V1UWUSwtwhO4+1r+2mg12sMSpziy2yapMsA/NgHQyy94e9hCG
QnBMTBi1JRIOY509yuFDWhLt6C7umMGaD+d83kKEdIoilT5wDfnMF6TJ893xg/RN
pBu7y/ckI5p2RCxEGIFns7iclfb34nesE6ryZVzvB67aRJ9Lb7jTPs+uG0HyPvVs
QFQADGZQzl6woS1Ta01bi6NIzBcio7Srub41pyTwjcrBnZcaYqjJfDFxhBAItUDn
0TgUMeH7FEii4OVaa9w2NWAjHh0aI+Ao5CZeXRmOeUMmJ9oSDYuaPRmoYMGa29kI
UzMhQaPSAn1cgje1gUAr0AH2N1s3yjH+3zbO32EBH5351r39eS4WrZMyAzOCCaB1
JdpKBqebWwRhUwxyNwRXNJJqIdCaW71sabX9GsdWFncPKEGi/RwfXM4vX4x1UMDV
fMo3T1PwMEAwVBjHaJzv6WtZPSjvtSp+cKeHN++cI3KbqcknzniAfAGEtwc63OoT
eXXg20KMDJU9Ao9mT55bMn9p25oW6pyUjWqg0HQ60IuQf/JvdUnRi9Np7YaC3vu6
4pHP6V+FZhZJtR1NVRDrWsXDJoUDmGwP0Ztavheeniq5lbXPEHy/boWcNXZqxmnh
sB8fflWF5pONFxT24STxloShjYXJu35/E8gC1yFdIPAuHxrtz0mExQ+pYnl02JM5
zxN8bMXElnWELxIC/qeelCiW3Wf2mKjN/TGDNGRGlcOVBCjSoJam8o0GkWd9DGOV
iyQmsUPK7ohePqNem84ovwwN4sxVxcot28ZbJ7ht4LtOvrknU4D8Jtd8W7oMZRUy
tev+0S1i6AcV/Zsyi0ryyl2y0waFZhWK5Pc1x7bbqRaYuElzbH7iPptv6c+7k4oL
Pcx+c5RlLSdnrR5fTgCDxfB2OF5L4ipBSzqbYHGXihENScaadDn+DUR4ZC6Y4Yn2
5VVSz66oKoMKosxmPGqikJaW8pj9nEfq5GyQ1fP5ij+fDBydaaUMj1h/Ba8pmxIr
Tpxn1FJtTt4O2oDy1fXXn9Iff/JpaZbcHgVsBTSW6xtJsM3JKIEmgsi4X5TTF0U+
R44u5QlSUmvslb0+kqDT/5xDN1njumbZpGF4a92xAtwyZftSyNj2YEJrL6tIuyco
fAihTbGi1fiNdYc472AHr1TOF+yozQKeNHCspS/I7ke8Bv5ZQUL87bF592/yh0Rj
2X0kOJt0R5Wa7jtbXoUe0SN2+TQV6lfk19WLYk0MKuvuJ3EpiWoXSWuPJuI2NY8c
J2R0KNm7s3UFFcsUM7U7ZVWWpzew5iU5wEcWck0tuUGszgvj2WLZcZ6P3zyJuz6I
vZneAkF5cky6roJ5hnVdZXX3wb+PCdGSBx7KlEAhuQyqWFG+oOrasn+a41zjxdUX
teym+Gu9K1tdH9F2UiWc71lClR8UXS/xCPReQgkQrvrG3ijsqVvp9UlcDzT1wuXU
vS5PWz6WJuS9FV7jme8BcwmozbJPzAB+xrL20xD+lv4njFMJr/0AzRvgpGKQtk7s
lbBLxtv4LETGDRs41eM5/cV0XqUqELEutXY++J2wyWHfaymSMQe7tQOGr3BfM4hw
TBjZ21jXwDqn7dQoxWFp2n4OomwEBHDNGL+uuXWmOdxacd19gAwq72/EFuQQIKFD
Y4ns8J7v1v48jaNUrL3gOlJRelVeorlzEF6YAGf9hCyrB7uH5Hw9Z4iPOcn1Urmu
8ZVt/KvrlAkVe1gcwa550h7VRxAcqp+geAVd0UM9s9hOPwi7gE27rUZTafnHeh4m
LgoidDNDjVTDsuddvjvrze3Ze1Abz6mfxMJiNdP5vP/tqAJ4T6J1ZI4msVCKwkQF
xbsDWkZwY5Dik0RYqDGCf5M2Xjs0AgIRQ2m2AjV00V2mX2VVa2I6SDGuNNX0rvf2
phYqrwg+jbamJmGFhWXs2deFJYqmVaUZj6BwsJG8Lt1Vn274ZGG3zNqpQT/zuNI+
ygx9ZJebsoQGhBgBQVwuAYte3EP18AxNBrgIddWv680aPHEDem1PBG5nkfASFsph
XRIidrizAoDweBAyY32s9uf0CA7iUUeAvO7C8jmIBHCGG1eNBntiCq3L+/aVu13t
b1bM5aNK5A9VvciElnr6JwS+iVdQfqZKWg2DX21iFhWzPPZ379LNeC4LcgrZeKUH
UWSQuPwZSBodLIqx2aFJq68gNgtr+Jz1zJ0tsMLZ3R9CckRKMBML0yZ1qdlycJrS
dkT1arbOBjyc5vi8uOtzDwGviMvgX+YmqPX5y1UHbGDf9zjMYG5HWdlXfLvr7NeF
91Bpxyd6/Rc/QkslkpaVARix+AkKLp4XhmcZUd0gHpvmJxhwWh0kb5Zx0h5PVsAO
rGPMoO75Lu1/4YplM2GqujpUkUhF2zNwxPfY8yl7zPaNuK6IG4yKO3sZbhjSm9Bv
/cfsvz73MTx3Pv+OLn8pnV/oS4ELLntXZJhx+zyP4eDVimITVvbihfGRVjEnBOj4
TiM9f/YUHdpavJASlHW/6p/Df75oVZHEb/osjPHJztTZOiwpZlx/IPt6yF+iVxcI
zfMLeTwE/7/WPybB2OOgTa8is0fYA5He2Zvf0mjSnyBlCDF1KlBawHr/4QRWW9/R
1ps18IRh1iuw8L26/giKmBADbdGN4lHcpofHFroaPyFj5dF0ybCt5quQkawwhAa2
OFRze5KN34Razw+UcJdg9Ow0rqj0PccY1pqKEZX1P/rDUMV8aSQbAQm0aDCdGfGS
0kXBlvSQsg48SQZSJMGAVyn/sNQgStfRnBo6A+2lCeSex/Vc/pE7oDxze55/QGa2
Ym+cLhI8jWZLsksarv/1cnyz4jSYAaos39LsOPfBCezfuUy/H01eJR1pglAITS1I
diaziF6M8KE//ZfJW+DLKTA5PJj1EQcX8ta3P8SC9siphinI9E/LQuwG5D14p/9/
1xiVblEieIHZcVF+Z4pVv3J1snxRdDoUk3wvBFWdwM7W8FAO5/GUMGGsBX5W6Oz3
96fr50/z0gEjRNz38SoprBzH75sJvBRfjYSdR72Uoh2puzjz7mN9W7dPRXr0oK5f
Dl+BqDIw6CygiX71zIbaP/c8MwsQzu7tsyCDkds7H872oUbeaApfFeVOyZG2i8qY
GsoxaQlkGFB4fSkIO/zUCB4tO5MPCEatRaf9yPGHPGTeAfIUWkV0S0BnjDJ1M5hV
DNmAFwWachbhP/K/qoeB/vu2FltaTXgbjNcEQatFGAu0fgq9r68Se9Ez5PYLjy5e
CUQVfGmxgJARa327ms2N4VRWBmI1beaOlEITKK9s1jw4sPwbUQpPF8Pq9tGs8/+z
EfVFGRHofuRISlUkcVTrBfi9gj1d6Q4iTZZ7v1xaOe5gqZd001WYPj6Ij+Z72zeM
ByRgLPJZRL9T312eWzVqkS+0EdgG9KbdeYZta54kdBvm9/Nb4acZ4LYmGUm9n240
MzziVZLhT/qy69Oeplzto7JnC6XeirBtBW5SHWWnrUV2BCtz2NC4kQst4pa9/1s+
qUr6dAN+rXzMyL86Rm7/Y/AR0WjYh78zLGU3elBkuBeGU3pv8FkRnY8qHZKGUHnj
o2SMgOO3eavQ5KKzC3a4Y+ZA6LHlxh//Lbq5DTOEsMYlE+iw0zNA6+o0npS/+VYq
BWpM+D0cif7s5ube/8x30HtsW9htNPRHMRVsoudjhNodcdCF6T/pEEsqqsFv/dUb
IBX3QD2lo9UAvUFBc2ROawVACi0W1NCy+eZGWT4DHD+k0tsLTZvXbRRxWMARIGav
ZfTtBmA5uO1FQAZqK2L8R/bBykrwOEEsDrf51zA+HNQK1YWDHLugoCHmvIoDFh6E
MsfOasZULKw9uNp9A38xZTIK+wyD1/FWenvkn9kYZc3xNRSpNw5j2YeLjJgdYfDz
bznDQMprHSjCaJqfnskrCyP4FPvczzDslH06L//3G+HBGuRjdyu1PyInz116RCYd
pVadnSxzvJ6Lhh4geMEBYO0kZkLOeRV8fgJK4Z4PzgtLfC+5TIzvBTzY9VE0chLn
XAx95IA4n9s3viEz86KGvCtqXCBgpf5G7t0XbFpgGC9sh2rCMeJeVPC4C3LTSkGN
8Kg1PULVf5e7rAL1DQlsHvyJ05G4CfyK8TK6FJku+5lnRWwGmovQ8J+Ul2ohgROb
`pragma protect end_protected
