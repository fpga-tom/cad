// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:40 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gN75nwQUwb1O7Z2UHLkcmfqVoslFglSS0vPVVpT+o0P6/pn19f94ZzwWoID+Ni10
7XfmjiKtNvm4eDeO8IzwoeshUbEJV5JbFBwIdBhEyanaPeD5eQ8K0ZL1e2QLsyC0
n3zT+ggDJ0DxQaoNXtQMINu9zAio91gaUvp398YWd1A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22448)
ulatWzyOprpLPV7a2IfCW3WypCQOmJqDkfEvqRutwFOr+vMQP2zqNEC8z+j0Uec0
9GykAMTFXSewsUxpwEv37v88fezWEmFgjAxJAiYfKYdiwuwrfcbT4ZuphxeK5xLq
t5BguHLkj8PO/GTEmV7NiszZMPx4FFnN1jwe7OssZBux8Rv3YfISRvzb4vX9BApt
IZbK7LhAQ3FZmMEYXF5vQezTOWVQDXYgcMfSI69aiRgUBtDKdbBmiSzd4LnoK/e9
nDpYUwcZV1vyq921JxB2SWc/zYtyWexUW43t7h0gPOWnk7EKFwXuQ6R3dKbH4SFJ
k6PpzYl/1vdRlnfZ3moRRg6O4my/63Lafw8JEhhoIumpY3oMsGXzOg936v8cRb6W
qa9o+niDD3mJzx7oDA8Rp0cqZA6z6phWjARHKxbYH6CxKycu9Tv24SwPLD1uqgeh
yKtKwPsKS7n9BMdN5NULSBjYtRxKNWVGYq17sV0py2nwiVvStlqFG8313zu1zpD1
Q9SBIFv1XWY1iSmyEPyirLIcc+8wm+1z7vQI4rMerCefZLYrjAUbK39nok/Y+7b4
4bRoOOlyz20JuLQCbF4/dbmEckfMdyqo+KcR8/UXwMnelWBoHxiO8VuIoLNJtpA4
c3bjh8nK2XuW+tugSOA2wQGc+jNcFtBpBSLAS9V4ZP/6bSEn0FzouJ+/zD0hDiOB
2eGg/TyLPkjQwHPzgvArWlQ0XppURt+FtCCaGmGHWzljPdcvhbj4PelmFm+TN6AS
xkXCTGwlOJvU5gDa3j37rZLRtc5wgeQ8Oly4I0vNqWdI3xdZd7x8TB06hpKNtadd
Ql5DjYg5Vsn/01fa2fMXgMSdofkfFSdlpDR6+2U6w008UuS7b6O8FGmbklrZ9ZqF
VVHMwEHvDCBp5thMMVnJfkVDVt0nsu4XO7/xqWcY5GojR/bR/zrgIBZO2xq7uvQr
kdb7V8QJ7+3+Yf9nST3Gm4zmDTHiIGCJhGSBBrOTY+fRGfh/3inlEYj7iFYP0jAv
5Eko4WaKOrukXi4hjiqSiyn23CohLWIO/4IFO2pzcLdusrc7kX6WUS5gnTOcwBb0
h1Pv2DY2VzbM2tNDZ9ic8GpkqVSFqXxD7j53/ugmqzO5cNsmmXwVxXBNSZwrC0h9
fpZaXWHgg/j9TaYCAXTrNA6QrnWT9zt+8v55motJJAdYmWuqjVUeyGp0rfHFMMzG
+IZiAXZ02Uxiliom4zpAGqpTA+WPcibQyHABFZ5EAv7wMIWHldwVIWIzzRwjN/sf
vLSaI6SfGjxGHDRmVCmjG91y4sIDmd6yHdWSLUwMvRVi+s3w/0mxxNF+wIwlbOjP
RQuDfuS93U6Ho7kfjNfRmCCce5oaxJ6C1+Ucw52OQty02nnZetmtUszgyHHkZYYe
awt4HTwN7Sg7WzwNeifCOU+FB1a5dU04vHk4wmhe/q/v4oQI+/UDbiPz9EgeLntt
eda3Cm/2vZ2xdqvIYhRk5nCw4K4V497Z23uf965gqpWYAzdD/qJExU9BCM8xLbKg
g8u0B7elK0/IXE2klYmWPZYD90SLsD8aIjTYhTVLPhMUU/ZTyhyB389TZvHcr/Fn
nbioJtas9m+jwEApQcbHXjZaH0ZZWByob1MSlu2Md8LOXvqYpRIQst2PGyV0Pdeu
kh/p0nXFJ/I591ZEyI5im/6lI6IFFatBXtLJSnGbioxjPAWXMFWqJWINrNJGju37
+L7emB7bcR4ddAyZoBqpfLSUVbwy7zqFlxZvRpGO3r/k0gPKJNnfHn3GjronVRc5
SBTRUESVSGUwA5E9W4q8VAKF5I/BJ1Lj15TLtEJMSNxkY4zPqla7+5dDKA66meRa
zTGDUtLZ9A8PtERpsrX+yK5hiAOEpotiZvmP9gCwQQZgxrtwNEdSqsvfif01svQ/
KW2yo04DLq+KH8NQe83BTgg8t+DPHQUC2PU5jCHE5a/Q4l7w0ImLEDTr8Oidm9Qg
bfvNs8Nptoy4j6LFiQZ4i/70QpXUCMIXf6UKZJzZ+w5FWsSMfCDM2y/1XERh6FMj
ae+LALO9ynN6Vbjeashho6jIPTaUBEehDyqpi04C0ZrGYApT3hc/IWjpCXlb65kf
Xy7nSZ81myEg5G2iScrLdzAuVLBREX9o/SiXwncvdyzUgKVgljcnKQ3/s+2nLq8O
7nhQye7zOsw/fnGkhtWaq7qSeKqoxQAvqi6BbrruoQlLsSJwVesRyjB6tQVeC0Sw
87AW0aEK+YuRi0g2NooaXQBc6f2ojOw/O7RdqU4xLtb8n96d7nUUZ66dqS8klYLb
GNmTpdKovBORwxjXnMXwUEeYFdUn9dp7svu1hqCuy21KWGl7NqTzU6NeWSI1JUW8
SG0kBUOAigx6TnCoPX7ulm+upEJfl087rhglkz/EUBQSgH16bE+v2JnBaHZDPweJ
2XwhbReHIacoAyCa4emKB8U0xtmjEP4fGBLYECLS3zTvij5vBp1kQYTotGLxWXFo
N9BCQQKfPykzHjQ52nlAHVKJmkZXC/6zizBOaOcnbXwGd1yV/ccn9TRmXRGLqLyi
kvOU1rnY7Gl/mGVret8LM5XpranRbMRGSTYF/z1exWk3SgsmMg/LbycC0oqTQ0GG
dEfIcSK+kYE6XS27b5QHP4YLfgm09PD1Mz/L7QlknTGB12S0m5hCB71R2rJaPCXm
RCDBERclHoeW6EQCJOteS0U4k65RAtddXkqwzQ+G+aP/PzuSctx9T84YP3bqG/D5
EuF6NcGRON+y6QU8qY7l0EDeRXwxEbUtVKRKw+KU50Lt238fWZ9LYP/w9UXDjwoA
GrHWLbAFF98u6kr4AWzI3Cy9jz6pLR4L5hCjEZ7S3K4j4JXa8VArp5AMEcTcGq/y
vV1ShGyw5vS+fAADzYefBougCegCDLoPUJU/QCBVLdCGRFFyXCswbRi1n3AxkBEo
afFtvp/d8rB1/ts0sRGVZEXh82Ouc+SzaWky4v5qthkPAq2bfcbJI1v8XhKHgU25
9IyiV2jmnAWdJsQFlkdhx+HlBQI/JELUwbiUncJwiKV5tWgk32LDJ3oRAkEG/XNQ
A8HtNJGkMRqTSeUZew6aD22/vrC9yevJrfh/kDxSxDFlZI86fiz8FCkN6FsZGWX0
DvCDiuxy1JgWrXHLQGIHO58qX6xlHve/RkRUALhmyHNFg/4Jgi2UL5u/YVXGI37i
x1Bwvo0Fv1lC3RdrfCcDpXgf3BFswWlWboE++ZhzatJyf5azQ+/E45mynRAlsCvO
eOqk0QIt4hiuwrWQp0Vfpox1h7C3kLQpsxCwji2SrewskN0OA4PW7Zt8GjkI0/IL
QeeFU5J+cfXC5ovvXUex1Q2SOqR2T3t8+gG3iL1VhVayakFbIW979OJlKg39JX6f
ktXvJr8X7XJW8YD532dDPtDg2oiPLY9PSwyRCeP/E0zUX98E2kMeWBItKbFRBeJi
ggvVqFs8o17B4BY2wN4USJ/Sppo8H9rdkhNFinNKMegLbI5saoYZaO06GkBrvCM0
MoxaTxJBOPZb4Nbht6GObEKUUu84zxx/1tQRUTfS/mP31fcC7pOwSNIVWslYjTna
np1P+pEix3tMahOyikFlzYeML8axZM45tSAuHqbM8TrpAiffmdQ+8I1L33L5wqrB
BVoLBPqde23t+m7nt6ef0vpfLgkx6j6qtfLhyoc2woQYCa3BbBfxtgYj+NDEXNfI
Y8SPLsBDdQ7V5DQOw6Wlu7ALkv5wNr9UTqo5cs3iAUhnt+1v8sYo7gFeYTFl5Qqe
75dX82M2qxnjX58QJBrYFhnFDRc8i8gDQ+Ns2bRPU8DuVY6VNSxVfduSuPzoTEMR
IqvftAqyciSw76HPb7Pp6GsWaF7/pGUXym/stoLVFGkmpgR1mhaAw8F1Wzn8qWTP
bieTvuITX6NWHso/LTrVsRlsbwD/Nx9UG12Tk2+GrVuTYFZL8ohiHMuXBwNWNNR0
30y8dhUZwWAocUg1fr+A12B2pIkNf2t/1mpWw5wFBqW0UQpeb3/QHiMH2HQiQwEj
I035SSL/C5WFnhkuyK7ZNtODfZ50Nvan2TW5Vp2XM3ni4jvhs2xLxOS0pQnbTyQu
35oQa96V9e1cHMvefpurRWsIBErEBI62agfDgI0X8+e7gZHy0TMkJR65AahsUqVp
7enwmzOPCoTcgDfH25yI3s4BMv2vTlmihlGhSod7NcQ8yYRsTzT6Gh3GGG2Ezm71
xYlk1O1CFCKaPQETpd1J03+A7iHupowRMtOX2r4azXPZ0tx2RD2iQE3JoQvSHK8y
ON45a6s2xeJvAXsrU0CiaefvAxGnT5uOBiONWskTlNCumgVPM/LqvFw5QOfhkq5d
wV+fsOG7BsY4aenPgo43StF1Ku1g4xZGCnO45dqSYSP13Gjnle4RWllbtdfniwz0
CoUEiKyRKnCsHSr2mT5bcGnYxgB2pOAC8UkvYcfvGjIF82XsHowGCFn1UJmBCbrT
Orsy+2Qf40r9wkJ5u2FqJY799dbh0N67cjMIxln/J1ENpqql1w0ojlvxZAhorG5c
v2S44QE5VHvBoxMuGJc+3iOfZX6s/IoRPIHYh+NxJCWopTJpf+DTQIL0sO/+e1Ej
3WJarGGxgocb4id41caXCFq/YpxKM15Iv5iNuehrkOMFL15XpsQZ64ji8Ql4KGCD
uFPMZkxta5R+cwGEEqjaSBTD5X5PMe5n+gX87LVqHZCwt0JtCw5LCxJByeDgcDb8
W5lyo/Jrs1KkEU9jVLlMy+qv0z83FZi+jemA4Nwr2VlvNeSIO4V3VrPCpgDE46TE
+n8Ew9GBrbw6Ynre0w4k0Y1JpxAAobE7birKqqBGJDP856cZ+f467Jk98HfC0PbW
Hkjla52k/mfgM00PlXYCAbR/jvgd2MQ8yvo/8uyVYeH7Ukm2EM4o99kuo502utA0
I2HvolSqfe0TwW8hfe0EXY2KUKDw/w6IF0HiEQc+f8qraVzBgrgyxWBQUAkhO9oQ
nogwUuclZJWRZ04iSvDVB4DuCEhQ7lvuxqhuJBeAqusBRp1tLJvqWJHbMLY5+rVA
yhaaWBR4wjrMdidhfUgukwQbh7hoHxjx/OExW/ofCsdP+/t/ZUxapB4I2umIS9vU
kO2Z0+0FsrvBEoKzz62aNdt8TbpFQjWq2T5SZP77DMMaE4BI9kZMR496sbrd5hEL
wtwgX2yhA9ht2xfyseb0hS78hTm0GaeWJjelElotfd6Y78NaB2DfOm0AcOPz7f3/
jBZzIaVIyE03RSsWjFbBSlHVQc+gj3tp2YFy94tmX8UWDJlTspw6ZK8mvG7ZbqF6
KX2Q5+fTTvCmka4TbZbsd47DZQWJG5H14qpwlQuojdr0ITqZWEaEBGLYjUfmN4do
p6BCS3lO2zWih95c9wbuYUWgLNWgTp7PuG8EHU4vElpbe2cq6uNc2X7EfINCZ6+z
T9HUZPdlJj3QCJKIjlc3xTvjgV3wU2Ax4fy84gzouOcOvHxhhfQeRiCG41vnkb72
grMtUrngqKYHa0GmtsOPcSHQI2K76BgTW+XpEAW/TZ37O0yCEQxbMvWcJWXZ5hK1
k8twCejDD+y2Au7tF/zGlA8dXVqVoyuNidhxabp5gMqamcc3LFNpf7asZZqVux+E
fz6Ee+AD5yMgBrPMMx3nuTG+R/5ph1aTH8qyhVTJxnPO5E1LP/58Gc1GDl8m6TWd
Rn1C4I9Oj0B5EXognzY6yJdoDhWg18Odn9+s0R8qySCo2cW+WsgOEPtIYqSHhn4E
lGmsIuOxhkufJ9z+UHjloKwP2Hx1wLS+//Lr3SULPQR6gKhj2nK7JQ3CMMi6qUy4
/vPY/TaBLbyKdONUXmFAhNNPPE1kXI1Ig+tzZh4b32ECAMWhcopT68ZnJK6nj4nC
znkesKPkhlnjHvy3Lo+uvscYnA4a3uK1vtFgzH2OXpyoNJEJ/c376hTuuOCN6TMZ
PJQb2zgI6GNWNYmJpTPaRzLT/Lf/0XG/DbSV+3b5Xt3jAwkHTZZGKn3s14D19BKP
7f8wMl1N6gAebhLrvRtysQsgax0rYg9GPjTsUqi/n0RDt0mLREbhb4ZH1RZ2Pfy2
Y2XeF8J/7N0/Wv/4mlY9fA8P4eCSbCH0MnqZdJC6bb5ZMopKNES32wnuZhCNdlpK
ERWEXS/1nuygCnqZZJ/ApW109mI83/b15qDmNSeOFi/w2xLH1KMgRhkCv8szs5+R
crPYUgg6n/ra0lqFnzfqW88NtXu6WIry+Ek6VkxgEXExjnOXsMuu4JPTiW+RV0X5
huaoegJ/peNoLfD8nL8Pd/kHdppV6btsU/X78uLwkZyiQbCEMLorpON32ltEM+Nz
JvivMeqq9NPOriC4UcpxZ5h05o9SUtKHISfgUBfhMsGKa/9DR41gZmZMqoKJLVMm
k0zBQOwJMe+p0USpFvhZjIsYAARuU47NJVNN1f9X5qktmERI3PtLEYAtV/1j8FkT
M95RGGmJnwGc2tz26e5F/cpiZhbAjXwFagQYuKYpFnvGSXuLr/eCTuGx4wbE9LBs
6sUerzl9Q/3O90yDAxdFNIEzwIay75w81cZv43DJAEy4n9d4AHm22ExYRn/RdecW
RvUIPtJoOV9VcYpp/5P6KvoCCjwsDJprG0i+HdorGqtVgNpi1CUlOS/Y8yE4ia7N
iB3EMZ4i46T3oKF9FtKpgbJeHSZnum3fnL1bxL61jKOS0WB2hufUxLcWuObiVOrw
QVsGUHTHJhEiR5V/011i4PNz60z31M5sOm8n6hNYtC2J4v/Ww6NLr3OWnrVNNXrO
cHCjrW3JU8KO/TN9imjB+1e+B4HJCz2NGGxwA1/gTuuEJgDS04kyns5vpt70XqDn
MlX/4Q3Uhu2qBTO/fMJbYytP6MDoo9yslpSqGmohkVulCJEPzEbt7cSl3CXFxUNE
jJtWd7Q/E63AYgXHA9Xvo1WvK4/cx2VlpJpbFXmIz4MtND/0lzz6XgpurxwlbQc8
ToqQibVtAkXhEAj9MPJLpiQRF2StgLzZ8Srle2h9x52jJTuTiUkUTmcJAF7QTxGI
uWNVBXndHkbCZdWhSbJe2yID890XFe8bYDmy9UBDMOTIdfPhZWyfbFn9gNMmn5H5
dXpLLWEqCEi7RGRRMvd9333VFOEWz4sHXk59Bqgl0O9RAS9TJ/rh6Bv6GfsFCZIk
1IQPqXmQrYN5SjfIgXer+8H7WI1nwpFOfLmsveFfkjvY6hvNCs9k3zKlXkvz6Avw
C6BqOuIg8QTESN2ojVNs12E63M3oa5fznmMYTnIht3NGfUz4wg5yXWeQje8yOd5k
mRRuqdtg8jMCk6fSheTSc36w8J11J2Kxe6kSwoxYvAAocoHNefX1s9n+B4g3s4wN
hRYlTfHrKqu8r3UN6giSyeq/lOnsEi8tuB7ZG0Ky82X6fGb/lj47/8mJkZdU1AEZ
cBQF+eYo2TH1ioiU6RPIjV9CD4KRK9l3Jd5FVlm0N5s4ziu+Gg1qdy4812qZni8q
fdQelXribtn3QfyVFJHfQcLD72NB4yipwbTVrWssRnwZEfOgmuofAPHgkov4Ut+Y
jh/pWhRbUlHFEEfRnjqA2JlWHVdm9Hm4YfMoQ9tiU0HYKqx4UshnJwSlw0NwDaIF
zWzDHGMBgQXLn2S3+mjY2CvBYNaVFp7aDwjdwkG/5Q7YaSwgxQH7w1lftJAqS7zo
QqqefKb7er2iFxwoKVMH83wEu8/ISdr5AMbUZ/SuMQOrxbnHJxWjxYk842XmAlgI
CkPmaUhzulmCf7L8UnskTIrMiG9UBUyTItGWJ1MwXoP7W7eZrvzN9sSEQSiw8l3/
2XIoA10is5R8fQ0reDht6MCpTF6gT4mkARSMJAxt2EH9zQyac/MtEStZNiWegeMt
o+MyMHIjLIp3weUpIAppxEWuyJeTclVCi7UcplTQQx97fEgTBLlRkIn4ri2DY6xs
AnVeRNzZMdlv1jWgaj7qE0k+8j1oLVIqkb90si7AAt8NIjljnNpYZpQF9mk9Ts+k
FkHJHPmOf7NzqXtzJfrTquZUsgjgpZAbSaSoo0gjSp220lyckVprJ9DtlFyPnruI
BWW7xVdx+FnFO/YTAfxYOgNsDr7yYrQknE5zYIlyQEO0RrsVMJ/RAP2WiU8N3iY3
y6hm7u74xqwYRbbqGOffA6IhBxVysz/3X9jJxi9XkMv+pUng2yhN8WbgfJYBHBpm
9PEo01fIs2w4qM2BUX/zbLliPwkCV6hz2qXRHhUJNBWPyZfJxnt9nsP0+tOMbW5k
xDvhXQYb+I0jQ4C8ht++7LGur+AFGw7tb+12xgXbTtfptda4sj98HT7elq7IBCSY
zCctOuP+xBi7uuIxGzFVFpCbQZ9pMsQprCDOnS7/xFg6bIsBu2Vk3sgdQa8KJ/qN
oWDS/cT6Gs/jyspQ6WCM5iogPJARBEJmRW0x6ZEfSl5sMJprICiQ0sTrLxeDMw7k
UKVMMrH+YHCmRprRU8oFy7DJiPfmtRkTL/mVdG6HX+I2MLkKRx412yGbtQ2BwgeQ
oAJ8z+wEccuSs1kVCxNxhR1ulrWex84f6ZQRqoagsLVq75Vceyl3LG9JzlTvWzB+
V9AlOk7mvtZWQvGfM7lKQNxAe6h3WYEpWbDBNLi4IcCHC2lN0PKaUORYsoc18JL8
6ENlHiik+9B4YagGc94bW8iPdbIXt4E9wzQ7RFBv+M0uhOayBDgCenAMfFD81MlM
hWIpli9mLba646xlpQf6KXZ76DPFJkMVhulNf7ze9qCfc6kVxIRNwbVdnGiz7Kru
REPOLSyU9mhzVITQA65l/5Ut4ylhzkgJDmZbEMONMpg56NoX6U+KJGYhcNs45d4+
URKqPKKWsGu5OKtH7zZgvbBvQdzOZxkIsd3Ahf1i2KzMdqE852W8aWmjhSPquhFw
HfozVERjqMVv9jG/ycUVawtkklD7eYDt4lK9Th1USsqxongEyV0EgDPNltwr1Di7
LZOQ62FKCY+kBs/TePF/PAukhhfGb0UxWoVSIYANTXPMsnJp0OasoNdNB8q02kJo
tnfs4CAL9W5RE2seQeAB2OXZfCB9tB2d+saULZkoAaQk7/qg++oQxztWhY/qraqJ
OY/SIaHUPPs8KfabCW5U8j7Zdiulrp9e6xwLvXb9PzkT84Z8ztTHSRR/9Ys8uP9y
+s9wuHwBWDJ/Y+GTQjg0IoZFOllcdoqq4B1VPGwZYipJSRBU00f5hNjTjOvxSyjz
cO09lG7h2wL0lHPx8xXcPz3edRe728ncXZWO2xQnDxKTF1llL96BA8cfL0wJUSjm
+JJWiOOUgAwQPSbJ/MJUhKnAguVVuSWhG6Lbx9B29w+oZh68p3ySDmA066t5SPSl
gOM6GuQoCC7QIxd0TnAPvSZE7w/yH3DolRiwYBVcnWiViRwNwryRn33l1YTZX8pv
Z8RmRqnvlhnTmyNo5qD3Iw1/Uljxb+M3V84cB4BEtFngHUK9gLtaFYoSIUcb6jy0
7UuSSbRp45bzSHZUB6hs0R0XhPf+70OYYmFaDX97yx9QFtDesQ8Zml8Lkc40rL7Y
YVMlMV1w3wFkXA5N/wpnb0f+pOqrz850cUvYKwfIzWDxVAWUj0VBaA/tJgBKEmLZ
hEpHc6GsbqQam42kmuaZ4iyMU/ZXdwBbAP/oZMPKurjj8JwqmduAkZVOJX3klzX/
PCssBcsLKfKxzvpgDkFsaoNQWoewANgq6X7As37mp5YnJwcwvx0xMBzsDq9Kj/3M
ZnOUL8QuoIszBVZYXMoLTGDof6xsaZsDRcafBXVe5sQKGTc49mVx2BqVjbvEDJdB
Vf4Pbg0pNe9EC0z0lGv/y6onGha+M9HMsjJDQAjpkAQiE3w01c1qnHepUBwDo4EP
f6hD8XmvPnth0svpTRAil5W98iGOdVdAvnS3qcgCMm9kgxLo4I4pFRBrPAotCgzM
2awJp2yIcckbRpXLNRq9Ux4cZxc+874P5UKuGw1L+kQMspOKWZ7GEgVWl4pc+ZtJ
K2oF1wNqnthY4VukJ7VnOApiqMcgqEGRt9UH6TpcIJFQrWoUzoiN7lL8zXZcRoNZ
RgitVxg2VUBLCj3V3VOXylpJxS5UmeWzFJY7X6uLzl1YtSw7hP7haeYzDTPK6yA2
D81V24784Ry8/hIUbMDcfHgF547y3UIm2T9jli8a8uW2sQNZo+DS4rldMK1v3ulT
yoKUUbySB66ImxIATYSl1xiSgV09YY8305oBRIWNhIMFzvow+iB7DWjYM8csmnk5
lAvPgi8CjGvhVELAKanwlPy0f9eY5cZ5GYBUu7fbXO2X4AzvesQB45X2t56cSY0D
28LbkoxJDAdTWWNqa+/w55b7kMibuVL0BBEDu1W8tCQsKV1GU1lDs/CYAou37XaG
uzB7Qp8jYAzIbFTuaWvBtxYzWUDb4rksQGL59VKOpjX/33OOYVgrllER6XggifZU
x5teuuYwIvDu/D2G9f6liGMWNydcdj8sq2ezbh4eC7Ke1/1bL0NbXSqxtdcaxdt9
KwwTAwI8eBhmEXIth9uSQogHEfqmfyPXZcP0TyYD1OJB/3PLQnf6nYR9PGa5pyLu
wzyNgI8rfmKz/lIb65M6y6uzUxsdCHJxJ47c0brf6sDhZw/VCMixRw3V4Y0HCyCl
2Pgmle1uGrs/cXMKdPpnG7yRj59Ld732EvVkNydgGQcvuQLVntipVuH6vrUMzlCU
O8/s9I0bKuRM6i9HWjB1+HKg39a0AT2ueptrbpk7f6xLv9stJUnG5BGNBPYDOSuQ
jisDT/ILshzI31rMTzdZ6mpDYjYCdOBBt622x4m5JdyCLmexd592xmMkQsxTqXMw
K55BpPRZLJHBUuU4Lp7A/yjTUKJc/uHiDm3KknKEwIolFSOz75v19JnAF/BBj2uV
ODOw8r6CDgtGrBUDO13FiyH8fCcbm+wuHiB5THuJASQ8buhFJIp2c4cYFa8IPNSr
jpl7rWbw0lWN87/WPFExJD9yNvhK+FqT5inXra8stlKzc54QDiz58zSgKLik9rVW
ei7wEVxWLPagd6WpRGxTYZTLp8IRzRT+heKF2GidqcF9epIsOs+mbLP3PXMMuEIo
1pS5api1aoUoWylZAd9MqCzprApQts+Yp27d9oOyi3B/OO6fdKo2g96BcR/gAJLm
eUfskfpqrVOqr0cw1pasug966u0U847jWDPZvG9Yqg8HohzQW6Ew8kmf1fmtOx+E
MswRGWMIslyq+jiV5oqtpb6zuwy/ehP6whXtiCheuU7Up/1pMzE+6TOUERGTOL5g
MCI+S3EwOt+arNRVxvW5ZDJEPr8JsT8NV8mQF4m5pjICYRytNw+o3/gdIGCWcfcx
Iv6rA1cXak3A3pkhi3TOCyjJvTdeB92QM7cpuqy7Senk+IqhBcxB6FCS13MpuuX0
b8nzt0glvQzCo3DBLjXdx79nc4/dfSLkPiJ/cwZ6ReZk62dCxLqlMwaUgOuTByPg
eQfVeySDjB6nes6eWXkHZv8hGRGxF2C6SvEyPapxd7X4mndwpyKd46MaaBsoPa5g
NLEsQf1jxpnih4boV/AjZwII2BPj9VWhgfHm5QXTHEcbhwu7pBoydZ27B7rLJhTp
2puSNZmCHVAa4edwn+3NyzIrVron8r+0aMxVQ5PaBRLviYEj/dx33COeMvt2SsTT
swh1fn9At8Yduc1sMAXvj0jKVJzRMoaPxGRqpNrosA+F1FGhJXqyYqKC5aA8/pfk
0JwDJDRlKpuEV9alnPwne1joHuGy5A6FUAiMv56b4ap7V/yv/cwJYXwsHDNOqfUJ
lHX6BuMFAIrFbh4TAyoRLc+V0L3IY39/0bT46Fq7nFSGs+/hE1ahZ0GQaVZRWQDS
nPmtb7/wMnvWNVtr6zkufvwO3jICwKvRAJ3+JyGrvb1wirdJLVpukK2L+LcMdqip
1wDUn17PrpmOhjTkl39YT93+LQsyvi9V9Bn7osPCh1odXn6zn7aTW+sOLNTKJT6H
3DuDOu5Ph/mb1E+wbKYuvVCPWBqUd2N5t8d/F2oZo7wN5a3xoT+sukaflejt3v5O
Fz+JR5q6oLWAhnXGqn8yON+TdtyipnYXy2/dKjDRnac5y4+rV0HC5mWsUZBPcoBu
ON1bNZB1fciyiloq/C3XzzTSpU5GYy04YaeoR+vAnAvQazK9TRwZ35qMGtET8FK4
bvL6wDzNAMBNSPipvrgjiarZ7Al1h4WQ1U68oOfENlznVlE5V+srMwQqcrR0ONNw
0BwwBPnE641cKS2AlXfUGpyJoBb3mJSvIGdh61bbIGARXOhWaQSS1JqAOLMcnNKn
scjGE3JU5iCDZ66HxclXHOPELe7IJnbJEyZMM7YX2Y/4dlGE8rYQZeJaZOj4J02Z
+uz6/0mtU7u3XGy+zngR7iQ/h64gS9+0nKiA2b3gYSznxqC11hHa+hbD93T5Fp2Q
J7N8em5taOKTDwmUv4uBpHqrwUMtLKYWJUlyQziR1Vue2bXQdAlI3/SUM3abHhst
jE+63eL7DoY+llCIEHFJt0lsMKVD3Z+/d4gkOQZ3z0xsLFCYdqzHFwq77fU2Mh7e
g3yQUoQ8FzdArlHZ+V5CbXxhk6M2bfQYq7e90V8d+1FgeKxH9gOCRL7nxMY3wDga
E7nwTknP4UyzksLGmKA3IarFmPJ6g9z4weQfZ6c1s7HWvRIh3LQW6d4JRwwaz/a9
0l2HvLrSY01w50UEQY8vXtjs3lIALdBOFpd+0M9MmyfQIyHZwgCp2vRc/Qi/h4Vm
ZmXq+G74LfMxwDPd9lZrfEc/RSBVsVOrHt1k1L0zPlKCuUSrWBJMNDbYxsmpkGOd
hIFGjfsyt6eC/QHWGxEY1yKQ96/bLEAUqC005us5iGjorouXNWT4Kz3ziCL3f+lZ
m4u7enow/AFflW1/devJAy/vWz5Lac1rNyzHM2l/G9noO389n0lMOYdSjcCjdVjW
QFxw5ShpSqRtl6RYs6JfXcTiiyFWVEWO04gG2dMTUafAMV3X1yz3W6GEkWj0R3O0
Ps1hXEosx9mCaeZSjG0hLSRC0hy72CPkZ0l7Rwf7+G3YejrFfAQA0l2v6V3b5El9
LIG8N3gPC2I5jKdxRYJS7i1G7aJVh6n3oHb9gL31HoZY8OzFNo2XtaLfwUvpSfVi
3D/WHIPng26InOB+TjUM44l/XdWSF8IMxFQ5iuiA+pzUseVXWY+3hVjzp6VWVxiw
xprFB2twhXIRlIRqSFR8SM7Yls1LpuMp3Di/pH+rgKU7nvHgXqq9ZRvGB8esdVng
maH39CPAl+lbdqZrVC4cBBaz/G+UOpHLMvvt1rrv1Z2AcXxIaurJZCJ7kEyLVR2K
Gm1OcRXjoYoggyDqd6JTz/LA736ksWBUnC/RJLc1MWVzCkmH45BOKltVHOJkw9Ar
gB5KA1gLin+Xs1h6AGIIhKklna9YZszbUfX4GWmeG5QjddL+ntenaH1s+pqGJ1zc
TaVtqbK30krCQXJx4BRwuJuvbXfz29r4xhVh4IqfHuYddAu6AqRwxH0YS6w/MeAT
h3mkle68AKjr/jDYMphy3tb7EJsi7ebjMeucCmLtz3FLCHRc/6HlKykprTru98ZB
VEZDTnFcNX31Gg6a5bReKmg/3qm+XyTlcXc3JDjwoEtAPvC7BoTDOX/XvLT+gj65
mQ1xLbJBkfZIeBzOSvdaqfv+h6C6pVCE4mZzgkdWlOx+swGAV4JqHkI2J162/rUu
h5Y2LnieBZdKu30Uiy+eex9ne9aX/msi+P1/cRAnw8KeLizIaJbg/LDAOYrbX+8N
SbVWcvV/fU5K1tVJz8UK/HBnAuYxgtTwNBdtBEGl7CskhRDCwIgatGFR0U9NDB3u
PSj0ijMCWwHzbWtcl4RD16YX0SbEOpOH38aGBVSuUCo+1tJfgJnC4WdU6GQmjFNi
t/rzOLvm51+OPjS5S+MVpGevS0Zh94hLyMk3x509Bce9y0nA3kd1gvQgsmeIUIws
SGjnVI/StyObxRz5KnLbfX7grRL/LgzCaYcHuphHWUpAbwGI6n7xG24DFpzULfPb
5qnF2Hn6LcOkfkYcYkEdOAuoa1A7euAnR6k2WxAO0e05mFgYoN6GLj1DECq/DCFE
W7qfdYuHrU+kLSnJvlj+qE9ezeUxyzprFm1l3qQmTcreQccXOMuvsspRInokM+Q8
ld06avdowLNoUeYhEAMZn67vhD3kyuoHyEhUjNuVwCjoz5qk62kWOxtrgAkzryWk
vuaGIco9AXtbRNxw47m4iqYr1v38d04fCF4FcO+gwSl/Op/U4MVG68Uaz9zsljBI
YjYJTWMvJ5Iw9WNI6RwTSJkrieJ/VF6GIzv/+yOLAcyFYHKc8wK0CrdOh7ZM+qxn
Ee0y0UFfigvdvpqZIde0IT+A6Lj/q2ouLpHmuuC7Gf4gY37b3Q9t5oEI9AgJnWs+
nP5vnxHWXMN5RCwtvXSMXORSdsRbqRAMghW7FVMqHKIVC9r29tFsG8F8ywxl0eKY
Ceb72FfaJiSrJIDRspE17bwcv+S1kQ/cSM6bZ38f8jflNE9N3JA2UEr7scsoSuob
QkNypmE7IO+Yg+ePZO4w1Jo+KLK5rfX9LXyus19XsnvQmOHVPiCvDDEAmIBzW7rM
TGTBtJY9u1b2MgUh+tOywbOtzzZdf24fdsRbMqVZcBck2kNKgV1/margZZT/k9Gy
Krg+HI0w5a2rWr+gltZsva30F71MuvJK5ayip+VGEQN1wlHxRKsDO8kyicAFqCvj
hnJAN+rsXZzVPs7NvWVoge4xUrHyn38vVUyaDBZADWtsIQ6C3dZ8DclWq0bG1dPT
pEJD56YnDP0tANFrnM9Z0XQwBlCVPPcnW6y/s0f/2jHFW9nbCfxppVq+E4KFBksJ
lDJnYAK06CNWkDVxPVblHBFr/+JRznwGa5YD7oNbkwR69pwiww2eFSqoR0o8qyx7
dKIkWmv3KFttwShc4dnpw6A8TmSeHgkGBVwUWnvkHV1N5UminXzRV0AKVD/OyGFh
Vb6AHcumh+nq3BndRkQ9yDemFoW6XjgkwkbBWIQ2rgdx7JaQPOwLtyk5WirIlovd
U8hB5jV8JRfGQj9gz8VBnewNSLsdmfqrmF3c5PSiCSLsUyI/kBfQXjO/8XUV6vgG
2jlks4aKXSArrfKJx2a8K5aKms1V8AHzjs0QOJjU+GH2eXHK0ZpVNAbaLsp9InGK
oFyQeLU6dJMKmkMMB2a6wMLwWlaYBGu8M55nelVr4LN5v3XLnCSfAjjknF2ihBdy
1pQ3hTvv9jcWoVOxsGXRlK54JhhbyVuqAvbOSdhg0WCvvSnEnY4/J/dbbvf/gnv3
aEHYYYnYY44dbgpvz3kYovCliqClYQAuefq2x1YZ4JLfREEh+7vRKpCyzTgDz8SB
yh/NBL2jtjNNyYbadOpq+GM8MiFGPDqa5xNwjul2ZCbNkHEFF8GsDLIBY4J4DPMl
ay/cw9SwNd+VW0M/F3jFnd92f0aSTlfcJj0vD5SnIcOmP8uYbemfTZ0lZZLVOlaV
jjVwcGHQ9coLkw7xACC3EC2k6E65tR6bG3bDDcRbUkj6VdjE0RiIDWO+dFjabpVG
UE2SDUDdqPTn8/qGCV8XkQT+0DqtjWYeVPlZ2L7W/jmhsOQK5TuhURkqzUziKwjB
7ykfxErOIDox9yAEGqx3eMM/hXX20jcXXxYXiH+82e+aQTkeLVVFac3yovVdIa3Q
OHgvCob1MZJt3Gmp0I3KA4fIYhIN6YbGwnBRV5iTEtw12zFrjxDZto7xit7KcW9S
hwpItQ5ehbPuPBMwU/cMtLaFBOxIt5jpLJZDVtuy89/xKvGqJrYQAzkClP3mj1p/
DnBhzvkt/37rtdrqrpXGAfnf6QkHnieAYWNlL5yCp7e7pWaTmf1ZP321D+4q9437
WEbsE075BODnA7s2fMYHu1lPQUmaCxDwibkJ95IRdv5ZBchGamerP30pypJXFKjk
OnC6UXv1N7q1Rm5qfyhwknf0majNJ0fXMOdEhLhKHGNfcHfIDrduEoFIM2vOM2e3
wUer+JcNXoFKIv/FlzK822CdmchDWAiitFZ5zkdR2NfSULI//+ud4pii/w4xen2H
JpB+afhXnlcbH1IQLFovziA+9sJFeVglcoCmXddiuU9kVe64eL5DtG0IQAhLCR3k
aIjbufwj6RY62Ysjk1CJPlD6s823lq56CADtT4WzrIdZ7tRK/DT519+M+qsP2gqS
uQekyCQ/Gc+F40NgWjT4YMPCojmkqZKgrnwzBQyefw3cLoPlDsspuzLqatvdT8gL
ntqGXMLJdS2qJLw8K/UaaczgiDfDf+FwfAJtGbnj0ZA64HWB2JOgO0/4Qhlw7r3Z
f+VksUtA/n7ConFj0w8RqcjQRi9Ng4xdbbdgMkT5yO/rPwP7qMcZ7q2h81o6IuhC
V9BlyL152YM4F4zaX92pZ8kt4H53Y9/vwPKmQ47On3tYxwyPHTZ6RoPCVFR+AQ6F
UePq5wdU2nXMTV6vpb6B1NcYLotLHUSaOvVrLWYIkPbdVVtaP7PNezE5U+qQrHAF
o72Vv0HuvixeF0toayub90Y3w5OcOo4YOA+LagXBP6WQ8cV9oBclLOFcJWKDh+Ki
wiVmKsT3in/iZNpXI2lTXVTO31xvq2qaUMbk0Bib1914hlyqPhPBgq5AEx+Lo3BC
jL8WMJYesLW7PuhDCatNlyuKPKyKEr1dBKMh9BePTM05iqIQoRSkg4NhQr3sdo7V
uP/aq7PykGGAAVypk0V+qwhHvAiFF/GuUAK6m40XCYbBKp9m9qSoqjL2DrTZpxk0
FIB2v+7VNEvo19H1tTWP5CrKb2dQTli5KNRP0dXmmlnRiaPIjZU+D4qIxFhSruwZ
FCWTV3vhGtr33KdckJgxkkMoDYSIS4rQ290DWanhIjryHD0SNZLsmulvjMa5jNio
/r3TXljVXR/ZPP+A4prL2gj17my0DoHWk3rkQCgXTGIBe1p1WUAlbqEbgozzaWbK
MD7sTYRxvWWJ/mk0plfyCxIPLzKPhkQ496sY+HbbG/n7DS0C+KXSOLl6ec/uicZ/
UQ7qYAfx5GN1PmZHdsqTDpfp0oPWBVdrZkdEJXGj8kymxQW+ZVoD4uvpV1MS+H6e
xabelzefmVlx2zotBr0mMCAMf6t2J1MkbGOUVm0TaASzs66nYz4U0xw/wzt7hJp/
7AiiVx7Yny6m5elILMZq5NIBh8wC/6vMHqRdfIcG5kBtkIXsaqTE1FrAUVYPNdy+
7l7w4L33Hb7cFjvbI3kR2Sm0MNjznm8q62lgvgVHA9/84fwhbq3x8m3jVgWGnZ4O
HXQCmiS+YRkOnOjYZ5kaF++deUniyN56W6fniOabdIwx6vB6fvH/5SOwabkm1Ewd
aEu+LXcLobHmL6gKMA9EOGeEKmgTpR2EantuSKnCWyVKdNevcqZ1o3A304Paeb7y
ZMZ+a3IoEVgANN2C06j3JAywMGZJF1km2l49pe40fDtuuGGkPiDt7ylppuOd5vdy
Q53dpz7mqnbQWYoZ1wmrBrQmNdWfHN9L4AoxmA+7Npg9pU2SZdU1cYv7LUPjXszm
uxVSehsn9fBKbht+lJcQo6KrBdc2zMj9WJ2fbeoAQx169dgIHjkOFvhOrM7wKZeQ
zFtMwKbjwyrgGHHke/slytFL15UZo6Ufw0/4ziQhesdOcJxlfs8nPDMYYMUxRKKE
MZMB4lZ/V4vnYJXFDtoUFMg6TLgQi8E1NmJvqAWFcVQLzQ+XV/hMtSg0nesGNmEx
fAnrWrMis4ep6el+HdjQtCR3UJAY+LPgksIbIsp6o+6CFbVMf2+4vj43ynRqGB6g
o3T6brPSKHGbL7O86mtJshpgvuyczDQEwiCFv0Re7sxK+DTv+oF6a+y1y6j0ZE/t
GZX7e9yR8Rbp7I8TCGqPcIECy9QqhBkhDVtMKsHj4v+1hvNlHw1gfEWRS+HOHhgF
72Y/AUpkTC7ttAo/uVO35ND8EuQzH5be/GLW89lJ/XF0s3oAt4RYPxd5iVWsEq1l
kfGzsKUX9r4iQQYMPo3Mm8JXrvpejVx6eWsc89O9aPbMHH07MN3SAkqSPUTrrAXn
XEueAqO1/jrAFrClUWtbFyHC1tIhubPeCdvN9tHtIBl9chBBcztsW+j7dRzRwCGc
UL8o9f9zwUveqRii+C3tYDL2xNsKjV65PJdQlqjjRc3zjF4uCPSXNHo+WkUfU+A5
IlcB/uR/C7iv4xxj4RnfYrNicF+f06FxWOm89HQDl7SlxLSPhf9zM11WhZKpM2OR
9vP/IDNhPbGo26mi4gZYflnS+60h9fSUWUJLQKFWgbquTR6PHefDjF5sOgJBjm2D
2r3BgXwREGDtuzU9LTIjfjxemWcRr/mD73dmlj0opuXZaOjFcqTRyE0ObeGPZA+b
pZQzDiWTHYoGiko1uXDt7SFj0aceU+MRGJP0cnImj0qYfS6wcDgpD7oj05AhqUkV
190GZTUCU3w4lrElApNpq5T0CANUfsn/Y9nXyTKJcLpsmE31nuUGBLEsk+7UfROn
Zwbn2oOEp+cIx2tWOoMrFg/4vwTYGUg2ybe0d3ezXHs5IuTd9gDjxXxzaFCXI2h/
1r3j7jZXwGDj4aQHns6kcVJbKom+92/Exwo6Qal8PqRBnuFnUNEmJK7zFTWdlUnA
J5hhE/OLsUlztiSjiK9jnlkDpLEs4YAt1wvtTmx+XDnMtjoFfVQ96aewHrSRgH6/
Dlwo5MPslJbAl80uvtipxzDbs/7Uh79p+ip456Bz8g0iB/QNpW7xP35f/EmMNkY9
2x5S5HCoOUtfBM7kTcQIIbfJVm7fyNVLZSYVYV0UfR9v8BrZfDM+BuSngRxUO6zm
W4BIbsW0zP0XoZ/N5O7o4BbH6pd/aBo+WspkpcxrSz8HE3S9QSrAbKD2GiKzRCZX
DJZ61z02bO2qvNdf4xVRiq2D3JdeXhlMh8a4s+BnvGvQ2d2WycRZ9HYhU+wiAUIN
RBz4VC0C74vOREulJKTU+1imEqL6MObH2qm2hsCQFYJavGDAgbiWjeMx2rGRlv29
XzF2mM7UzbriKlumVurI7ezV1ma4vd4W3vUg+nTddncfw1fau0i3HyKDwrdSKMZ3
zDvxjJhedQzE9tJfaDiK5SN/72HGnwW+CvdM4PjN1HGanzxnVi65oELGiZukOyiL
7BU6nHo4BiHiJQNWkeEcz42RxnAO70d5hNMK2xqRgTANVqhzsdAbboqR5hjvAsVe
rqPPJ/WobaKoCOLoQzIZ6Krg8qvVMGKsNdB4rJAO2WT9KEUD8kpC5jK6/Ni2omsJ
AifY6OAFr/KoWrqqMs6dZUWmnx1hsm2hg+22eD5+KC6ODkXFttysLo49zePWaU+G
hosooGuhMiVlqoESzyXY8bDVL7kHet7xY4pivYcOjerQpJojuDiX9pC6XSpqUebH
/oj+iJWMrYg/WO9IRK5vpS2ek5R4y7C/neY8SsYmO8Ne9MipR3V1Sh5e74N7mlgB
GiZyHgIeO4N2hO5hHzj9TvlivFOpkNlUElypjNO8R8hOXXwg7i5Wi2N/kTxAkfZT
vQwVmORh1WBKQSvEcIdqXfcfWNdtrTAeOtYTa596S2krEjcAxu63ehMSpC3L2hyP
2Fwk6OwWrIPk/cmA662l0hYqRTvhH3vjViaFwLoIzTB4Vl19YCuUval/y95Cz2c2
u/XTMJRKsDgUkJxAQzw4hDigaCVXYakG7oCn2c0GBz7lIU7dSOLY00S6se2BNfQ0
UTPB6+jBtvcAiTmCcXlOqwnGgTnLFuwhUfiAan6e3NwpAIXmVLmL6hEvu53NLhTU
ZMiC18eAsftYiUjov2a2ER7N66YbITo8uFF9/YpIolzyorChGT4ICRTe5K19RaaS
EiUXsmrlbZn1HO0sO7Qu2vqE/j+AUKWNpj3XN3GSRxADP+4dvu2uzNX6sSIjzg/V
vVj0iGGKdU1f946g7je2zHXOwr0Rmc58DRwcO2faRBAXQ3MXKSrLJvUXdkBwI4y4
JwZRDkWxkbTUqH+vIangYm1Uhfpej9My8QZeMqXeWEmhGPlMVAijeDHq0HWTiU8X
6WdSsL4Je3gDjTLg0jr2oqCSITuLB2B6bIpEen1XCH/YCzkxsiPAB/sNw6VVaOgO
yxdoICWHbAG1Nsbl+zL+7Dk33cwHMRzf03EYaKRclS1RnA39eUR55DMlI9pp4wnY
KvQWcAaCAT+p83w7JP9ldldVGe81dJRTy7bO2RaRhu+phiXyXT6raBbz6vbcQzJD
cv9LHq8DepXw5x2JuxGtobQ54XEq6VARxFHz5CEnUqex9C8hRJrZQGSvJkf1i3cN
MCY6e5rvFNLMPvV/zRuHa+BWGsUkT+3CCX1kE7PokdDajIIO3x9voknwfT52HI5+
wa+9GLz72eTbkgguKjfoU4RFLfvBT40x4WLFPObg9LfOsYGucIlJ8JgGGtLkg8Lk
h/pLKwRjUtJcCjFZLHMbKalHldbbE4nwyxOUQtWXfjdjY24icjrp/PUdOrLucC82
XHEMHWwaf/rRMA+P1d+ou7QyEPcLwUd3CvPslsZZwzOKK6CEwfo0eUt7cQurummn
jY+3iokUMvQx0P4rUMFhi84xH4ZgLBiWb6o5qVRADM0sCoGLdylyxzdjH7AA4UPJ
QnkQPwsnoFnCnngtDJXrNzSJZEVpxtMjT5OVriaXtdszEalVpqTsjq5yWTaYxaPn
NRqUrlNs1Jz2lWBMGlrP6O+zFLXPmJLL6OVDJsy/YRs+yzIxLS+vHKm7+J4FXwL0
m2ZlOziUOTsVpCCciwYin0ZJxG1lAbf2/BvJYieNpmOiRJ4IjnX+ji2amA8YiC2G
A/C9ah3xGL8qzVr5mhBXXkO6Ga4chDeY2Z2Yjayk/ywBCnTmkk43v5jvfDDzMjxf
ePa1WhZTp6j588J614Q2av5baanYDWEReqqinhsZgvOE/UIkslY2i2oR6zjH5IhU
vYzpS5KwIdoyPdaNYFDCrpM0jokKwaXntieADmHdU83IiIwA5zWmzRIpkLpUtyh5
9SzYf1vqNwyexdiYG0kzHhlVC/JXkXqs0+u1RT6tVgttettN1zdl6wLUbCAmmRcT
HM3GfZj0VJIjEag/tW/UYBR4L7D1EXJvXh44O1iD4VYssZoqlXR0T5ea9KLD09bl
pVlJC/WJxbwhGlOtI+Nu6kfeseYerhKYI7OpmOuSWlDNHw3KBjUFQ2OHRTgnlagt
lEN4dF+SXX9Cp79aOciAzYspAsCLAb304aU78nk/cKdpkbdwgIgUadBchPU3flTG
PnUnRKH4CM4VMKmuGthcvI7gtIkCPDQFq3f2ucSMa3kUKAsH9WIWpO/xAmISLZ3Q
+A2F2Bv2iWHIRyZ1N2c+Lw/u+sIzxCXs/dTgSGA7jaKot+qpDsOFFpj15ZbiNtp+
Z6a/D1XuF/sdqaw8RFY5v13W7XIjWTAzGD3qhqzkr9ghbI8d9TuYZ4/yPM9WG+kJ
pnILmX5pPIIa1V9Ov0fMqQ3Wi2UCMUFo0Vmz4FeM3Gjt5rs5Z84SanZHrQjo/EFP
t1+793R9fn4IgT+ixttNNxIwG6aCBVpIUtyAgJCsmr5JoDE76un3Y1rOdxNF3APQ
/9zCqPNuw2s0vEd8lZAfPc2aSOOy4YgjSSMXT6jHWSExtTo/lFGR1n7u0m1Gk0xJ
iKIzNiDf+exF+2gpLJsJudjFvB1D3Du33tKBlTZJA5c4MlkVIGRuHZyTUvWfoRpy
Ghfbfs63wYrZv3QIzpmSt7JHIv/gK+qjbAcoJnYmTY3mQdRHA4eVbWGMUWNCjRqm
Lw0+Im7HfI79L4cFSKvVDZV5bubw9H2QE92Rx7mVzlbtwjej4ngzsxssKIdcza25
235G3A5MumIwZkmai4e1Ot0leRcZOiDeSzTjFQMRc+ombvg1OAm9+z81X4qFv84d
N+CwMvmzH3r3MnGYt+Vg/8kvr94rlAOsha3W7fN8GFFS9M92/qYqpeQ3VT2Vjrlu
TsW2tb+dy5CuaoFBed5B5tV//xGiwo3IUpyVfzWiooFkxwsIJfkfomGFlCLQ29M+
hCRudoSRqIiJvru//gSGMgc3ys9Y96yvDstyu+Ukj3NVsl+FnlyjOiX1dYZgr9yx
sxJmrui+T1FSyUEeVKUnqjywzg8Ci3NchP/wlf1CgmMrbs0Xs04eVxJjk/WaK7Er
vi2r9bcXCrHoXm21vrifW4LKXGfpbmO6SG7BViHXiobCPfkNkMbkHiZZmbrKk0N9
jkXR6gQGxKqKvr/QcJZX5w4Cu86i8ORSuOqWUL4Ixe2T6bOTi6g1l3P0ORwkEVAE
jsIq5hF/j9dtblSR1WdLuifGGQQEqd0OE00FfGFWwejzVGvm4Bal03RAF8EtvpmN
a03PglnHQUi9tUgZKZ74BizLVg+xFkacY6bWrb0AMdn1y9u29J0maSNUl2azt7nR
7Ay8wdI8ngT5tYEg4K/QOB6eTUvrZ0qfjOPFbIWFNBimgozIPL7x3GtTW71Ab602
0x3A8wVRQpdmgxqd5PuTTS1KDHEEf5pzmBrptkbmtE0Si7fEu50yaB2JRiVmQEqY
MqHnnvn7vcapUheYxFpx89bTLMxDgBAU44KeS5nJB6ptl94O+1vblm2DHL8zI1yA
6kMYBTGEy483ZCuDvHi+5+QmrQT0APteljtbUtkpKVL/aidjf4brHl4Q3rPTwmbR
v8Pez4m06uTGIUbmShnJigqBjls8LMprnINXnRBa4Rrl2HYMMT3zMynKLI7klz9X
zD+SvI/cufpYc3wv8D0p1FUzXp2RJCwRapnLDIGjwe1KTV26DY7UXrJIl7fGXV5v
FChl5g9gOL8TraYeFU7/hMR/tOKkJTqagk3eOLVRU46cIiAQnhnxL9+vW8tdb7vb
3ZK76+7j6moF4cVkmIia6M6kz/6n5jyT78XbXW4gEeFJHWsQtFHFI0uCaPWxs5TN
fuaZ3dA1iqBYX/6bkK13iRgc482b4PCE2dimRCJrMlg+RNo3mAWADtw1Tj+a5Ssx
e7+l7+4jJhuNME8e6MW8R4BpMyL4NaKMU8O0NCvLjLFrsIProY3bKkiHG+JZjxsO
SG1VmCFfjDDY1XbC3zWqjTVJbmYV4jow7cSEmz+ZItKcXp4pviRTsUDMpiJ+Eggq
kSlvKUZgzEf3iWjR2SGkWBPy8o2uKHDXcU/8Qg++FelsjwuU9Xpb1UX/xPCf6Z8J
rwwAoZXxGWpgGXHdz1OXMVOjNFLZPEfSbUVyrb8W4c45/9/6tG++a7ItnN0c5PoA
z7dO7Bv9QoP3yUDId/weRb8J1gqLisoYU/TTMgDPsSvT6MrEUS+QUue9R7ZaU6Q7
5gVCA1+oBs13QVqgCDOv4vMJBw5IuGJqbradX6+/tud1brK4qVv7fTW2kvLEIH0N
lV5h5KectPaqnbeLNM8oG4FGbHNol5s3+lKdmF+19/BE2E3alxL3GzWiiuvCnAIx
bhkWmSBlpb5rJwBZU94KISdlZj4JVc3VtPWWS38uLQU8fg/9Xc2fYjMNrwUtBjax
mnkG0cjnukJe2AlprTParekhXRtuTnL32CIAiP4cUqSDH+l7pDzY+X5N4ZQE9Oc8
2M1S23yi/5xHbJJjvUOTbqC5Pqx+cSjqxS0K0L0IuTAOQK4yesL0UmAtcnkOTqJS
xG1yqfoDXcMMCOZBgfIF2qM+AuV17LAcT/CMgSorwtszNo8RYmuhEx0BRY5kFF6R
w5QgfM+xWIkTyIQwVnThtjPbtu1igOWpp1I+HPXtUpbWdf0/BKsRdoFQ0HCFn1Ko
D00smjfbNEZZfzSUkFdUFI8F+G+Pz4NSo0V/OUqA9bcdLJD6kJE81QQ8nZrROp4S
568YrGhXHWfr4Q2pAFPcAvJEF3ujyEAQ47pbvWUrOdNLaLPX8tz+SMXxFBJE4M6J
eiOTCPoX3A7kHNJywdsxlcQosRf3BisyBvPevgAxJjKMujcVHtUwbTcmfr8jlB9w
h9sBKWjfgbYhXvNrcR4SJy/0A/sinwjl0dDTfz62YHqlBMipdx+MUQz/8Tog+i7F
RwMbrbTGrSBnZlV7supwADB28En4j135P8a/jhAjdEXG74ucq7JkPjnRYhzK+NTl
xjUL8uc5SjdJ3lHlNEt76R8hTWQgBch/35Jvu9Wil2+e/84gNmGI4sp27VYrEnFw
+gkAZzmQTOjGnkiNVetJDzXQErd/DWZP/uFJx7idNBHzE8GlPbrGBLNVzLhQNOqo
Jxoo/54uphWyw6HGjhreEwZXSnNB2tHapg3JCcinxyZpvKugyWY258ccDRM6ECac
d2AvohjbKx+UfdokgI/SYsMGD6+saT2SwCO8ax8atxsZoe1jsnX4t5sqa8Fu9U6y
pc9itlMnpotaEERwEeDh1yFGdwyvH6oXEVJ3Q1eoRRR/E7ydOlaQTO60UuUoyD7/
z6h3B3wTQH3ijS3K56p6wDtswOW7cqSvE3VwoTs02U7KqyLWpsKzyTXnbYzaOs2T
B0GfY7IzuCL2yCcfWLbj+7qK2W6gPQEAs7tcDJQ138zsIdMZIPoBNUWZ9fsXvk9z
8CqpZvChTYAJ/2+Bfb6uTGuznixmy+eyzoUXVWzLhXqGgwL9kL8Uk2bjcwFW4kLE
gCuBBCU44Y6NGj/64kqi2FgdNlhUzYsCsR9ARRR4FMcFj/SGp9KXsV/zOiIO+icA
rrWIFmMQ1wixCrA1k539VFOtmcACbrD3KHYF8RNKL/ZpU0G119ycRYYdFGuQOyzW
P3T6GkBWtilrJbTBC8mr1sbvizzBFgXCh/j08JEKY7Bts6ZYdGRd1NcXoZ+xGAfc
uU6ehXq5hqgUUv55cSga2Gwlyz/1suKAej6wIE7LgwZp3YcUUQVCJ6oOztnqjZ2D
wxvrg+bFc3nRzC4p554mXTrdwwI5t0YVWF6nfXwBOf5wnuWY4liflxLuK71urkU8
ooEp0bVQu9j87lZjyvafSVlRjYgubofM/F/rlsquoH71b+Dn4+KUB0T8FqUqSp7T
hLUwLPG6bbVJuShsXykWn0RrY+WM+5m3Drj4s1O1z8vfkFSjaMrli2L7pBXVwezT
bRGbvuyZ2APEkCmTl+OHVcf6ly6kGdgfonMFqb+yw5RxPXohCWKX5ahTbHbA36iS
e7jog1ym7V+Zs12UbKM8hYsX4KkxidzYJGk3PgGdVv6Wlh/pB576D61rSIy3Fp4u
1XGs8pqXQdq45RGUQs8KqrMaQABqXs8LjchNEwEN3okJTKTQPULD4colxi5fHcVh
y0YpuBs5ymGQ2fMxIsdKXbRUU+WeAl4DUb1dlvdUhzC7uq6OH4lePqYh5foE914d
UrNyGJTKFVs1HSNZJDSB7U2NiWGroRg7/HzJ+pxWTh6h05hdwfhKaCd0Ikj24FX2
vgmuu2xFX9izddyVNFMWc8Jq/OTWBnVL8OemmxfsnjAwkm3J2dbMfKraWx4Ij0bP
pk+O3TzoTp0s0dXehZziO4AI7ldqm/UGtZ2clLB9ZAl34LkSaDpoJ2IAeQgz2ZhZ
8ioLeNGbpAvIfMwe8w7jninCGZDbFtFqGbXGjoIf0ao3DlV26gy7tvKgyUeWJWEN
cFVboNKSWK1YVrIR98rV20w5n7Kgxp8qVNOPBaW/4UDpr1LoSzSEwP7yUNovpyY2
LmnOzkaMl26/JSrsqoXMcL3IBbDjyo9UskSdpE1BCat0K0kA56+9pygYakIOPige
Q+L99TQrqx22/PxxSFu3twz8cJ6eUPlx3fXUzDJRX9NLX/GPObCUDVc46R+y+Gjk
ws21mS4DoDLJhcX/7RB7NnD1gOVmp8b3Smqo8KczQzdrt1tfVXl8eeLHA+afCr8O
f+ewsAx+GmE5BBfhyb3NAyJryk5VAVbcfZh6r8jIKAmJDVIZn3Z9CPIOHtXl5wD3
tqtb2XN00xhbiLZy84jgaDfWZ+atRAkLm1qxUGgb3t5YTv1fPyLqV/lOns4mlhKR
jxDK7xOX/CpXIfvzmR2NBytdtQDtuPv5rjsJVAcX7Cvto7u4X4RyuCkInj/sAvTN
99mmuxYjI7AKA95ZbXt293IC7MuKbZOE5T63mb4J9kuoDrWGo2YqSfeXIShS//Ik
RD2bgjrCnIm8u26p5XMDnoDTkW3KymIQ85XmOEKrDZt1QXwm8LL4E84oS/wxCc+X
enCSkPbVlkT1yl5vVwK4VIUOtKsR5i+yS3zNCy5A5szWbeJ2zdP6p7YFBz0jSr2V
P+UvmoZCYXmTuScIotaTdse/KKFdnn4WSh1SWZRQOMpZih0+7nws7MBMi+dgYKIQ
BaDoBGMBysmKASgw4JFbSO41r/d1xwOCenG1hia8g0UWanf+Tqkrdv1jy6wv5FD3
ph4xlwSnutPESBmZ2oMpHZfqgG2fnD4Me9bM7/egC1akMk5Ma+czrpSdklbw2mb6
WNLpBQrCV0aKJ164Gun/uMmvb87o04RcDD2khP0+qF3aRwfYooLwH6hXQWp44KZp
t8ZIaC5kx1Mo4Ji4XD4kB6SXLqgxlxgYsLgIqLArL+G9fchm6Y9gw912rHYufaxG
xmFLce+2e40QWKxz9ptk6t1kP0quoLIQaOJF+FkTFa0cPqp4q9cUKADJ5aYHK1oi
LToFjyuGOb5t9v0yZDzdTCtMx9smq7lJKa+i4uscpEpZkpT2Kl16mGMeSb4ime1D
UZ65h0J48bTKncErVhH4UWcv4K6ocXfG4qEBbG5MWhgfcNfl3MGz3HVbfiBM6bWp
hVeVM9dCXsVA7lSYhFQhTEcin9nsD/lsuhTFFqn1UXWgujo439t5fGn4ZdWEpiWF
Iw8rq+L74LkqwIT55nFg3c5EbdCoZeXf4uwaqnESD8fzDHbO5rnfWQD/bVpMkzAR
EgJj73z9yumVSdc04uH3Ts9Tj4CH5nVtHuegL54YD645J4DHBm8Vg5y6JXj0tOTH
YnT4VZXaV8Q3M3H0FugZNiC+JJqqecFxwCrMi1AhdLVpI/ewOrVgIbUxDAnaLcQb
E7CKYsPtfiTUaZ+6kLGi5xSfiKM0QJ2iIJsJA+SzOokWSu8YLJBEsennKZ40Fwu8
n83M9UvBagwNIqGfv261ELrspXndv0CEdOhPim5qkXvOhmvIbyaxaOrwOwTJIkx6
rNeOgmqUr05SPHmKK4TRMdF3gPuiv/CPnHSwtmL+0qHlS5iMRAEfTaT6DUk5eT7a
1TqBygNKaPyt8N0nU/4BRBkN/xbTSXSbmwpNsnaI/mwQQsQbcNtrUY0ZDrMO+6y1
3/C2mMDx+wREH6K/XfhJEBv1X83AGhrD32t6TofLQc22CheM5fnWAkM7tY264X1Y
Dp1FWRttVcmpbX2ZNnRflJ2+sPD0A666Xwd+tQ4PxpBUEfQmkVBlAsijXF9dIku/
8T5utY/n78SFfENHn1Tno1qbSYGNQtn2U81C3Kg7emm1fKaooWfWJ1eVq03AkvBc
xrxfH35Y0DZzHFqz0/x5c4f/rXS8xvuBJBII7IhLNvlwWhn+7wYiP/MxtcR3opVS
mz/hc7XyZ+IHaNCgRvXKQzWgZYyLZRB7BVrhvVjWLADtAKXbqq/dDw/okHRgtYt0
7Ja8NilUBcQumcU8a5JORqqNnrcrVyKI8qaOuZzWZm1we+1dxonfPL5yJSNwrwki
a6j9kQtRJbqP3mA9QTi+3KTSZtwufGKnbVHGIwJdNHNEi6plNv4HiqCwfm+oKh+K
6h64lTiR2dlBh2aat1FD0NWM1HddonZdq3tFWtxwLEvxFZfg55VNWET2TqFRfJDh
0RhYVU+M0zsDS0PUrJO4yVMkPDpbfzakPkzayFf6/qhKCLF8epKBQlqpqDX/G4dt
xIpNIhuEktDMtXrrP3gXgroQKOG7pgiMtjbF6nKd35hhNDhcSgIEAq2aRTh48coV
EVzIJ+PhqDrYzBbJ9r1cq94fNWyW2oWooyOau1RjWJtgm0wi3v/63jO/KF0supo8
QYioAJukv1Nf27/zzcwz0qvSNo5yInxDMhUjUc/5ra49jyOpV+F+PJT1/cfN2epT
BMz+U58MJiHPNSHpHQdzXHodjMbyQqVUbqtiTUGmvSfqSw2029zO87u6hmiuqHuU
A7chyNZJIq7yxLBbWTEKUXXQvVBoImgIrpehGQkcHm99+AdTJk2D6t7OATdtRnnm
OoOWkupvb24QC7MMe6m04XiCwvaj2fpjAyi/703oosuLwZtGBudZi2WS3U88EOBI
JPyf8q96IxqQdLNvL4GmZ4vUVetilnr7nJF2+MC1/qSDPAiu3PiKEPcvoE2oyLcb
qtODy9javhJAlStvF53sHA4umbzYfdhLMtbYamQvj43q7Xlvi+nQipwzAGxODLl9
wtYRKAC3OGIJUCofF4i2uH6AnOpNLG87Oo4sf21mGjbIuHAQNCSxSbuHZzWn3Q0O
zkjZnViQ98nSb3pMTe6V8eZl9JAUWBjlK0VHYnV96xngCFUnW2iG4Nyhm5bDuF76
E1/vVlikHkUo9u2j2IYND7mhIxfd18aDziQhwM0H6LQ1Ox/vS4hIkkPivIHU5bst
WKDJe6QZdPECf4P8xWEiEaqE3khIQcIckz68aCYtUYPbIAEzA+TbDfuO9Zl2NFy3
q4ufJuwMS9AQ5GJ0LNaZwpWZ8Jo4N1FtfZTVfUrn6Vcj/IS8dn4oBLbzfXPrKJ4o
q4TQOX/VFlcwFBZeGX6lOwPqRYZEeIaPpX9iI2+gdpVad5J/qALr14wU3U+G0bj6
cM2f8rZeVCrzTuIVmg+owTMQNM32ZNshmSmSR43kgnj7Pvok7K1CmCXY+z6vQc2S
w2XgLI7Z2xFXPa+HRWHXaK0vnvQBU+6JAdYhhHb2wRux3ASsq5Hc8pcfSGnFdtYt
EDUl+ZYgpUCx0PgfMNOPwyAaRiC+VPCJb3FndMXMHcAss9TGOe9sKIcUjA9vu1qI
g9zHyD4z/KK4DkgOCFo6RKqCe8vlzudIGJV9vUIxc/h3pl5e49S1X+EMu9oiONs+
+s2mUHNU4DLozda0fNq+1UdIChnwMm3Y+saL7fvBDoMfbnVvSYTqBC6QvZB8ejBZ
2CgFBiPCQd/RQRaXdm1AvbXg0BF5pMqMDFO0x2ewtxIxYWgRt3oqVCYV6RnyRJJR
kCBo0dVBC1YjuLgw8fZWnp2pXOhoYT+XK8apnPPPfF+bWK6KvEE+xTvLWlFCUCZg
vKWfaCyCak0x6rMDfyu7nl3O2VAEADgJt0jL9IHqhubJpjsv7Dzd+J5ExXObT3bv
FwrTXLJ0/uWtCvYNSvjU2f+I0rTFros4hLwff7Mz0lXDs4mvkzecT1h2iwgDDbyE
HHr/wU78QWQuRQcJFH5xwdQjYhQTjcB3MZz65EUImsOCaVUH/LRy4r0XXP8wL3ON
fwwn3ptw6ipynJtINBIjOpUxc9jZxEFZWF2QnEjKewaXjxEsnGVNfcEy590sRPbe
ND4m8Zje5mAw8st0eqpDqCBuPiu1oj0IWYg9SCCeleiX1Ztf9DmYYbUUYxj21fzl
H7xPF1fAbMiMAx6yKJuXx/KRIw/vc/M0q5vwprJS8ftR4dUsXpI6Pfk9zYYq2vbJ
qlJjSFnu4gqIgsZOfmzyyOF1dCy/Qtn+WRHZb1dz+ARL17F9KL5DTQcEUYqP1YSq
bn0c9DUAw5fP42KkqqanBY7/0S9/uFPlI2mbyqDL48AL+RzT02WxNR1hEgAv1Smy
NrTXVjO6iwhWpfCG7UppuB6t0OQmfo/q0L1Ijsv+m0Qvw/YuGe1lYKv00gT0yC0o
POaMyjgt58D4NI6iFCRm+hnMUHOUL46fei9/BW2I0KmZtDhJXJsCPsAsI7r0I41e
i9XWvfE3D5Eus2ef6lxN/MYU/t6+4+3oA8V2X8vZwkhL/pa+Di8oAT7WEJAFSZD/
SKT7wdvpc+QiOyQ8gb9I4RrNqh+ilxmpMm3l8NJhewP7uzNxKRh610BS+h/zcjZG
9asdHC4T4rkkFqdd5giEOuTloVJk/1bQk2sdKEzcrjE=
`pragma protect end_protected
