// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UiY8PHmV5czoaqJOmfuG8+ncaIXEabcuw6mDdz2osBSAbxejdiuldiag6Prt3Fw4
hdLbwh4akPgHYWaVj36sL7hIHm8o85p6k11T3dXF8vJcPiAjHxyjWF/gRtG1SUkg
IXCGHFKCxO4rdTBRau6jBZFUZ/hnNnBWMUr0A8o2v94=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15376)
IeNVEFaoxHzlIYuX13YumhHFBmuXjx2EvTSsi7r9LRw+ZRV9uABYdlJHKGNVSelc
jd0L8f+DbgSv3nEdtxMVj0jtWRL/WYhnFP8BArb+isuFlco8M6BSNDXc0xBd6SGW
K1snAZAlg9509DubLXYJtV68jhHi2YKHo9aaCI7+Uxv9omBdC2YobgdWfTDHry6h
K0bkdVcP9seuRzbmE/4wv9goTt26PMjTzf6fzUchHJYE4SIkGztVHAsE8kknTQzh
4kqhTtT6GKnH6jmHiO7dwnzlmBxaK5Uv6qhHvEAiVczmPb0cq4VuHp1LhSFnGfnh
1/QLAEM0Z3ahjnmc1SDZtU2edArNV1kcu0+lmj8nUcBBFb3eR1g/+6xbciV0PkMD
rGmTp+iigTiUH3/dpAbJq9rWrFa1frl7lSoWmNqDrKZErGpGbG3SXUvu+J44j7Ps
cwBP6JitA8qzqvd0aowsbpNsZNVdPc+vOadvCE9Z4HDhAevfl8UKF/JXOMMV+VDi
GX6Ts3HBavve1q/0U8avg69QW5jB9MIS+96IjQvhpA/GkDKw2R2cTR9oyj+Fkiqw
5Yv1JtfrmKJbtKpPFnVEhXuyO01OknJ+W0XFMEh+YdOBEjNlTvvCufxmp2wyEk5E
s/JLSOMM2Zk2CoHohyxqZu2oP8b2zP8ASAt8wcTt7nv8rUlRRjY/wDHdAYi8uAIy
bLGUkWWycttANVjq587i6ci2xFyUrQKT1UCgXFN3yyDYV4uKoXRXQBy8pBAhDXAw
JKw4c4guUVu/fkLwUzwDXfNnA2RYaRrgHTUQC4mrHxFL2edFHT5XcRiaMzERZkT5
dgQrDkmunpZt8ese/fIDMChAzAlRPZL7yHfDwmXmpo5cXatsn7X7JlGUg8XDRPNy
kf6rTU4PmlyvusxWOAHFfjyAXS6hEmsJi9ZsG9aJ1evbg6F+swnfqqqegCYvUs6u
RDqm7pNDSfzHGE7DLFq2mlMNJfQlIDPf4EcqRnGHJSfneWCgeD6njDHhUHkhiFG7
I9UxKFJY3PslKPp/2nB3vqYaKStFDa6HPq+UFjKn9StmgiVns+mU8zpyfpa3QnwH
YNVYsYjpYCQYdGvTfBTYrY/ARE72fjq61AdlnCH/JXRLn6BBzTOAthtT970KkfqU
Ia6KcK/umsU9Hg+ydK9ZaOftEZJbHKBAPq3HVcMWT9Uluvd8makJLYfnk6gK7CyE
XfT/7QDY45YSYYTm9ikfWUBT/Vg5x//JaXz+Uj0cTENSeDDioCwcL3JTQLjUiS/x
6RCtMtY0Df0TbkEZ/cKLIZjwenhEv+dR0L44jypVLcz6dfNmd9LyIhf2t2o/4GHN
eLAROWK/bA5hhPHAl8zMYX54qezcp22GFwo1RPb8l/8ExtFqtn/gD6kFKnKzJ4ml
hHfCJXv9EDaYcbMsqZb3uAOmFGX1BQgjj/OmFNwfgR0Xyp3BbK+pk6t2MLuxjMB3
72vOY/yWQmCkZWytii83GIggXnmI8fAizYcfdZ2775Btw8SivdJbmTmYgZ0iOlQR
6XT8/poaR+ItoNJg5XFAxRj0pOFaqCWCfWsTrKB9JzVSrEehR5e7f/0BpM4T894Y
k1e++4H0leoz69aQJiJclXvMWupqwnvsP3Sf7Wsq6mUpUWqk2U3cEnxMhcPna86A
YR0p+7ba18OhI40uUPa/mY7MIpVKIBJ7vL0T3rlU3QZ7ldZrzlnz4+kSlHAqkBp3
2vz5u5N1ftUSzcZ9r5MBr2pFf/BDQOnr2rM7XwcVm43nLbPYSD/QELgtbDiNCpij
Iuzshg2wfetwAi1NPg181Ni4HNPENQyBS1tDcY+I2u46meTp4MoMPP2sByoTVoGF
Cx+3C4DJs/O7C9+qY1rI/ELfQTXgoDBZs3GGIlJartnZyDJyuZyfYt0YjGDRLvV0
jO6FQztqQ+OSq1/qmlTis8vnpjqXYG/DpM/MFUx8/t7wuuUmaLBSu5s4gg/nVujT
Spf+aln6fMSyQqZpR49UXAaF/2n3c2i7mRHaRoaS7iT0/rZXOFe8nBOWoFQn+SjY
8Q5syyKFzAy1Lxe2SeWPmbAw5e7E60IldojXdX3iRbWW2YsNnhAwaB4fdmFLlusA
9H85Sw2HxBgOoM8Li9arhz2fZEfFXnEHmZdFFmBk9lMDz3rdI1LZp+16i2j4KPEw
Y3XRk2o7PZ0FH2wzc+LGGyHyGz0m/KC2FoUM+lKYSmBXC8Nyv+c3yYmlLy7pCSa6
ObG1Gb9pR0eP5xTDvztIynZXnPoTvV55CG3HHvQzWB6TZwxvFYJQrLGIx17h6CxO
QuB19fVOSh/EY87Hxjdeep3rpZgBkfnYzr2FfQoEkuDaQkt3Ogngyv7n5UCWv9je
OKRvfQKhOzXQafWw96HNo4UUshw7gDw5wj+QEW3ajLaJYVzrHmjNwgiYfuhup1FE
IFHGOufGkUE+MIK2Pz8gnzpzNCFMIh6OaZgh+CnutZfZIEfj4+J2eo2jeqH7laF4
OqajDJ9NH+i/CNFe4PGk6X3ACiAZgZH9dPHHW4POybvo8tBlg8J+3YLLQM2n3Aau
Q+jMt/i31yx2eH57Bacf1JCcc74CSyuRMPzz7dhOBDXxSmII8NGjOjlnJGizJeA+
hPgl2qWhJRG44fizyUMw7Ton5ZacYx+h7w9niPY+uCS6lVdFl3MMgOQEpHpJe+Ah
2pK+8G+4ExWhRTcLMdjt8FDeHn+Xw5PBmir7ddysatJfN+75X3HSSGE2E4SPNnFX
/vL+VwO7SdDfwb9642yqmQZ+I7YwxRMSdCSOazClAxuO453/HNt6FTBjLr4BxYDU
1OKn78zy+bqBO2vm5YMUd1gZ4KGQ83xiY0I39SG8jHLytCSczqHuU3wK9HIGFSOI
T1NKwhBDx8ULfNYTlrKx5349w7c6YXheTcud9sS42bU/djHDNZ/Lduc8BuNu5INN
rdch4xCZRXEx/BELuWJN/EM9wqKG95/PlNfv/RRsbqITfoRHiTJ1hG3tdDagCXU3
w3hEuN4KtAGuv27kcVtLRVcZrtkDduOQrD1l6E8GalnlBFnRSnIBMrIf9woRCYWe
kN7oz3cJEq6xt6rMBiv6VMlkVoVDcMFvi6ZwDN88dy9sVVPCIp9wA4B7g6cGaio3
fY9aPoPEckyXiQOoqErnVS5ygTPC2az0k0ndH0ijSmaF5pYK1VaqofXpnWkOwfqF
0vhduXdxJlpm5CNU6jQWUQZoUdnLFMmYhE8qsyeNnZUqyvtJgwiYnnQTKTx0GdpA
F0rOFg12mXLpsGXSHorEr12yTL1nkGzyV2Ajg+CQKV9mt0avDrCKIYynfzLb9ogy
RUBzMOVeuJahxfR2lyc26S2LjEB7vkVFFcKh9MfUQJXtOexZIsBQAnJsnBWgV3s4
HNcKf0eA8H1m68gpNi/vmemff2ubHQChRP5reGnnisxD/ptVs09c+eaouRfotTZl
OsZKlECBh+pYrwQ0Mbqw4oljX7/j3pcsnBwbqbMzgfzun2IFuDJJUTI+04dgCVMU
vVaDS7uBl8nwpcys9sY+XFTgf50xc/JSCD9d3cOORVzaEo3Y3MFf3nQ5UmgKE6fK
JsImaWsyF+V2MKtEX2HxMb8vKBLChm6PeGNa5wEzYtwQ6Dqu9v1Vp8Ogo6xAA0z/
xE6bHAVyJjVSj3AmyBf6KIlyDORA82dQnAUAcfAPE5tcdeSsUFphr2HIoNmYhdqo
797H4BX3yCP+0jujDiAQMbcGB7VMEcCYpaxtk4VPvPYJ5XltOL3z0dipHp8zwimH
xdBdGilEgEo2hhRFRDd4OEPuIJfL8s1oWNafDJsH5gKIX1daABk4dC8BdE0nMoLp
GAtsq6K+6bx0LirpUP5iAh1WbG0y53hmzyZ5hxLC0c7R9I3eAtlzWO0Kdv3PoH6m
UBkujpPiMwa3Xbaw9j247E5btQZbEegoVoqVnMf3MYntmE/rEOJ4JqU9dzNNShit
nBOCU4hKh9RpYH2tcwbK3gQwLbq42Eos98IO5CmyFWznQItKIW41znZjnpKrYoiT
SNaHGLgzHFa0bGrbq70rKEkZ6cFUvs/fZIkuG3zV907s5+1CCcutMqRdmtHW01ES
yHUnXXXjRXxi+wEUZqwh9HgWS1k51d7QdANkmE1c6cM9dQ4SWvFE9C6iXjRRrEqg
e/h2DwbVJdOCkYgQ+j0lIkr+8PQ0ohbh8ftrSskzymwVHpdm8YMqeBuu1jcV4FoI
i3DvnmlcWfm+UAqM0SokhY8qYX6ouz8z8+RHN0cQQq0KZ5E+GbXP6Lujn4J7AULS
X7PUIqvuoulM4U4/j8g13rf32wCZrg7m0Mo88tY0kePJ1UwbxADnM8KxuKZkfHPF
jkrl3t+Ftt6So39ivtuPAcAxCbhg2qyPLXToJS1+2cRxe9599zNSVbbmEn0ekvm2
dpLqX62o6T1R1Zz1Z4rOKqvxUl1zFM7z7xRXr3sKfEyxc1TDQxSz/D9n3yZBwnW6
s7umMt3mwhc5wXEzbV39jklYl1g0gNA3uIDym3hkOy7jrqMM0yWuRShz2OxSCSxr
djgq/9m+mIXjPPyWP4/GULKr9qxDErbjXtIqr06oE95pqpofI+7dGZrGg3Z6ltyZ
UCHTe9ZZt11SFeKyM3/pCS6kGMQXxwdsBeM6RrDZy/SYABc1vfCGKPqSnZPmnKDC
OZbFOxq+1AXyxWpeFTAs7E0y/hVjq5NhqYYEEwUj436/C4La/wqKymTl1zI9vySP
PszIOIA0vd1W38pVor99g4KgOG5MW7Oixya5NZ2LesaqOLcAg4sW957dAjylNfJA
4Cc/dd3n0zRJls+ciaecCZTEGAy6QZWsuZMnRleihkwW8/6Pcu5mPPZC1Nn4tSew
2DIPKwN5ZlkC+GecogkTKtrR1D0WFP6iLTzDSbY6IIaMqzSLwIQ9qw7AVUGAwNgb
w3On8rXYUwb++ZYjTYhJXL+JbmqiFKPM3v27snfiwunDK39RtMQV9edXMef7MwLd
CONu3/iBWozk+jq9yN4AGTkRRt6OGbySF4HBVzDCpnm6uPdg+NdkNAlXu80+rog/
U/ghr7tr6ROe3IrP7EJTsrbnuJ4gRc/w/lG2FIHd4PEwmSBsCBIvLb0PvqieYhrd
s2zfM/Ok8aMnlj8hcf264Hh4dhoNh4FPMAb9wu5VbAQL2s8Xon05Z12EYKBCgMgo
+NbfV/a70f6XvxTTW7oEJzh2NGl0Zm+jbmUo6dq80R0reHb3uEVOjGe0prTV0MN3
xsYPbxh1A8jMBcAZc+//aH+FJflaFotRnE3ewDQPNK+XqYoAnv4Y6rtLNRo03OfW
6wyo2Fn6XuK1zGkPLL3lTNm68GdYKmrppPAc6G0REsKzAgClFA5Q0ebIr0abK28G
LCQ1uj45/UJp9bHOS1YkWdnDA7o0ZyWhSPukDkWO3AJZy0bsqgJnxxw1mzCEgK6c
nwVaPhOjbI1XuMoZuGZYv57n8s26Casvl/YX9MWtLw3rfqbeF20pPumsdVJEaSKi
wBMG/lsflwkuAoXFO3RlupxwU/pMYVgeVSXH7f0vzpfREdydh4hP3fyz1lgdggh8
0RF7asoLFuczGfjJTUmEageg4QI81aHM7MORo0cG63iq4K50Pm5y/Ik8yAdmVEkn
hO41NfjLFdsnxo/QNLuAFlswCSVXx7EIgBaGL08WFWaVprUtDf7WXukrcOJFzrLe
rkvlIySfQ6dIl084s4fgOB+gJkXm4axO0WsZjW1ekp9psdqcMicTSu4Mt7PT5iSP
8czY2CrY54cX6mbFbFDhjXCJrevu0UY/i8ScCXyBxdsh33A08Dxaqo7x47QgX1Mp
ZMkuDf1ZYKPIQfCfVJGZgJES05ZI3Lq03mSXTS+2i9FRKFWGfgO3BiZDay2Bo093
7UI+oNEJwoqFlNuJte6WUQre0Z+xF/wotNSzDcK9qeqThpaTVCpcVMmZtAfpk+3d
wY/nWR4/zLoY+jz1cj7nQan9itTORB0QmXMQxaGIJt7NdmlB2MMokS9r/PrTSFG6
nJh27XyWmNFPz41JmLe/v6rhaagv4pVVEGYoMWkCQ9KTXQzaxGFXMxgTKp8t5ptP
7WIX48id+H9FP6MoMV+k43lFKWIzwrLzbSasP1zlU3oCkn+C0IiqtUlBDNIu2v/B
BGc+HHwgeUxg+cCdvDfMeymVuohKCIgIG+5PtfCQJcHgxHrKO83RgXn17Ub8p8Wn
BdgUEWGRv453EGbAwzWwe47UKotmyS/M3TqzqMRqo+hwsyWGk4LjSorhx83rPz2J
YmCnlfxH7leVZZ3ySraKbCcbLNJa9NTr5ERhvoNnJWZedxfD4iL76bRhWSVU1kfd
mj3ZeHRO42VPMEowwxKlszZUN3SwwVe1OoRa4Sofv0jqSoxcLJUJbVC4sIxOVY7u
7DkaTRC6y0Rp7eMckWzI97UZT+O7J6YFscdaStzpMexYbew9Oimd0waiifl3VhmR
8tGkdVJjfW2hdE++DyNXZSx6VegJ7Lz0Q7+Th7ZSHlK65N/aice+FAzfw9huS5eI
vydYbeoSZRtPrYoXowLXCPk+WsS48ffi8txAQNrG39keQ5gLG5QUAZGlJ+Q2oWy5
y1tdr4jKi9bzTBNhLgaF0GXWVFa9Opfg2UpZMfvmts6NbivQJThfq2KIvq1IW6ey
gPea4hsaWZDzSqNmujQka2nXutCkA43rAVCZTEzaj0RWQba/rhxs5d9O+OoHt0+H
LD6M5HN2e1EDSLWNxeFP4kr9jt8N8CQzzahPrvt/UbbWQADD8EY5mIF9g6qsHO3Q
RPX+Nrt/32ooWU3pETyFrxkuWStbUvaXwG2O4x82Y+w4eIrtDZfYup9WRHIUUmF4
AFq9q9RY44mkT3ci51TMpQjTRUCG+ectyNOZpum6WfDMLfcLBERKqSWGyOYwGoqz
3qCAgxeCrTPDmk6KR58+AywGj6YJUGF4uAMkGF90IrPlOKgJtm4On2JpXUUeUn0m
pDhjC5CFsYJSj3T0pKtaiufEcWEK0WC0s4kz82COKKiGc4ydXGcaEaLgrDVu+ALT
XGfThN0E1aIKSMwoNIEY26VMmHrZspNEX/4buxv9SIbHY/errthOrQ289+a3PP9J
trnXkpganXSppFYj/niVxKVGtpMWxQhsqAte4ztsSIsjFYAy0VgU1bW2bhFKLO7s
ZMQGJOH4AySHMTy970B2E8Ho4clliVNp3E5zGGwj82wk/ponlICXEYWmVmc1ntoJ
ddX1voAcYyZiZI1KN4EWmmFlAHhoDZsNGm0hPzIMCT3RS6zBMJGstrfqf1P5EVrq
YVaiGbdEatRxhEuUk2c4fjd+/1OG6ZMwD0sOYlTGV+Pua4omix1yq1PVmRfEi74n
aSAZm2bI/fgX7p5eNLFmoC08FkELovVAb3dJmVRzu00KwOYo3vlWb+ksGM7POl7E
vmwItmm4HHKJJXy0oGCGgQ4bQYJXTK06drPasWzFyPp+dFBh4avGalW+gqRakcGF
Q/xIrSHRX/bqQIyhUNcGWqGBVFMJUwwzx9obydBY7YCwpxWcKbKYfRDM8SvijqGc
+fcJU8yLK3dn/PSgkVuuPMKA/EF85JcL5ltBakSuLHAjR1L0517plMVAdhPXo8Pv
9UHGGHV6E3OEdjMa09PqGbFrp76fB/bLvqJBf8jYQMaZwi/59lAtSG3ME9yCew4o
aSc6r7Idbzjj1DzSn3FOgMoXHTFGrsXxeX6Imbas3fM/HuHuEB/aSKE0VtDcQ2tR
ODwcyN9a0YMzvB7cGkY6gYInfbvRlhSzWvPIKQJpb8imIEJILcsl1z6dwYw2h+j2
vx8/6JgPvQLbAwqJYGIJtYBSAlmnNjWPvUXqabqmHOgMterx9SZ9U4eRxHbJRhZ1
59XiDsTTFuHOpdLmCWmG6zXTIfZa/ayLxof/Lw4J8FWBdVz1QhB/mEeWiQzWVQtH
IXRk26gZCyjDP9GA0uSTYHJOY4Bhr6U8KKv3dmempTjRaLJuSnw3M+IqWGTh0JEb
rg62l0f4D5LAHfSquqh4dcqnCy+GlWl61lgu4k6gyudyrMGiP4s7xE36Ijl4m5Im
lag2bRAuKK7anZ/x4bEVp73L62UlUbvVXfqz6l6PXxy/QScMhfVSzArlNevEh6so
nG500HlPPqgZHz87+zA6Rc7Lzs4EuiVkdvqMYzRXLa9Kb+/dTir7ZP1xZ8vNOvxS
LEnVSwusgGB1+C9sozcSW+nJ3g6y5tPCQcQBF8qXYhLF9QBkwg9KJkisUJHpBncb
vP+Ga+TpEtx4vejQ6DnjuYOPz0gTIsjaWnvWTxgioeSxOWJvqKG9rk2K/3Vjon+3
qRXSFfvRbF600NOtibFMvUN+N2/wVBSBYnFpXzIXOZaNFf/SXzqBEYUYPIjeAJO+
87+CdbjfOQLqHwnBoL82t6arThPi5Y+DjWvJHy6BlcaV/kx94ucRIumy6h7BeKQR
+r7x8EZqZttOE9zLYfBGLJG6v1EYOc88hbmq2WTUE/CMpISYEjYvq3nDVvYAV+lh
GC1wuK9vdkFPG5PwYD5KkiLcrcGYUpl6bcC8vvnN8gfhwb4KzmqlugyFX9RbpAaZ
NTXWioP+8qyFOCLHH7HBanBLcieZgp3MIVYXOzzDLpeq88LOjXylFXlPt6AQv3TJ
pOieLxs6f32JJvPqIqg6pkuBuoBm8bBnUcg34phR1WLFo/Br5BT0fl264OuVcY8F
o+FdTWhELjqlmLNv4pFE1z9KAmGAQ8mtOv/d9idjeJ3ljrxrJkkItj9flZsHpOTq
7qoZHm1njEoixVRN/ngAkTdElPclYQTis3UOKJnzCUE630Y88fXHKigWcIsMR5W2
/33JAlNEJS6E4NZn0pSwIntEuQ62IDbYipCad/7VtivZPoskjn+MdZWNohNL4Ozm
fiXgTCCWhiE8h4zayiimNC9aNsAD3wY3qo7cRT9CZfSq6l7Li8tY6F0O/zYPHGds
LomBPXcyp6DLJOORJPjxlBSphV5OJnnP+dmC3YvfIjNCvjGxmuMiK3pY756gtxVF
PRTl2vsUivXjlPfkZqotJBoZLemm99ZN+hn6niLrWjiezOGWy+vkMGNbMMKMg3R/
gHlMpsVGTF2IYRisGPWwcyuNZr6LXkazA6BeyY7xr4on7UNz3Ifkv8gXQzmBXKCU
BILpeTny1Ihf/FpUIk6GUtr3sSngi26RFHkYFctNqBEvplLYkQQiW3Aen8NH4F6o
Qx62m4qO73kP22XBaM5L/tMJqGN3VxkW5QMEsHp8oLi827ZIcKeC66D9VXePQaeA
4A26+C4Hz01L0DjTRHzI4Y7JAI1glj+dHdU9rEZ/mUjNNdpe5hHzR6nCoau82WpR
Jf3RTEKh8H8jMltymCJAr9rmNdLFfHjDBo/q+KzlkNEfCt6smtyT/qOPkg2jVLls
PEtRAk59542AmgHc6nnUL7Ie9f0fMXLKQYNIAL8zTND6xysHqXFnAEJ2M3L5XWaw
Al8LJQBHcvpjVxAInYfuubX8gHEmCOtVHdGisj8D62qE71FDLzbfmh/iejcdrKNT
TOKJ7/tZqDAGL26mhyzZZRQ83/JxKQ8NzP4Sau1FA/PZINDB9vcVhG9joZNBJtZY
PiUpWKu8xflmff/4rchvdEKFC2bxYAV+N3JN4Jkq4op9JiIVkVhwtnbven4GwXmi
4tPhnGOV+CXaI2Y/JnktMLWhRccyYvtYl9mvWCFq00Ix7MPDIXTroQln+T3IfrUC
t3CZqX/LROFrsQhjEbp3SVWTL2aRXFb7HPh2T9jnzPq2W9KWLTYPWfmhoB58osFR
9Q6py/6I3zPvyYFwxvThKAj5lVsza10YuqafyNitOqvVsD8J6I+QT9I9wzB00nUd
h/D7OYhJZkDWY9+ySBm+PvCmbYzhPsNODOgfXpYAGt78vqTmelbAiKhHNmnnvdGp
ZTlZXxbRi/0nSEdISAfIARJ2dpAuSRHqNgMZLVAuj6/x99aoAr9p0w6Qup5ivarG
3246K4e8lIoEp9x/ixf5kP/WPXTb/FCViAQgx9DFe21oP94T1MXga7TOlJAurJdF
i2A4kfLOa1LZ+M46LXyf2Ah+avbk/IfmXKH9jumbSXHmppZp4bkJH43/yl+MuHr9
a0etfg+UiO6bvHZZcgKpYS5jC2KpEHQ12f4rNKORsUYSUhRPhM7czpog2dQKa3Tn
FLC+ol4E+FVfrom6mVS8sseMDjQgdwOFte4/IPneliooMuFUcHF+TjWe0mQVNwoS
Dy+VVrkkAA28CiFkxwYJ4v9XL1Fsx2OHvH8Sw/JF3ho0ceu8xquKSjbHKIVBi+i4
mPD4drIfl+rKatOKlJHVE46buyzjRkfGixF9KBVQgPGy2NrYDUCNZM/+mUJj57ti
ejGOYZMoGQgpMO9W1zJALng7Z2TOGV4enpgQnYwrYCTwt1ikphxiiaRc3z2DP8wt
ML7Val21buCMua2OGae2cpJg7c8xsg99Tmw8njHlxC06YVzht16mcraw3OCzRjDr
74dYJZyjbSpeuLX1Hsz7mxkxZnBlZiEMevqMEyoUmuh8aGUOrE3sL9cXZhAWiIiX
+JKyATc2KnHHxQSBIaLNctW4XewzXFjajJ6KMx39JDywVfKj+d3G11sc5n5sBvFN
nZg4dzrN/q7jnpMnWjvsT03NlHZoRzKZxUXtBbDv14MLKHRr6jgHkCZGwUBAYC1m
KcQ8uxw7ENWuz4QdWgdi1ySOlyas9tUV8Qqw/AwqldrGrSYKN/U/3x6l2n+ZsUsS
38D+G4rtmcP69DC3NptSCeXnd6q1k+NcyE4vkql3TNPRa7xvWw/1z0ce2veJlCyh
prwiJ+vPg1FSTxw1W4GEW3zHjhalvK/75MkVvqW7gFoatq4OK3MIIDWOLS75fn3D
g2tTX3hniFsW66rOEoz7Qtb2JvkKu//8O9avOB8DOGylYdOPGHBezuMIsr9aZaXf
WPl5pjAEv8LpsCiIvKbDqTo50yrgYnzpyhG/btBKnxzS8OD5rQC/nem+44Uz+ODP
xa0b129AIgwN/n/UlRxbhKHBe97goy8fV23E2TQ2wKLB9hlMa0jUyaK0sKYoPaI/
+/OwhKJDqnL4gTf5f5dsdrumSs/cjosk6SMUy8Zeda/N4e9WlHHSAuQJkb4bta7m
wOL0dLx30nHgH7YpUBAtVWRBmRgPzGrWSxgkK1lnoUYXiCVJqfgFS2Y+vV2cbYIz
MdgLsJO6z07JgCr5t8IW0WevExaJ/XpoCQZ+ErMBSsrjc+qISxOe1gxHlYv/bRhJ
TtshmeyxhGE7YhTC/xqJgpyM8AdqmHDVznmLdBVvQ+EVpcmraO7vkkh9G3fpWQEv
7rrIVNCovAuQfIosrVanxdN83hds7IBGfqKT4NoEyTFSXp+BEFYeTmCQG0kvy6pI
VwwftVIBQjCrBuGyoR3Bp4INaDv5+9U0TQc6STuArHWM3Agl8mZIpu9yhzZ9NOYY
HuIq/VJEK+GznE4pMy5dBRwewxAGUb8vI6t4MbJ+k1K0QVhL3ycCtI76YP8yoKSq
sjqSnNcoMb6j+z4LwwKsmVEHuThsxuM4FumJNCbmlJW2rxoSpCNaRUZY/W3W2/+x
h9+5kT9guLe/U8YUv4x4J8v95i2og9DputB2KKOLQPSWYaxf2yyWu657FtWowILm
GTBZNk5hWQoI9lN9xWl+UHO/Cw04ClxeXzbw9zIa7WSK8XOr5TVrOiNjM2/CykNY
25KHWIipQMCSRfXepuJbKCkv+6G9UecFIPTze43xggkrlKRHdtNLGbqJNQcRFzkj
a0B2zUCv/Y3YCiDEwm7hsbvp5btYMp9x7UQKY6p0njSp3T98KBEAS85Lxy4d7+O0
smzAJoauH+2D9CTqnCD3qRtLDZhURTQQDSw3pndrbp+L52XDqSUbo0bt4uBLz1F7
J72+2ovNwz3koxlQwsPHkVCkIcUEviWZ6cW6cxwpMNPsdF3aS3uGK+O9EE3VsBC6
/RQ6QB03G3H2aeE1t1452IPmFv2BWtOTiY7m6EtteNIm78Jqjlub+YuuZx2k5oVm
WlLTR+uqjSe1N0b6Q39ytB8Ww0WVOZaZm7o1SXPY+mFsn0j10aV+RM+J7vFyax4R
J5sJ5Ov24c85F34ytjHzwv8ptA03U03fPKZK3Iy/8WX+xH39KTOaFtvEV/lQeOT1
qQwlE4P8exXgt/bmaQhSxS/PiaTRXeX0bMLbpW9mtiY9O6V6CNZv822ib7va0mP3
spITYFPKa5E5Lr6Rh5G9m7tLMZBOthT6QGX8C8AFRryTi9U0g1a2JG/KaxfGrwIu
+NnkyeN4I0jCBOAKjHHIXaC1RjIb0Wvg2gS6Fyk+ucOtj1aTXx30seC0xyNZTUBH
mt1Sl/+heLH49UBfyQC49QHhn1IIz1H8wDqV9erwjNcJduJkfNzZBFD7YsernTsF
/I2A0MkpEBeGOHhupoQ/YopkO5JSW9NIU9zqF6hEi3A7UBe3YfHFjV6l+koT23VK
tyTmmkBHX7XhFeT2m8X4VozU9jgmC200nGoRKy/sWTrXNg29SG+0e9Yvql6Vs/yv
1ulCTvl2hwLy2rygCwbZ6g1i5yTUW5k5Ju+NZbqnhIHcXqBqfy8xwGBz+Mh+dgxa
ZEPNGA/LkQUPR0qiUoFqMOBG49e3tNe4Q0xs+aJ3u63evltH6j8Baq1wdKrqbr8v
a2H3vPG5cXuRBB0y2treGRjSI71ElI5leIihNY86L8eb5cU3iwRNl7o2GlM1pN/y
DOD2GDTukzdNhF7UazuBZhkwPE1b0KycL8Qo+cNDAXNzKS13fu0yTgdN4Bjc3VH2
nIZ/T/gvX4qtL9EqCLcz3x1v68OwvpSwqcTG9iR+6g7+W7qpfJimakI7cpl8+233
Fl6J4jsFIBVIwkA9BAYo6b5PX/w3FkpeXbQqKqnFhg2MJ1Jrmc5DrQGp6+hEOKu9
WBMKX3ow6OYUiaqs23iMVPhZYzqlm+UG3Sc2Y8pgPXO/cy8uu/nevcUZa/fgzoKO
pf74OcBm72i0wESEk+3ucBqS2CXAEz7PQCrGVBoLaccveb4dHi7AM5NNPyhjLaJL
N0rXelpGrRddn83MMDWmSmoHl3VIrrZH5Xw5s5lS2Bxb8H1VNBxdYxg1i2p9PXHq
39TuPBlVfthl06ABytFAmozMol2dwqir5/yS17S8U4bzk0R543jfJuiGFDpz4DvX
vOFE4aRqd9jAu9lkDSA/iL7CxyaVIrbJpt2jrfWXnAEOwsvNo0STH6PhgGQVSyDB
hieSs86aNWHmGY4STCuYqqv+rntaZjW1BJXqbVVfRSXmoaX7y4xP5OqLFPtIAAFp
5AhdMLvmSDmQAX6efnWACdt5I1eIwK+GeGa9ymr6eVK2nh5/5/s18ErSvNnTHMEu
yEktVObvPggzt9XOs6xwp2vwCWi8gwW0vKMfgQakcGiyUTG798ajaBCkPokW4BIr
92iZifZSu2+v2QgLV8Xf6SSKYhxKF+dzdMohZ/GWKJu07bjALT6vI0gblWwUEEtn
6ybHfZyuUJ+j/DIOtyJzvhXRkxxFHAKyUFOHAk6b5CAvCGnHHN7NFBf559DsEioO
CHaTars656psqxuoNiELKauephQTOuOhJ/is2LXbtx2iuODpTquk1HR6ijXCpjqx
3hkObtSbkfQNPPUwOlnVKrRK74g/rYX2AjqCSn45Ez5IpB51oYb4IByMn2odE5LR
aN4XBWW569ggkWbYOlQAg3eY85DOFRKdSbGzVzptZIN+NeszGooVIjvs4iQE1TKQ
iwDlfTke2nL92xX8YWNfoLcVSoCQ5Alxe3nHcpyUJNWgAtBBYoIu2eESujqy5xhS
kzDu2L4zNukCqrXHBeUgdJz3KwlmbJDr2/W3kBWFuGudnpqaRpSQno2v20LsjxYC
xueLriYmHlghe37tmhDPcspYFDeDNZuZRVnjFoABY0Kq19LnCcOU+JtakwFpMDAp
b0nmwkTaNhv35MVDxflRXJZH9Bw4vY40jlvTsf+QVY6WGxO2swMudRw77Q3WiWWT
3zD4/ojIyfq7Fy+Ir+JHoD5i0Vf+khsOtRmzFR1dGyU10hCAq5qgWFXv4O7cxXvz
AmgTjjtxbG5Oy+VyAVi+zzvAWvGoVwEO8/cn8Czjpe/Ar/a3zXn4dFvLit7L4ZxS
7Oq5eDRA7n0okPv8n7OeozMef+0BR4EZypJ2M4oNWxZkfbUqpto91cEx3MtckR1H
aaeq2R4WnVGteFrg9UftMQ8VHOxou7mL2qjWrTIfjN1Cd47WkmWfXHFCywxx4hvX
L91TQC+OT4tYFeTYEhuxbvI3y7hEH7InwCzrpsxTMt1cuJF78Y4F462JPMk9pEXh
cG4OmYd/LhYy8bDF+JoRCNXqrgh1a3QawR5bCdcjrNqgmTTuw1T/iUTzfIqHUNAw
LqLDeOyCAV0Vv6qiP9B6GXbidH+IR4OCbZFBjYvE2SsGxRKpw4E+QfhkDI4Iu2ZZ
9gOGZdyb0iIwr/SH2D/XfnOxqCB1hQ9EZOIBpZgeBvVhdHFWbdWJRS2Hn03pB7Vj
6ZrhoQRo2c5bBqQNLk/l2sMe5ST2Cxi7QdUqQpUgUYCMQJzwvka7degBJM4HytIn
BZmKyeWS7xT/VDMlJhLIMFtDLMR175C3aPQU+tKsXfW8qIE4Ik/AC6C4Vr8Cnd+C
ovwQQsGhXzK+qEhDijUTLPIm5yBlPQpwt9Tz1lYxaX0SJJogab8C6Tt5SDtow4Jo
kzsmWM+xSSUX+pipr6ucbBlPaaJa7HEJtilhrG1SKuU4BRIMSftN2UlErpxr9jZE
rD6Ydzrft4IUSjS9N1bDs29pvDL5v5IGeQkqec3VOJjQ/LfPFm2aKJkswGu5aZdl
Rwf2bN0wfp98ThxygTV0mwQsVomckAsoZSUAH9Q+gvmApAMy1YSzMROaQ4CasTj/
yckgwrWcYBFMKA69gnZGLfu9QL7m9B7oXxW6Z9L106PdjW8Tri9quiMje6s1OOOD
6xrA2ucXXn+4dys+F+WTaFSf+aXq7c2M4NzWtUwKe0X7L5G2t4AJNdWaVxbkSYI/
BCCoy6RNWjoh/NnP5KslvR3qOKBLKMj2LhoZocA5lNJG6dIOcNUKlJkRtjb/UWqG
Hj+Mx/Fay24Vmz8oaRd9wleaPN8AdvfynUDFY+7gRhakVIM+U0cA3Oyjp7tmkNET
1M+qk8LA4VHzr6bCDDfWhqpi6fwCskB7mUEkUpg+s0mM3KhpmR65qQqKg/j8wGf9
BxZL04kLGZrG3reeRxmKRX4DMK7GQGdbsO2hgYoDgIOVgEh/WQxKb1uPB+KrIeZZ
yBUW7HtfzuebQGUMw/xRypCBluZ0OtvPW32rSwN3Yq8JN4xvIWAvkGEBwz2oy7Zz
bNTuRBhzUzqgI/moANZTqbpV8dMn9q/s+T84rhUV1Jw/yv0CTm5o66OkJzS7cEHc
da+lvFhAzi7I4UOExofiDGzUt7dO6VYJAP4BbLkTSe1CVQUFW8EaqzRzVAEA2x7y
GWl2hMztQ9NtaAXhCzBachB6Fh6e9Mw9Df/CNZCaqAWxjsSb8JnFXYLU49lHuWgo
H9R5hxtPRlNFn5O5zXYDzuZ7+v4IXQpjebxb/9ShA50UVLUiIl754FQ9RaJZ1hwZ
bs9HHsnU1stDeDMuZwSkMkhbR4Hy5UI5Zi4QJN621NYo6ecm1U3GcodHvgbCRfQI
emE1cdWPsJ1nEOd7KHQJk/A5tY17cawDiKYFLjGN+T1Fl6zxzbuimbMk5iWwFRDI
maUV/3sQuGF+8hA7xaWxLC1BOZZwkcToDD628MuxgE2Ll+ZlTVehH9iwKqwJuLc3
OeeFUgyWdg5EtdO3qF34Bz7IuPIsBYGBn8nu4drkqtbwttHhXNVrNuRMcdtDsw4t
2v5WUBPtpxCzS3hZzUyhk5PUTKXS9aDU5kLgxBMpz3Qs0G+TeUFEXsZSNYp2MSyl
ey0HyR2yxR3zTssAZnwXZPlWo9xW5izqAjjlRaXV5n6rm13JRVs0KLs3HBWno6nX
aCXAptnj9Xcw0aiprTCwRk1zK9QI1EYFsYvNKVMdL/XT2epBSM29TJlEzI+u/Mfb
RGlNQi9/nlSmhqblo8Rh+FCdHG5Qg/3Wqn9qvIaFbCXckXC4yPbbCvK/z1Hu9n42
HFamG+0sRxO+TyWMoDZw3738z9Xqm4BdEh6NxqyKlCYyDkrZVcKwbcYzvF8CY6mR
EnaNHLg5w/sNk6Na+tAfRQLFWepmVhSQ5CHFq4XMYHuYw26rrX6ZY+oZBqa77DbN
riSPryZU88btXfG5GQcdjEw1ORY1F2H+GxFWyiyqFl5a+OqUDDfqS11M8FyITg74
Vektc1apZdm92f5+vykZ+7HyD4eP8Czc5IpG0kO8Ku5jnM52CtIW9S24h6GZln9/
sU/ZI5ZOSjMGt6K2zmgEMHo0+TCkrPergDsyfnRYYBNdWqd3YHXYjPRzuhNob63W
D2ddFe6Qa9jutiw6svPEIJcbo0vFatevrIq+NzbxuLKjCxOhGwGQd9THqtfF3Frx
KuUxiqKgNc+N07Z1DH/1a9PjTjdToXxyEDKzR4B+2NoI/TX4mOiiK56Sfszf96jK
UtZBhGLClqjZ6rPTNekg4WvKvCkRdid7KVpI/fPIylwP9RlV9XRjkR40fU9YM0Mx
fKU5Ijx/qF4yhRAR1ESbRZNpWYQUFHQTGhdq63H/SB5pv+CI2M5rMf4hQ85boyw/
ysqNV8BjwgxdwCO/GZdJrjrIoEGnYu8Vxoyqx39jFRMfBXyag3CTQd7RZvh+LkMX
f14TdFJMYAxYjNq1froHicp5w5anGtAV8V/jvjG00r2+UbrpKmuL4uSxMDHXzl6X
YTsVIk438njvZI7ZE1DLoxo0P4W1EbALtSMF4bDKuZ9r4Pt9BLGgzVXzO5mhRqTp
yXnF4UfsgjC1xjgMyJn5qs5DyCbpAGHpjdusdNr91piIRJ6JQf7gP6cEWGndDVVj
2b4zWJYoep4iUMV+Rc7l5typkDDqZGWYEyLeI+PZ20qrCzmusDBCRHWNrZD2rQnK
av6f1C0lLKBfHIJVey6EM6k3JALDVichx0GQwF+Tudrfx4U3Mp9I7bc8BZmdhL/0
nXNT+UoquK83pW/0GZJXYH9wqxDnNf5QHqSWzTSb6wy4uyG57Osx+vZJVdeer28N
uyAEnup5+f4pO7r5UwNlKntbjxJKLfXo2iI8kEK44mo1ME1fccVYafrETTt5KNBo
60Ik2khRj5RHsaq8SSXtnrOjJ1Hph8NI09+/dE6SCliS6xenjKRsMcBpSXhRlzLF
v1M4fUk/YP+Xna+o1q8cPnEKOQZ8wYN5pqmjrUUDE1yMbmmVmwFsTqZGF3yBagPe
524YS3eEWQjKs7lrcZq4uRo6cZjt5sq30XmtYVD7UQadjp/Lp/N6EwC/hkaXezYG
EXy6UMQs0m/nH1AyJY5pWMOX09VEn7Od4Pbn9nqfvNnTEcjmUwAm9p3GPsdFnH0X
YC8ezQ3YQsDLTExns5r7SDkGRslbFrXBrW4+0wnOS0sKeW5Pgn8m4XVxTQAY/E+3
H/lqUWxFZ8QriVWoFuxyE3RnAsEgE/2gYycCgnslw7APjjvRy62MGBYfKWBUfUeC
8seeseWUZttBxAr3ThBn9vKDWq8gYJuv7J7DrMzu2jO1Ti6axOlnIy51TexY0/rh
j40LAET0jEPOZWfMOReIJnZftNdX11+Hz0QO4eNxx7S/3CGNWt3oN/7Jifj15Ooa
eLS6iaf5pOmKSV99CvXsIudQ1uo+KwXkyRZF1d+BVe28fzxkdXMezWSRI6ylkQEl
o4+zwrC3CJFA6l5DSXyOdlY3UrBpoZbzNoqsl+rOlsudJvBLrmIczTKBi5gVBwBg
rSlbOjHSDQKFP5g3s4nxuLS9Q2LtvM/R1yFyj9mpUBbet8919vM9DgkOpv+GXQDO
deNUL55pnpEPvZjm3Fv7wHy9k74MlCqll8Xbw5TKEd9+ecfp3eWS72H/ewqHY6Tt
MRtsWYXQ24eAqLuCc52QT8/+nSV387ynvMGvq7IcNSq701QCr0bcTa6Hr8cg/+l2
ULsGmMFv6iBhVf6JjwiSGQ+BjhKS2j+P/qYfnqilGzkckGXTl+E+J8GRDhJpgcY8
/CbFVuw9lOeqbWHd6Q1Dpu2etjrV/Rva1iyJ3kBGIDIH09nepOtjM/bXN/To3wl4
b+YtOlzYlNE7VfUs74laEPwJUvLpQOCw33k6T8Nz5qKRN6NhM6wniEKm9sWdD0Om
rpFKqmsqDH1CEE5EuZHQuMWVHHZKhsMun+nCcoCV0mh9w/odm3nxbjMYN04Endht
zxNqbRzVUHNc0InYYIISwxnK7T7181ZDGvo1b34mNbZSOwbkhrOMzYtMV7BUvyO9
uf1as+hHZn6odzLXrGeVPv6JeA9jU5yClvePZaV+7uwzfOvKeTQa90U2pqkguZJ9
I9K8BM5yXF4/E9uDweiK/hyFj3WAoMGgdd87CI41BPDXF3+xA4rbGiZERCS1rBeR
dgdobeR1X28hySWSAol7p2AtzDzP4u+HZbqdmYm1Pub4G+5tEDIp4m9ZTVTg7fqf
hfGx+izP4/05wVKObCN6AMxDuKM/bpswzj4duQ7I5JZCAWuQQDUF9k7DdFYQjC3O
cX9u/NcWTzztouEJnwtzWu9HZTDsoZKtcNc6YFRGT7emTs5bP06+VFbicc5hYxxq
TLFX51rBJ/HEAL3/bLN/a90nAVQD/110uVEnm0wR3CTrtbjSwKiYEMeuUcB5CHAF
v30cSgUSJfGIO1xv2u9DanxXHRAQqj0kTYcmKIuYQbKRMPPJlqWn5y8e8bRb4sSb
QaUKbuN6HqVk9h95vCC//+3y+tvET4vIkuPCYEx/2ozKMsIkWUuBg93OZZq+U1Lq
apFPq6jl3RJ7OBf8akGvvHdYBkdSuMkuURlCaF2gbhW4qaJ4Pky7aZGGOPym1uQN
KF46/qMjze7OdcvgH9Ef+xOovaYMZEjHPBM2Ty6eyzZhXkY/SlcwzWUqxPFfX7qD
pyiHYj7bePrmu5IvQyW3Ex/sVuIQ6YllAkp+IKKBF65WuZ4da3hNPwvFv9Y6pUxw
131RFwJjzgQ0jXKrw/pkIjZpc0SJUaPdf4XN8OkbEM2LsEH9pRycQAoQtVTu2Vs4
s2/4X/sypPgZtEu4IzGhwigrXSw0O+/QMQt6Qhg4oXedt/Bu+AcKU4z/YPLtjH/N
Jfv9hD0oRi515Pzwe2hxFAEkGJe3wIqYDc/68fDkJrZKwQzs9SB3FIu47jiXDfVN
TCFEjTWnJMdxhstMMrflENb1V7vgGyjbaJPJ3sTKd2B+OzkD1eI1dEPCK2NySH3U
K9Fz2kdmDoAb392mT0mVZGeaYKQ534bzazlJSMPLy8olO5+e4rHxk8kgRuRWKs2B
1+MyrRto/xa6WfoKDNnxMbaBRRmYonyb728eLD0GtX3MjyxDPs3Ew3A8WUXYQcZg
C4Y2x/DAxUXEa/SMs5ymBZoKkcY/WAJgd/OJbnRXy3aaaEb+hVOH6Z6k9wvykwf9
J0RYFb83ab3weUPv5YQfEPu1HwblXE31y2KkywPxXRcw8CTdaTeYHO10RmMR4Exc
mMlEGU0YtS5VJT3VpsuSq0U+QSZ+wrb/PN5Gzbtf0E0oiCTrJxrT9iNOXZNE1s4C
Filwa0T8CSOvs4sOUDXzy5YR/oAaFVKj8U7GwGZTCxsBE9AbB4/umB/DagninT+T
kZwQTPaY2RoZfPDKqo7VgtFWKsn42WI0r0WJQMJRR8kjayYqIB9N2zSh8OFY81wB
d6C/VsXY35vNsmDO9E96hO+zOv7r1DcU7IJItDTvWTQEN9NMXqDKNon7yYCvq9i1
NxWeT8iUuXabLYoxqgLOldXGjtmkrfW0JNtq2PblGQ+1qAY5Zdjvf6zy3VmNEyEd
FzH1AIFPsJF3w/rwftqpaDYYmSzs3vECIPHduIRwJ84uvsgJK+djaBe3d9QM+Zbk
G97axPYcSPtDCTE6Pe+a6vysHcetSFtUjnG2zBsZ+xLTeAocw3/wCx5KY6zDxIYq
0c7z8jSM2tk+ACHBrdkJl4XpqJSkJSfdKIrWFcw2GuKO1fdXK6UBakhbpB9EaL9Y
jqXKFBp4wHZwQGvcq3Sig7abuUWfoienDpVU4nsj2ODZewUbKCJ5JjNf6OOO5isa
D6kjXCyBboLqexhVTe21kG6oy5s/KHg2OTybgGbLav9lcdYNPbVxuJh7pCdXJZqB
egVgwUpgx+5bV1iEF0HkT+A48FbpK2jMoEx1bq5/98txo29na/7h9eApSJxxpLoD
8ACDss0oDcRp5r0dTW3sj9CrS+35V1lMUqYBNw/nw2aI4z1fOYUqX0Azo0C9ofoP
GCJ218eSE4NI91OVcrH+fsH81hHW6W5J7hDNb1CsWXQ6eCQDNwRTzB1q6tHiViFf
tPJy5GnWs4fzaXZo/I4ac56eEcBimr12dG6wVnyOVHDQHidNiduUrsPQ4bcIJqRh
aBWhjSo01kl+XEGBG8mZAA==
`pragma protect end_protected
