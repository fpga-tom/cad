// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
afT5ykvHI+SGk3JhAJfh+byHjYSVqJO7kDMLr8+elzHrV3GkWvfvCL4479lakvfJ
9ZRcigD00QIDTZvJaTqttbDVG6eilkpsx5pisRLB2I0OqCgEpbu2xrurQVXXtozr
IwRJ7w5iRrVMQ6sJn4T/97rwgoTea8D1iOfpTGTa+HE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11072)
UoyCFEJM/WT72JG8wOI/nAUkUhaAzVhKkr0wni/U1RHCUnd+uNH185dQQ3B38brb
YNIFUTjyZ14IoJv0KgdrOwDzZHZg1TIj3EwSv3VffukO72deYd3lyTJgXF9ApY0J
WdHDxUijlDIkizsJUAPFnmJMc5+jPCmm8sYSEVrHHe8U0gqFa4VFKDqg/8VrCirj
1bBvNReBHqleeNYgBII6YPL04C9EoEe5ifILqBq5aPJmzCLOAshLJ+YKJxrbeEb7
9uaDiaA3NSP1tbBoI9WU2rOubk1VoWz1BTxFJXN9vTLy5HTGSS01y1M7CgIhD8cw
sm3EK/agKtyxQ6asHhSpcvuwSNmx6mXEXJ6RQ++Dk0k/YBj1GnK+3gqUmq8bhSnr
shbyQrC0ac9cnN5C3rpVAmuf4+rjj2ZnaKhYap9rzXyV+TBi29wTzoTxFBIiB6Ma
nWk9heirDS8r8eMDhP+adSK6RluI5f8PPPhaqk6Ga6DlxpLnOoVPAzEtqcuWb8Q8
iuBJaY1Km15lvns0LMnStLpqraIDVxWGou4bS0AkpaGD87LCOUmkU4emQvWVLVX3
f9G2qijTdRKts2tVXKdZjFLugoQ6R1nYeTHNfIvxSg9KRYGErLf+2b52t12uvFX+
A6EyiajzuDvRQde9Qg0zts56k7s9WmRAVB+GiRgtmRz39pkJIiuNBwOf2Jl5O894
5sjFS/F6/U6dpwDgyn8lXPUj5RyJgWVAGhqDTdJGZhf6a8qxkD8zctT25JfJ7uwD
tTyFZ498y6O06jVc1IfFocYQMWUPzb59m+anu1lHd73FXtdmBSbLyroYnsfM2Xkh
DHyx2W11hG6i6h4pH5JBDduQMoHLRB4gdZ2fcohTi35zft9BlgaWK6GY7P6Sl0dn
gY+JJbF3DaW88RVAe/SnWxKA6inLBM24jYbuPeCA5lY8Cr0rOxPuHVXojeFAT/5y
iSkOTCTfHqsOvFOCsNRXexjuXAdigXjNWUriX/DgZ2D3visDPU9N6DQcRlicD4gs
hN2EqNQkYpWeK8NoLBhQAEv/6CnGaV3zN5Hj7w0sXqj8RBOr5tnJac8foikK3LVY
WVHP6jjCHwFSIi6EGD7JEVU6btTPSg/mH/kF95XZ2gHT18wKW5lUWkQbOyoq3fiO
/kAGLZDnG3EYzrEL5YjEc5Lq2yQTx0wC6BR/iLVG2vZNoM0epiv+nQQrUIXYKQ2v
bKdgqx3iVtPIZrN5wxh35z42/FGUDE6XU7cmayljpoFnKFKX78M2hqokWmd6I0G0
UbFKZFIML3zUJdaMcQRA8TJpRC+1Ufozgqs1Qs+y8ZbKNdxKSW8OLm78zZA+/BI5
PH1AeswB+zTaPnFVZwnTdKF1ZbMLRL98AjJmkcKB1KgwE1xgRCKtXbxbSXm9hh68
zguTOMNXwfw1S9YG0g+0A3HUPEJ4qacWm7I7JpV+1UPAOOmNrUEwiEQIiR4hnt8c
due9reUEm2r+L5xerVv1sfl8f7dyspcuuTM7mqsku6o/4qRC4ysmRPNfPxqq2WQ1
HnA/T8Xr0YebiS4TZ9sc2NsfJdDI7Y4zCOmz+OjR3PAELnwQUPASFfHOVugsoDP4
bSYKURqsoAW2Z9cdLLXuuewPwsUPtJMlHWQl4/QuaTnCgYefo5+tDckjz9tDk2O4
ai4ELNsP2OnOTUOzF58LUwfcLlvrw3vdrlMZCexV52ix6vJvC5MUJQZg1UbfuUVg
25rvuCQq+ZrgEbHg5dpMXJFcoYqkeJpbDY/N/R5qE+9dntY39ZEj8sSr3MmLUYM2
QUcdQcImzCSMncyjKcsLOFDU4vd8d0RjYUAV2ipIg0AwThhu0bi7y7Av6V3eWP7x
eaaYRxnwSxJ5JCgESUBnvADfiV9lij0fdVzaHYQ+BiMLZ8i3BbWIpb5om4ursT4G
3niggDG1W/c1H97vEcaBlbzhzubHCWbk/EdZP1vuum8G0klEWsKvXR7Fh7s3r3oF
YaVqbi+OoQLNCfgKMNGWtASCELB/nZv2PBhdO16gBeBWXn9Eyauq3O9FswV7QbvP
T5+aKeqUSlalgCpL4/GxElgwL2tdSi043sN6W6nAZA+mrjaasD8I21vjkIdgS/qw
J1Km2qTOh1yknjs3dVAQZjT4icYu8UFcwlwflZbxhqankq6ee+fszY2DXXbjtMA+
S5yl5d0y8JOUOMG7Gj1NruMIT4cJKkBacWl3/PzlAjXzOUX+wtE3gkCKQ5Sv7sjs
fPoQ11aFjN+zACsVges4fNgwc3tiiRcv2e1Dz9tySJJCJxXr6jFwp+sgRui91vi4
gL4JDS0ABp1Pf7Z6hsjPja25d4GokJhArsoPHfEkRmNIRYI2x0Qh19metWlZkpsg
hfc0N9SOsS0vyNTpn4ZrPoDRffpndx36GqE1v7SeFhNYNcWZZA4FXTijhy3CLq3f
hS2s7yPwIE7Z8G44u6/9HhFrdNs9XylQru/izGXCa3v4XTj5iojOxQ7g49/kxj+5
oH47OKvwIhTNoGJU2crydyX+xnT7rCIt+nX9/G1JX9BiRxh3Dynw6Oc3zpA7YVe6
f8TPIxthBMLsLmqFdqklQD36I6MZAqvatyCqeMQrLeVr+6oyhvoaUVX20HIKilhQ
DotqZbow5I7rB19pSRaKS0IlSUGJNtT80kgU2wV9pPiniVAH9BQN7P3Vn/tDGQUM
jvBW/WayQC8bh9svoyaqzej8HL/lR/C/rzneDwt8cj05hocPFwMuM5lk9yhYEe9p
lZQ5UfjRTahN8mlVhyAhrEpP129R21nQ0cedR8yGENDWpFnuz0rRMvMaGAvOIsGf
6nvX9ECRc61I3CMpXQSuU7zBGjJfxSTBXZU0Y1xyeZQKhmoWqceKpjoWlFq64KqV
fZxlXDtoIfK1k5LWpQQKM7iSxGAtM7PJWF20nYtKrLJl1GJnB+LAeZlfUMUuFuEh
qWRbu9ov0px0wELJaz/WviixBtC2jKbLk22gLP0Jnu6IWrXSJ18FUKin5sFJTtcA
eQWv3bGaeIhepvtfNyO4R7OJQbTHbjp3ggPyi3Mn0ExV8z7x49xuTd/DymVdk7oT
DVgjQaPtxoBjoIEZYfFr/703zgSJCKmT1xTJ6jLgxTXRzPiNIt+AqPxNhGa9Mr+F
fuXWYcnh9vz/X2wMgRcmjvhlpcveh+rTCG2vh5L3CvRrfdhd/X5udHX15gmDZyTE
K+uY7YQmgkyFn6/Z/H0ubxcYtIje/28hOhXQ+zp98rSod6otlwyupFBSxERsPLef
GulG8I0X/ZifJEUqBCcH4Wzw9q5UKj9IdxO/ofpqU34cYnSnZlTiOKS7XgFbBS+V
aWWRi7SvmxUmlggn8d824zubZtPPF5CqDFoWmUTj9In9TFVmh/kIHE8fvcog0LVr
18GPmfwNwButzKuCnOXvb2KAHXKneZqz/mMrzAHyeiPPCfgcgO4IhPS+qLP05lRu
/zIonmb3JIUSMDQ62q672XF0P8hIPqds+/52NQcIhPatgijklgAcseed4S5VkNhV
KTk9Y0zLp0SK7EcRbO8phLHsmSlc46CoelfYY4OLJDEBl1HaGpCMMfCPIUEu+pHe
cGGg+QG2hiAC+37rXUl+XsnPyeiYVel4XK5MOQknHFizh99ohgmSbHJtDcbtOJJx
Ra+vIkoatKFHZEemg39a6wZc5zxoISqkS8DpsaQ/XjvMu8NLXpwl898P9D/ucauS
tIwuBl+/1dd8iQ2vnf1Z6zDHXOEX9iXIl7p3Jxj/GenWxFfhwJopA5KDWLtsnY6y
wZEbnwLMiHAO9RCWuBuJFe7iwLFF09t1+Kb9rmkeVwdA2fQQjO5ca02pBHkZVbK9
O1MLSIGmDBWOZDH2iCdfLfK+WWPx8HuBSnCl0ugDp8g90Km+lMb9cvfBec7vmSPw
warai6uxPCi64sqeFPV9zonFJPBqvSaiK/a4V5LT9fArvdB7OYljTELjGoYnPWIT
Aiczua9zY4R9umvbAnLPth+TYSee3BvZT5EDORIKtAC/kbdWnIdZTJgup7W7xidW
jVssfTzE0ho2ytyBuslonUlnPo43iUsGrwCD8eWkfiXBjZelvoosXOPSHZPu6aRo
C9FxbIrzs4Rj88vf0Iv8vNHBuxGl8W0VHcZTMvVHJUbq7rZkmumslY7g3sR+GxcH
+PrVx3YEy72U6fkK6jwizx/60weWeezK4am4DA/5Dfw0emMoEsyIx43HM2536/vh
kxFfkCrikxm2DvA2cOT8r1OOAeIeni0uyORvmk+lkq6B5hYSS32AcQ+qNhREA51H
g7hxehZIesEc6Hvocey5pS+xoDNfOkm9dCWhWnEbGM/gnuPqGOze7s2kLfifOLSJ
Cgv/bR4G+GYw+K9fEKzpF07wwyAzgZ+hz6vdVBzCSMiMpmCEaPWLtDSLzLucaTnP
ll1CoAnhv7L0nRpHKBBMTf7kf6gu+GdjqNcxAve1eKhIvOCpUAdrzVHuCRyX9+/S
c2cTQbMV6np3uW5cdFgqAnJx0Cc3uAcT9ekhMlFtWTY/FlUQ6BpaGLiUZ6GI97w+
zIC7amGaU++rR+iaBXtDb/SUoZjh2tJ2ucxHc7ypT1y5CjJxV7cX4tho82Di2qrw
DlUh6R30Rvpbo0EX/J6BGbxSVz4Tm8iFn9qlqk3+Cqp4RLcRHqrk/V8Xt4Fc9xzQ
wbkmK4EzhW+o+72ENYCWwHR0QD34dWCvNSbQ/VT29IgHG2LCmWPoj9RyHSa8cBu5
WR3Eok46tcStA7/WBRV2H8/fm214U2mltlvQDZS3Og7e1iVLuZvPPcanPanZ0rru
fHQ0dpxhoiAdqngfLR2IhRk17G41i3WjVvF7koujRQxM0xvkZAfGE66fIrd7y67n
qkImqbqCopnYyEgZ3aifN8FFvRW9xslryGRBX3rJ2ru8e6QGpDbP7bDsmgE3jA5/
8zLzIywb0A9bvqhyfyKGlunVRgfVWf1Zdvk7RDlIZTK6uILUC0vkOlolB0/mE6wM
6RWA1xYs4B51CeDwXb79/iwpiuNY52gqCDq3+k3Ab5bfvCYAHxLCuWPcFrZ9kvwc
VJ+qmbT2EVTKCj9PHo+72ctzhyiE3HkesALamXsWcPZF9TWMmnU6v6Zn2qalWtPo
SS05iYJ23kv5bYJnAdRn9MaoeY0nmdr038VvnQPLZFPnbexc+rWZS3WO8acHHxC/
l/KAQBfaRZwx2EMnVkHl6TR6KpOnPsalWlC+/tydmu3Eimjqv/zTA0n7sC75z9zD
Vq8pgMv/hymFuy5eAW7vBd2IpuTgjWjeaCBgj81IOMINfy226T4kCrNg8+IkpM0n
mYagrycggEG6dZoIGB8TUNAI6Y90nEuZZ14k5IWiak+/61E/WI9gK1XDP/t6ALiA
QvNd1JCLVRcU1dLuyhza6yzFvegwt/Zb3DWCxib/dU7H4g3lQJ9EqCC2KGc7C80r
qTAs8I99XZiIQ5Ak52WsUkj7TbTUKg2omaMlo3Jv6IkQD4+6ifZuqbW6wmEMehYs
nbddrczv61bBsYw/S9MUM+EPTYslKRq3H0z7lqD6GpsmThsLfnZ/ul1S2TnX+BLf
vaXrAWGdKjVNkGFnVcWNwDXht0CS2fVHModr/jP5nPmecSsy/MPt1ERkD1fpdGgq
w/mYcK4xl+aPyfaxPjQ86CWc83Ag+3Bj4I7Q9s680F4aeXGL3snU3wu6LtsnAD6X
7Y4dWYDzj0fMZ9FCPpvXrVg4tgLH/Aua5hdcIjqFPdllRD4vf+lipYrJhTjIbNaT
2CLITRoAI/orEDXRNB2SZzevw8HG7qFlCR8ScMtahpmAxShdI53cA8Rspj+Qx8tz
e/pYV+EQ0qNWJpI+Xyt48F1tdvaQDIF5Px6q2J94Pcz34/OhsUj7rBHCd8UIqrbR
9Bz89pynz+j0b2aHCW4pZD+tXuHTDjr4hwDQCm8d8xMu6HGS3OMGU+e/EGUz01x0
fzEub5iMHBQh1/y97V7PxqbT8evppUBeyykj6YXciB10/DPDhgnrou2M7BMjUbZ4
iPg5rS+U8aIBWLBF/VLbsbW7r/dtjTpaERnm7AFyHfGWFfnoVmdjdV3dgBO8qxxL
DHCPJUtpITTyoctpqTQ+o24JUez+zTJdkK+x7FzUPA5IwRSoUARo8tjhCccN+3rc
GpVIG27o2AxNI3np0sA93gDFX91+n6JW8d8kzXXCjePfu3nEU3M5lCW1Nl1/rpV7
rNRoFPPHYva6ISqzhoKmfeSXNDz07AGJ3AjOEihhT6QkH4SV+kQ7B4Z6fdjSSFhm
NwEfarKsqAZCLA+xxLCE+5PKKvacXuarFsNyqGXlC95DtskTZ6HV4p3uQABr3Vrz
kr6nGVnq7tPV8R/6Qla2AD0qNVP1WqJg84Uid1f48WpbnlvXiEW3iMnlDPnk0ps5
mRtX0+dq0KAYawAeypPEyi8SFGjMa3JpuGHph5Ahkws3O6xdQWOleovwraNIcX7e
6mQ+qeo+HVnWeEQXNIXHGb3gHV+QSwXbcFU9wI+IAjR5++1p/CD1iUPIoKK8aQiB
cNl2M/MP+ieyEXiTKwTTl3N5OKqszp5YVj14JD4ieEKgCXnkD7cMC0h+jbw/d2N4
2AtRrzgZh4Eop3FAsg3acoGujQ8k8K/pAi/7zwQmupoP7r2BAKbYDj19HqfITAo2
ioAUdX7aPJ0klnuuv4O1nxTy5RDQqVG16HsrqSdlvz/ie/KJt4UxgZfhMSYu0lbt
UNbYLBduG6rwSanlrOBNZwgVc95Ge70OwqZ+9Sj5ZSEYoHURrajSVK9Ukk0uSIvB
2twJmhC6/8DuxVdDX4Zvcb9iddW8LerPVwL/FqmFH5xNtzMhNE4mL+wqsOrMRARw
AuJwD/ItukI7Mo9egXULTVZzUO/KNj6i1sOFs/c4YibwVXogcve4Yjrsb6kxw1q3
xUqKv1IImMxmovkwhdh1UrXlIqWDEU0Lh0y5+wHzPbWnXPPT9qevanPPckNqVRxQ
hH1msr1xcuCqmtpMb3dZWCW1Iqkm2X2ySnybdmzf6d5YBDuYB1loS3r9ybBek0M0
Xzu+Wrhf3gaTTFrX4G/9m+cU7+3b+uDSUlsNVAelM+QsqQha+c+z/GJpTdPOTpU4
gwbuxuZIlf4RCzqsT9R1o/YkmCG1yqfEtPaeR8YiRGCzLiUeWeLAO1ID+eY936oq
KVTaFcYpk7aIul6jgb42uIgxM2Ve1JxBGrK6AD29MMzi3Cmq9KgecREzi7/Mi1jN
xZlVdYFG/ndRrzJ186RqOtywS4shIPWaqUXkXxA+Zv+g9SNU1AgFVtmnop/DKse0
MSX5cDEIZlNg2hTQIM1yfK/u7+0T0MPAsKeSe4Z3//nlvw0CtA477H+WUkcWvnl3
2Pu0bKSv9yduuMQoH9H1bjGoEFIEbBjMp5SttQBrshhlbYODZ+zNP7ly7hQdHslO
5vQXui1DoKiR4sIMLFhfbZUQsFyBciJj1E4jbn31mAQ8PQn1o6DJ246a4Vb536ZO
8+AG+lPATPqCdKCt0ScXBvpbpNALEAfIvpaBBAWckgCy4/rLb+RmZHqdcAyfvorn
mkBlvBrqNfMEh8dEMX+LUHRheraMkQrMhQ5+57o8mHiOo8U8YgHoh38Vh7pKRdKQ
ILxZmdmgPauFEBajrZ00x9wTOQ63i4butFzVX0ubla6eXImRnLisugkLynjaDVD9
6T9L1g3donp4cTnJhrMNdMFaKEitYM2HqSkQnZeWNj9+HFFAzYfKjhXKc8RI1rax
9zTNX4gWoHDtlJx527nptG1GShjNkk74eYxl266J1/5GWbLiKJNZU8fkBUdOqzt7
5VENJK5Rpw+Ee9IV4BTdeB3UIlpJpGdQQ9YTp5qS2rOUihCuIZRnx07ewhlm79bl
5/KYuXpTFFgFRGR8spB3SBHKkNbPl2vjmo6pLPtGOAVFNJTKe6Rr/CsrAQo+GhBi
7U1lqXlKWvSIuApl6tca8EXHJpvsF3N7JfVuVSkJpWKfvSQJcN3VwEUATRHH5UVC
49ymG22dU5fHdDjjp4fxgAc8Cu4iHJB/px2aOZtBVXPZklsV/gaH0pEoTVL2WlGW
OrZS77gAgh7GCGg0vDXHQLjo0+5QkLV+3eEyenivE08sFvgWH48VXE6f7xs1eXOS
mJUTpi/1iXMFbftM5Cv8tpUHgq/llMaGYnMwIU+oQnOoKl6vYoU5SrtQxinEZ3JI
VR2leeXXSmjgCMC8eyqwWzdS28sptgQq6p46TYPifVzfYvTuWIzBS4RIBvsDpuUJ
2TmOqq4AVh0mGWkbfZtm+z9qplX2xUfgKAJW7TJr1sVjCGevv9uaz87X5oE+6TVa
/CgnnPFpnK9haOvghikPgUVeGomgkV4ew7tlB+6WqXLuFyNJH/jRvj9t2n+FdYbx
S0ju0C/+1E/BupFUzdYs6DvmKhU8PxcTEidp0dAtr7adGILcz3YNmwDfHq4whmn3
Osca7C/a3PG9BEOzUtrIE2dap118nWLFfdUWuI9QbKRnOZB17AQktXR3i6sImXvO
dnuMtggughGlvEXg/i6rdTeKWN37FIJama1SxLtFlq9LSXCV29chla0Yck/repzW
lrP/jWC3VvcgBzzCi1UMX8WU6zzvj2OJf85/RawufyQ6VnkafM7IpjhbJx5U50cO
HVvOxu1efXJ3LNO5GluzdD83m7NbEoJvQ8kZS3KqPe2di0CNSOv6v+RPUxy/nfEw
IRXAfrfH+VkHjaUiTTcyd55OyjFi3SyE7egT88VVMgI6OA+trSm5YYtgZA7YJrV3
QtV0y5zHC3MHWbFMBzuKud1RgFozQtB2to5+iZlUHGtmwkhW564ZC7VIAFNBn60w
C4s/8H9GU33G1OIgKlFUyl5Wd2gy7Qt1xi1ZTF8ZcfmJkAPQNeKA/0rZzVTxWnOj
y2JWvpRJ2F54sgSn5jVRD+PbjrlDBetomPPWYov1IZqtpmtZuqrdOUJY2dpPuJLd
2jNenxXKPKXXFjh6XXZRyxO179EsYl/UbRwguPTxbgl1/YdWHt5aPwOYA9SbZ8in
l/FzYpMvCQfm51kgZbcZ9isnZlvk3qGtNRrNto8dEpkSGrvyUi2EEYxzF7CqE6Jd
M686Uc0WNJyjCnDqLJs8qQXMs68l+hKRU60kb3B0EmkSLeyogCPndJotVQqQbTMg
C/5lw8ZoUL7blbDar9l9QuUuDxv0s2srtZ4Bs860kppe62r3IzsluaIZps87C6yQ
7s/z1PxrRphOzSwbpvefa+4TA0vC/a4bE9VcDS3GHK/x8B/HjOzgU7npzIpG9EH0
sANPCjye7ZDePOcQvP/50tv0zOYUde7782RW95cFzqnebdBUbdV98zsncd6T4KyH
aW7N81d8lZ/2cgsl/Gcto0ruhMAmZUBRO9HsTzWP6xnuK3kt00RuqfqfTFjY40R0
2ZujOvCRIaEn+IeMJ2Rb3yf6ezYDng5/hKuy6BTqBhTk2bNaLdwDzGIV8S6i4s+/
wGwKXOB8A5/JzvcPVBLQN9JiS6RMI8ZOtO6h9BAmeS9B06dKxsLPcY4x02esKLCV
DoqQabsN+H73QnLBjdXN5ZoKLWTsu/z3E8M4BJ+70soF3xsU3EWt6DGlXEJnchSl
JagCYeyrs+mDIR+M4CidiAy1VxxjR0nGM7PExxP0BQAHptjrf0S2OM1mDJG1ewF5
qy6QJic33DwlzZDzpstgNMqKfDDOBCJyJ5udKsVISd6/fENmGen+ZeAlb3769zfN
arExB5oYAKfN2r67oMTeJCf7cSE/+pvhPf25OETKQNCN4jQfv+02Ap/D5sTXKwxn
5yM4Z0TJRe1d4RdHACdkTdjDMpxsn6sFzp5lIqj0yI/R/Bppy1LeqdR9OcbAm6bt
hIVJ2By2ZN7xzbxukqv4Kv9KbMhl8qrDdjG1dxE9eeBo48B/CdzKXx+ADPrAPgq6
lpDY91usLsqk5f+4CNZ9yGxqKy4FxhWLyZmSHK3goIIKp0aIEI7U0F+KjuCmTEPl
CAvApR+VqXhxNEUnG9zxlQcrutvFeD9n9FC7E7yvph/1Has7Drqd2QRhV2NbadKH
Wkl1aPChGCkjqqzqwzoyaxit0DtS8f0uaCGYUrCKzXe+ho7P05QflEZDVp1rQriI
vnARdnhHAF4ke6zkPTTiESa2wrADkhiabxk58PZFA5mq/92FZp48ZNCwfHzZODzc
4yjyknOe31KvH+rLBIpvld5LplWiUT3mBWx3YqEWBEsxerkFhcw6z1K0jswTXGYb
Y9cZCk5pFHbw7IgMLkVMBIxmsKcsZhBcv3UCUnOIqV/YIB/DpXPcc77c6AbcVuI4
CVsRg2EB8yWixA1/C9vq2qEU7sS4wcguiApa3K3JsA9/gt3VGcCpPgoXVIiqbxJH
hOVbjYdm9ZpRqiPPc9uUpajheWoHK4+FnlbCBdRscgRx8QSF/Uf076u0tRO3qIHm
M2CdbfOyvN5LHVpHJ6DvHt8x7FqmPYoYwoIfA3L432GP7PGVsXAAqAaeHFgIi03y
9cIbLg2o+IENtTphRSEplBs64apmLEcbHa+LBOojyVTKUPHbet/SCHQB3X+sqKsl
mes7cxuls4mD8Dh0MiMy5HnvSkTmh/K3QBB+yDPoySPabLR9t7j5di4GMztitIJs
FSKKECCdhV53qhNTHzWYEED2ia8MoUaCpdRfFxAxfwi+A4auaewLI2as4lVY3Gee
w4bButxo5pRGC/YbONb8mf2VA/FRw8mDUuI3+32jf0QIILZK4DpdNSWOyYzp3apx
mTiJ+odbct/zOqA0yPkd+78y5rzFUwPLr1d6T4GgxOgfSOoUj+xf0kaFZtUAluwC
GF5cKa494xfPnVTcr9k5mjCtXy2sTtC8VObs61x1RCYBcxWcdcw8pGHAyaUe1IXw
ZotHhxEV3WKGzieoPbOSfEf9iNfVEOHuk7fmTbV/RLtp0mZNEHE1Dzyqbyjn6YsM
tbL4AijARp7bohPtbFcfhHVlXOkRHJH0CN5YSl1t5NatMexmJWhhXAiYjwlWPwDM
K0vf3UomedqapyqSInAhcU4dNKEKxswijT4IcaNktO2KcUB9RI7rLWAvo6VCsJcZ
ky0rYd7FPfKkUgMY8Exzq0t4U9ywkRuSjVwwW/wPz0s6MOlw/TUn2s7AaIQrGP4J
HdXbS7UjtZr89De3EI1sWmlSnLAZ0+1HiL1i7/uDqL2yRTM4HXptTTWXj6TUGQba
TT9c3fhKVr/06fYfBzm+hMECiuRgcz9Tca1dEmgu6uR7OXZQDrN9FOelfrd87mdK
Gf0Gy2ZVye2o9zponQPRxg0AOIccK8naiMOXZ/kaxfhELI0ogArBqvs25Mgf7Ohs
4g6Vtd5QD+hn+lA/2f5EvxtBDzFHmXFZtbKfbIFB+xIbfHf+gJPRLkLfCdWOxvze
q26aWZ/ZoIg8rqUjj0RQYyVRLzT8L/EebY09S+qLhjDfdiKQBxoKl4GR3b/sc7H4
dxxXZvfdKHg6836wi0Gi6BklZFigsQiE6tMrgNXMDh5BUf+irgDwJZ8PWDiE3dSI
GmZHGl07m5pbx/BELJrXhWjGezqnJF2+B/0VXu5JBNYFbgoRIJ3vWc5nSBRunytJ
0n8IKfReR7ML01X5SckvfJtjdMwWZscHYLLWnWI86SdBOdKWfK4ix5+THozJfXfu
CVuHfDwyyuXqxyzBFByAev62jb/h+YNkVgfF9MzwM90K6h6a5PZeSrZfuIulN93G
PU35r4yaAdc7hS1VReBT2N3I60uWnZkjzPm8WyzaHkwrVA9VUSZy8tSP9ZW5mz2R
e19Y/suKnGDQp8StI94H1a4p2f7Frn8r2NMqBpH6V9Fviv3/L3ZnpNHWssmsSMa+
3WVDXJvdTgYbQ2mgvl7A9p3xjX1nj6VSinTBBcGazJFbZvyMyfon68OQp4Vs9zUC
tYgsnqJCQ6FtTXpPYJQ/Cl4mFMi77hpkCH1bTEQ4yL4d/iJtR7QTErvZuQ0pSbP8
h/Wnd+D33IGIsMITCgab6Dc5YyB0/fF636yO0f5NLmD0tLytN61IryIy31I+bSQy
mo49IYgA2HTdm6GWlXhEuQErbulJUJIulpQk+OZ1eXxTEU2jSuSj4SEXIVzW8+E6
HQ2jr+Qxjoar0hKs8T5UjQ/79yP/Oexc8mGhdLDDfs+710mdBcv9MPgyHynQ5Fuc
HVQcdaB1ChDmffMZHEp8wTyLZKT1u4Mq17rNg41b9Y7RQvOnmOQqmbLTbDsbN0iv
yXzteohWPLV/YB1rYoFvGL7c5WIxA9GEVfQ6W2beaE8QHUcIPLU5fck/Em6IERrs
dUfrmwgj33f8jwQqkPb7Dnv9FBrekTCxgtW1+RpdJhcZng7P+cMtJDZ5+wcgki7b
/p9rcm3b7mnPZczb+M02zxNbUemT6gb25RfltQznik2OmozIYATAaAbfqQNd/pYv
We1kFzIJ3vaEb0liUFSPJS3/oRU3Wpl8Vj4eaStGFmv4+PXkvj8/PjIDCO5TaEpu
hjbvkzTAvq/0ewRItmDNBUSo0KaI6fa7sLtQpgCWmMsEOIOKI7MqwOLqCws48LIA
nzQbZvMZrb1pkvcCUlg1RpJBzPtqS+z6NUuZj4gbKsrwVDGyLFx+/ypop/2m3GUU
EJ2vK2QpJKtauhLC3ISPn2+0e7vfFNsBovT0nHKjywM1tywqwAhYPlAKFOnmXnF1
wpgdTPVJV6bxbRHm63EAxrCyAhzo+28pdj0y4WAi/MTe9eBhM1c/4ctd8kLApoza
ERq667HZ66vuXSffwRvKkEgJi+hZAkM4IqUK7RhSUWrRdfCKGEIb2EIu/EiPVT20
CLGClbym8eWNXGAnaxQ8RdsTlmB6THywb6Z4IYXea1Iw4uwL/OR92dbbBRcSvB5M
Vmcw7aokDl5UeUfKP9/0Vf/Bl2/lbNFVgXcWNklga344cZ2QjfHu1wfXyovBpzG1
Qb9ltGjUYigEEM/Mi3UaPUvLOWJi93brODyKFXbO482mMJh3TDW5AOwoTUWR9M7u
ojJaloVFnqaF/aEzZGOieqLOxqGNYpUaFb4mi7JkUF7mBYFnBGn38oSWMxw3ismz
dqUyMy7ZH9dsUZ8GW2vP4QgMZByKMmtCSjAoikkOO3JDeO4ZgaF6jZKPzZle4aF5
QBci1cM4GdNjymUhchKUwwJxsSYYOBBt7DMkPa5YNC3tkxd189VvU2YOswhpUcqG
0tAHw4faJxDVnN2bZ9U4DrZkzF6YAA/2kWZpzrp7buqgUL/fReMWl/38mmoTTE7Q
2kyAk4Mr6Y9vUIiCRXymo/WRpCbONs+Cw+kBR9D9QthDLm16yGnuxZgKbGPXh/e0
DZP6996n8rx+CePsj40PZREjqvPNx3Dvd6tOg1jx6Zx3K60008nZcNc5i2rHIHSo
zUfzTO+9747SeP4fvdDf6TQrs9V9ZirB2mtS7eLP+kvOwzkmsqepD1p887U6bb5q
ui/aMpmTugN79n45MUe7xy1ZzsP19nwEzo4KF8nZRuZ3W6QEfQwmKN5caSz8LiVv
5A/uhtVzOuO+4H7PYkdmBbX0chX1i+faY0YGYDX3XpvJc4xDtc+NoLXjNfBWHyjn
yJ/POP9q77er618/WwMIet42I0Y5P9RuGwMx0f1vqfkAGqX5qEn4J1MEaMy9qF2O
y4DQYV5MUJWgHH/4GaW44Q6ClHyf0zN52WFty5NBd6U4wBKl72wfks9c1MFNjzQQ
hNgpX7AHXB3PpwFC/VVffnvADGYK9aH+LPDLEWmDg6auAp8xBuCukXtb8fwlOH15
viWi0VU1ZME5/+uYuGOmVssHmAb+UwFflzrhNDU34yD9NWFPIgCqYs657hKgD4Wg
YGMV6lZGT+8qzgsyd7yMfI8GxIcGQ2hDECXXVo/SdoKFfabmcd7aqruepRs8ODaF
gbxz11hmgoAOIo8BFu1wPScrAUq6OtUqonBV2Q+dFScp4wgRvC3/t4JTA64zYRq9
teICAiNJWUaya1mZnLlLj5tUKfgXoweaI+7fl+QjTj326A0IeQBfy9Xm9nwxDlAe
l8nnWXtd8ehR7ToCrdl1neVRQCcDSD0BrWMdt3Cjszz5QMv1q76h5RWi7zD5Hpvn
kmbSIEXhhCHM0GwILSKf8XCpKZwpua91Jp5hjBW2+VXaoQ4SST5LEsH9VtwPXb1q
FduZ27ijuykU8lr1Bwk7iIprzfYxVcav9BLPqdNmToXPd1MzJDQ2zkq7+Jkonfcr
RxMWH6SFVWUcKD7a0BZvdcz6a5WNUeXJ1QkuW14paMe9U8fyEh7w6+WAARvIbwIT
2PADgj6Cdyp6FlakIW539iyU03lwcAbiqOUTZl2fEnBZ2zHmZFDMpC14DHY0OjvA
Ye7ZOdV3o6PiUNeO0HQQs6bfeXRVqjiGkjrN1Pcme6vXfL31sq9kBZzwDjOdZoWI
Ao409IXHhqxIFqD/34klNq3Yq0N5d4t8ikjcH7xDF4c7lE5hV1JS1tYvyfn3GQNq
v1gojpLONTELgdKjjNTBOkrqndfk+B4BtyjhrnP5gZZF83Z1h4aIGtjivYGkH16X
FDlUPErnHLm/kF8n6zqeEJEYho/hQJxYiBj6zxGfdbjD7XF4rM5z2UcGUR4F1L0V
MnW8v2ZfCnH5VQAWT+xfx8R/Xjao/dt/UiyLHngrqkQeGVxSv3jsmZazsUm+cvfP
6sdm4JKql+yxzqbkOlEPgRnKIgksHf2KAFuzIbye2lSXkjTW0ter/tS1f553Cdas
S7jzCJ6EXvldkLruP3M/1JoagA9aDh22AJrlNiynx/I=
`pragma protect end_protected
