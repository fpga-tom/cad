// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jiMAZgf0JaYsa76mx6HvOLn3UYYWq1Gz9p57dV0FohXqRXj2jLWlyvNiLSLrdVfY
d/DD201fRNld5jYqk8ZNKmG6uUNzlqlNdoSm4kPatBg2BUXyp8QnG2AAAZMrdr+r
5kQsrxvqrG8xBPOscFbNVqpkM7CcxvaI15tKIXIpzrs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7376)
nJHXd/G79G8SHvVJMlWrCR8Va3ddw1t4Noa4f0cZaPX+UeP5LQJZ2FK8qxjXdthy
l4vIYgHugsUIh81J4ZWSDUIcr5raDEuHykcmpnL9TABSgOJGO6UZO681fjsoMHpc
WnQAmCk1gDY0qTdH3y56uuEbtuaEUPfj1b1r4NHPyCGZbns6w/sbp8Q7HlSxqI5Y
DMqHlAyFEbvnF3VpndldjiwZXWoMhoYsRFyiKRRU74xCKwkDj5cpovbBCCz+etdB
/5gMtAtoL/xu0M/JYa0NXxdlq43KzMyt/JU9ajpnWDo9f5l340HfgF4b6HMNT1xd
Z1oJSWzRQhmfWUEJkf0Tj55d6iXaPyAkYTYX/23tV/3xolbyhnSKY7/jgpZscddX
AAP8IBk4G24i3GdsmMwXVVovPW25ubzUqbTUbVqML0aJLaJdCVUyMs30LZp0v96M
0iH/lAeTsmb6tKdFuVjhv2UP1M5I/F53T5ZId8pk2bXN0XilyJl6EEtHEqtFs9Mj
TiegZFcVqdto2Lvrr9esszuxvukAvlEgksCwBvgtzK90IADxW9XnTIQRX6tE6nR/
rlIzMVrAlXrffjdJnf9A3+F0Kvobz80Sw55ts41MLFriY+C42WP1C62zcuFyfk2D
ysllhjvzQkFZh04naH7p3UacYw5jqtx7FYPWK/85WR2lK9t26b1a1SsfWGcBrZio
0VdZ49fYYOwfPRgBTAxyAjJe7i38sLlYwToSlecHbWnha6LsFq1w112HeJqQWR0d
Mn+za0sUo13VmOcT4lZdrLH+UL9kffWEnQ5Mj24ImXQCXT9WlxpwbCBoYEGhGT/4
7AAcb/vXzpI8wbh8AzmkfXwUXJvTV6mT4uScRwgEHzX4a8s+BsmQIqgpNOMjEAnd
NvP+1ihCtRCIQPXgFg5BitAl6bEa8bmSkGFJdqemIs9ZtkrqVs+tPKiYpdUBFZUj
R2KWBtGFxEfcXUBvjfCwcBcurAwlw7gTn/iohqqGX9DJaWoEWn0v+ditFS5pt/Ss
gaIJ18pZv1XsPeEEF8ghlM4CjE86H6G+lEi4Tsr4AUeFae8VOx3A9D8oejQtyV4q
vJk2/4wroUoK6ZHrIfcN91D+gjRUMrftU8AyVZOJGInE0NEO6ljy6LfVMd7+Kg9H
TTbIrsWr2hKhFCmkvj55LftMinw8z7IHGsrII7oxKJhIBwiQlDJR1BWwhYXbv0GB
iHzG7YYo14ao82rCAGzzPT6RW5S4lTYLvFR+D9rohxfrp3VRwumSkzz8/hEUkxAy
G+cxbMRdZf9ZrqrKSO0Z1D71p70E+v8orlWk0wmytqw9J5vgyREQ8M8BwDBwxx7B
e29wzr6SyXWX/B26C/93GXSDk0BrTKqQwPeD93+Fad5uPmEuEKMWS2GWDIG5ahTr
sOPLTJ+juYz55bQXD6+JimEIS4Rmx7qGLoMxirZhOkDYvSs2rlv8kfEanROVrdes
b4xpknNWLBO2SKZNeuJnfY7AK1iWcJx39xdYeua38Zex1S3NiVPQBeAEpsKnQBe3
6PutsNx78PY7cIF2HcHjHVFqDWQpaprZpKfVZgjh0V2xuCT0kOdYOc5PreHX4bmh
U740CQPEkjZMEP2XaGXSXePVI4Xr6t/hA0R5W/p8gnQ4I+Dh77Cl+DvTaP0QgfLM
pVqM2pYJTR0gb6mLaxmDAo144wW5QnKrflfMMJ7l82n+SZ02d5sfrM2DLIw5Kqk5
8jSw7EBSwNvzaRKfKgOvLfvHsm1ncmXxOB5GmLf9ksek9YYf9iPFOUbY/U5I7H15
NOntvmdFMBXo8GrTE9ogAMbYtjFpQLjocOE1xnmlQvhvA2/zPRZkMlkSbcdrWcxd
1TIbXs8c1vtQtzWN9HFy0ZB/1G1+V9QH0R53dh8sXsdyoxTNIs5MciNjCSdlv72I
q/RPEwcVfWOd/7au9ggfcSGi3O08a2ataai+Le7wFIB1fauC25L6nc5iJ6oKOc7l
nAQ/V28bXX0BwqWSBhk6ilDDTaYBr5mJox/y23zNtV6f+gTFh77xybYlG0pi49QI
GvkeaN3JWv4Y5ekCoMRiH42LYufB9f9Up87T/964u6Mnd+bPTbyl5EeB6JQlZJbA
gON6RYX6fHJXcKAkJozKNTn+R7kE06GgMfDxOMYx00/koDGvRFerG5VYkPbAVJzT
7FUQ/7LZjE9I6Ad0xpRTnoQpdELYHVh3TwhsqCW8vgNkNw0fpKssqIWEKz0h8i2n
YHOa2tWP2GG2GkqLQ4yiqnpHzJ2iCC40LetQOp4T6dhcAS4OJg0RDu5M4x3CJ096
lX7gLmVt/XMf6hixJ5G7q+/nqGY4kXIogTPltvPsNNKntqT6a7gjEiHdXCHWN8Kc
shT4Znwqh70Udtu5ML0PaHa541WahFAC/qMd8sDCWqYsF2Uwerj/nJ10srStOKXr
8eNMhQHMODRvuIjOywt3Qu/lJal5AgmAxSp56o9BkP9gShPVAc+ibJwCabnSZWd8
lvN7OxI6BBsQKxKsika6W66qFoTFdzo/IPiKLKqVSSgAPM5a9BeLFdD2WlkKlRUL
J1y2aBiWpvbIlwikoS5cSyCaOqIueR2R/bWuYuxKXc/Gwaj4nhSBNZqk5BLQeU2k
lJBNS8ywlpVHYC6WYMvbVI/+68ohK81Iqq5ougrHk0GCGxRMrYU1dP4nBOenBlrb
Lb/ulVqIsw+bmuUJI6ANJsxwoKB/ka9dIYXH/jnjYy+GUnfejbL9dnwKjmkzbQ6F
OdUrbZXyvFnVSGRiEhJhlmQBrS4mkvg6+h0+tlkqRmfT5P+vKMsaL23nIl1rciTf
0EZEJSxaQYx0WAvmQW2hfLRZeEWNRA7z2ex8PK4N9gaKxMFBcCBEDu7ETktIBJbv
nPKtGrbIWjcUka2j0e392lnkWvM3a82vQhwxI/IRIT4oIAJ32x/rMdprzMBFhImF
bTVQtTo9+QLMQmYiIeqAY1GyTvfm6T9IAknZOaX2tTYL9dvURaaKPAUV0RYAwndB
mhmEVEuN1fhN/EKg5AOkh0O3/A6hQu0vp/koi40W35iRxP3gvQXND11IbR/a7PvJ
0+5ZK9wD+ZtB9AGbK1/A9mxTbhtDFJ/U5iraPz7K8AVcBTl46jTbNMrOZbj2skGZ
C1sz5qvm1Gmia10n1S9frSWDBR7hRfv7LMPGW0a37lUqK/yv+5pOTRl8ZerUI1Ux
eamG3aaIrtdCVaBxwIgEj8DNthNeXQG2HORVld2Ro3dRlBXpNToz8QbhDgWwv6NC
r+oF9kWklwUqr56F6LlfBVtyX4y8zKl5p8sONFK1UZHvlN+DYY2N4f9mMxhIJYxk
0cCAM9VcuaoomZRkZG+k769ep4gXXPDxt3J46DMMrNhopht3SnYHUJ8e5RsNtju6
ZWtfFsroMJRCIXOxF+RC+h3LdXl8B4VR6nWG6WRbwUN09WW7DpHV1MI1A0vsvNcl
bkzAwRmRcDxRcxBO3ffJP3s2IUNQSU4lM1KNX/gJyuCooXtHrHnIvgZ0PuT1OzzA
wR+nthEA7Wd2MgyqhyaIJRH0/csIV2bsiGifiOa2ZT7nV37SDx15DIG6I5ZwOBjI
aHMjOUYa00dFteN8XU5lVAnyUp5tAwmewpN0nuDMOJhy0j1maZQDuJO8n9DGKZyX
aC1EV1qwo8cKsizRN+2S4GT02lYCzQ3LVJ/24CNsw1k3oOnFtKUAsdSnbTAGIAiF
ZZNIBBPCv2e4IMZmT8IDNRG5TOSP3SwCcbZMwe2f6buDx0JtwFzoEZu3mqU4Sg+m
6gwzgSUJdJNUbWo7lgm5/nPMyqtYt1VWJlDw8JA/lC1U7NfA6EOo7qDOCSXRX34u
4joqaebed9tIqS3x+dE4Bh1Y99gH9zlmH9iLc/MZzJjQ8myVMUJV9460P+XHa+O0
82edy8AGZllTCymWD22qocaS+EwwKcu7Gpxj2+wRnCbsA99EUG8dy4fpkFdtMqPz
oqpkPZJVKDNCM2nFj4iwlwfN5aGcO+PTqg77s0kR5YFDQqWVfIoMeqasUiJVE9Ss
MOaTzzxp4+4hpJfbCmtOUx6xDb/Ka/URpJI4qHpGwPB/e3JyaozGCTP0SmnkRaJ8
losEXrgFDn87QB/sxWhBJcAtzA7KJjiVx88B5etdMTmkfewjGlMdPjL6jJZYbvxg
F44/w6i7hjNwnlsvx8OiBCMNuo7jQBAm6jKDPfpHd4BQbvp9Fu3bbtUqOIQn/RjX
maIm9z9aOOpJAv+OVqK56fEbBbHbciKOtlUFZZZQm04jjJdWc6Y6IryO0+Er8gBJ
TtojqUKbP4TCcc5xZ4UhBPGQnirplEa26VYHYxUOKzq0yH+9SnXlzy2Nqjbf0lI8
Lm/kV66aI9fUsSaN2fJPMA5GsUkOtT7WD+nzN/i980X7qgmqyb32FtacX7Djbcdc
Vso8rjVO6vZ/8iQP+pRioS5sZnHDXrn/hwwedWx2FHSDLfAKpn6q0JeZKwbLSQA2
3rNuenJYJBX66l/UfXOPtFZPgNr3inY1ALgmi5BBaqP+TPsVBCBUJGbYpDnKj7Kj
4nyN24RxhYtXuOK/oYJAo+aua8dyz8ivhTPk5TdQ8GobLZ5cF80a7KzuWevz5BcG
ycWD0+DLhF44S0RqBF4+kPC1K4+JYTTskk/yeSsphUN/QsashdX3SRsOjiNahugn
k/Ib9yGT/rnEMy+fvlphKaMXCjM7fZPJ8kQAbS7n2SBJAwzfNhY+2yl+O/eQsG/+
UOrkcdt+/yFrWle8O+FgNvGzC7AdKOy0YuFkFGtJ3o5mHF9zVt7dZfka8OKbY/Nn
xKNNHpnRZ5iGpv/tA/VPHISTPl6VS/RRSzP254OR3qYJW3YyMBmCO4Xy1wR8C2B+
4w468b1+p7kI7OFo91+vtbM2kqjYMhhF5NasPdUn/sx7Me39luC6IK1kNeDAUUML
yL6o94yx4W9D8eSUvYnDFmhBOHm+iT8K6vR2lHlZAp2B5gqC8z/DTMHSu3/IRAIa
7iEW8J1CGg4+nleqKMNGZVZe/gKCgJeebeKC59tQbj9Dd4JhDGMfNIn7sDt6Gs/O
ojaFY5wmOOD+E52mepfRjH3bnKGLix53HMF1UQ/3uTxyKoz3y6TLctcwfvigqA8s
9BrHEnAXfKBN5GQIYyfI1ittrhH29v5rL1T9UZxRuU3av9r/1rm6ESMns47neqhF
DclcMs5fs7xbusM54nNhMAyxq3iVsjgNry48v84vsZt8tzX97JEb1jBhu56RpgHF
+3Z7/r8KBsNMbxXnwQuX5ohUcxJUqnmdjJwnWp0nwGPkXpP/6dJh6XBW4PnRQZ5k
0avmS64TCSiWtGfvBNHYyVNa+KAqcvH23W1B+y0oEurXat+mPoqsr3isppGfQ4BF
HDwAmiFc+hv9dZO3n2juG1FLa9CuffphawAZ3lEcnUrmdUHIVmwniH8LNjo2JRl/
GGyqFCelh0hRpoqduJj9gOz9fgoT6VInhUMVnnot8uFjfYUh1davOttDEyzAwoya
Eyp5bRWdVfQ4Z/t8nLz2mveP22xKVLiAv+jUV9CyJvEhoFlmzdG4cl2Ko9Xrb1iz
USZYS8PFnyfi56OGt2WdlIl3vUfScbM0Ja56HE7Jbf3y4TCbUKf1RUiL3KdBmtKh
0+5NE1uV61v+mnIkIiD3SgRgmNsSRS+b731WcBiMBl3RJPt9lGb6UeLgIvannV3h
ljhSuMZgnPvCeqIdr5T2tqRDMlJerBZKgGIs3jvgoqzBYx97BIJsetGmj5ctJYJ2
JmlvBFTGjUfHaT6mflSGIU1WG08iyvrmNrRY90Tq6V0UGBSYFfOy6KB5xValDElW
8hYORKkKfrFSMhajhgWiwC6YrUEZvMu0k+vo4rTBA++DOv2CZRLRoaTtyCK4ai38
p2CI1c5TOnPlLLelciR/C4RZDKByfV/jwVgsLn0+RGisHeOYyVmIdxas+ZYsAORv
9Xde6tMteT2XH82VhyXEcq6rOxVjEphM1TkkK7D5FTJxXKMP3Ot+7LHrpBOBp0c7
ZEkWrP+EQVIZtFoMXZMu89zmCxAGfEQSltnS0viZ0gr8gWbFv40Dh7HKr+jiL29p
u8B1T6ZVCIm1K5RFmBN8N+Dcp6o6sxf7fm4XMF3R2vBQ3OVEA/FYLD7Er5WAoYD3
Q/ZBN5KdYpiP0RqNkIbuAtw62rWD//DJgwyd6ISpurr1tetuY71cLCS+m5Y0K6dw
qL+9D3JENXVJaKXPspFUrMeJFpFBUfhNDcyl21EE6pPGULreUKCFPGMZws8FUmX9
XaxyUppr5z6GRL7qT4Y5ow2fn42LkFKsOqF1PNwA+hw15Pp53GH2wB058IXgVSJe
dhneXkJnAInqOaScWpYpK0Hf/cGrrmh2aN6ruWie956wULDylK2LMXxuYHtZ+/b0
8xeiO/+BbYjSV3RukoJtie83Y/aBsMvijf4MFKhCt1aO5C+WAaP8oRNpxjANDWsu
wbshXKEbuaOE7yn/MshRQSaXlam0eJGD8hrrtnzmoLt5bfuooyrMwaD0sKMs9vbT
431aTG+WWT8AC1KazMwW3CN0jyKwWKdogJ1HU56inwl69z2r/as15tv+wnIwrCFi
NaUKAsmOJPn9s8GAghk+s984Ug7E38Q16dmynMDCN/0FnO4o/mjpSXgnJf/o9+V4
mLV4KHMo7eU85ZOyX9K8RwzcwXkmexSODBK1LadEq6wLSL7od5ZkpQ0T/c091rgr
XOXULfj0hXJmF+D3HV49pZ0pB6AMAV5p1i8bwSnXBHzBfW3pupNhJbkk9UG7Lswg
HGU7w8yqolJHl/ZOOSplk6CeQSnSer3aegOMwdttNS7neJhvfqUSIWMc8ETZ3RRB
lGKmaKea+McSbstRxe1sQ/XPLhOmmJj1BppJcf/GMqBAQz6HS1b621DDK90DrSF/
V5UjtcT+sMzsfb1CjvpPMlHKimgmbUlMtVJ79tDwJkBTKmDhmxVfL/nbNXKTFQBJ
ZFnj70mAE5PJJfxJ7ZUXuxK+ioFhGPJ3qtFfX+ekhs0VaRPgw/LHFNdJDSzY/5w9
icpuFkorXu1eGxFTT34jx9UoCrwq5/EYtxLf8YKEGIJOdfw2WoC1P1CyxykYW7Qe
kgz1VGtPXYlTeEzTpEQrwsET6wxirJGMJiCEqpj2KZ4hmxcrzcL6R10A+kTQccZV
sqI/yR4GrIwrjXrymCGjUK5zpSeP1QbgGRkhLRRRS5uKemnr7rp/3G/s+0wpy5QW
pYJDOvF8bf120M3nRLFx9Qtvu2E9BEocGZcmFZKNXp6uL4lprxI3z4RedIjDqpfT
TQLkh3jSUcWpSn05KnzKBMj9LCMOr8y1P9V/BZqe/AQL/UpDqtwzTaARdaRaBoKG
LE5jyFGXWnlShq88EPBs5Q+9a3+WnRRmQvWW0HzjeRuTRYEVvP3SZ+4byziOfQV0
G+cE2Rls7soUCNSv5U1OH7GbVSC4qsy6Mwsx+UMVm+BvFAowVAHbwQsvqxuJ/n4F
B90kxE+XglrBAI9SJQbOj3Z2/IfIEC6R40X6Df5D4y8ceUCYWSUQQ1Kz53/tgjZV
NeZSevHS8KWvt49dldbOQr5ZqCMmENT5sTYGL1X1MxyAdP1Y42t+qD1SLlmFERLR
zjAwd187k9I0QllhurhE8Q5zXlaPSFtfZhVaV/GvXj8Rl+G9ZsNG81Sr7XyD1yxr
xf7fwhIa3/08ASz41y8QapxmMgcTLM12Y9N5e/+/RfdKCcgo8hLZEHfC4ILI13Z9
JEnXo/oNLjd33qeq7rIC0XEpEzv4KPCcSoPa0m9m80eXevqWGlWys2W5nijXqY/N
ar9X9E4K4gyxByDsP/7QxcjA34Um0KOyx5woQMyncautx3jsIAuppfuMY6Yi3bi2
vvyZ8gdGzX2McXUWNo0wHy7Mt0780BzjH79H1ucOa0EpeC1doDyzdIXFUs3mF0+f
3F8L/A+RkfLAgAGoBW1/9J4ItYG1oCklQvPbgm+BbscEZkIw7hfGDTSAiBM+NVwn
gyMrFUCD6AzqUJLVwfX174ZKtybKSmvafxmxTLJ57+evjFFocUx9l5X/qSiJvm6B
RGXOt6G2mKmqyRvZCF8DIVfi2/PCL8IF7HAKOjVumzHC3Cudo5Hu50cQBdKJ45cv
Kx/a++88Jxu9rKMMDx6p4D0tICLseRO+rCMHbF2/M4QPotxaEuahDjVtpuv2Pxgu
wXcHeGfCRESND7xnCaOvsfJ8+4nbYoLEBNp9T+Tdb4Ob8bCo0Hik7BjddkWVhgb2
opM7FHY7YOReTXQWT0R7vBGOSU/QWq5hFlvalPsgb6GlTFP1+Px3Fx43xs3ukNWr
3DQpcViWcdgBCZ/KDfPfTY39iof0OkgBy9hHYEO42tfdAv5ZoGSwM3vEX0yzxgmF
/iWScQ3bXRjqI491eOq+vkoAjEAEud2LPZvdE0L08LNFDGmS265i7E2AMD+ydf6L
sUQtkW9rSKOjzdhHwMbN5P7jj0+EH0rUKYdDfax2amZvwzgMlEwZR4vdOcIBvcpL
+HL9iOybzcC9xgigeahtJy4kceCnyQ6Kuht467TuX2q5bjiqTB5CELe8E5860qTY
xD0fobyGo3fGZbAau3YdgW9tz33nXoEAnVvj3ASqLPCSdqlHcCvrPohfrokM+YUc
Y2s4LaQvW457VlwaH+wwCvx2lSLbkIcXwh57sk8AmTQ/SVkFX0JcZ+LVCok7tLvM
h4CPAcODkBm5LjJoIXgg/o27q2Agol8TQ4WrFNtbNEEQbZtpg5KxwEupNYlCyZq/
NkBvabqTeSWuQ5VjFlfeFnTs4MkpBbZ7PZ2XTz2RGDIqYBxxOsnW2CwRcAtjpSdt
2S2wp/KorKj9kxCKUoKbHKrNPoFtRIep7ZeV0V5S5pedkb3XqpUBSirsNdyjraF7
ohuSrz0wh6YzUu9zuGViUxbDRAyuOlkA9A1CD7iKRzF57DCLFP+PTl+bY+60dB/v
OOBgT5Xh8ininlLzefQMB3AtmlYmdshVnTbU3bxLD+lDaB7n79/JIiGZxlB/BRtU
NUj1sv1PMw7kFIsxbMw6uRce1cEc9IMckW2ywX8Tu2G/aIDJOc+LdWofPvoIQeVJ
vjqaHZZ/5Cr98fn65P7BYUtXIifzIpwzCyqMRbdeQzj4USGALyCLbAcO3OH4MPTK
rkFCku4zc18eaLicJLi4yPHGEidMuZ1Vt3BlzSgj3gqWRBFWC/RY8U2jKSvE5iE5
jBqmX1O2UosWSPJZNzvI+J2r9kVB1eov5RPSwAXS8v/uzFJowtC8mzux5zV00Gbk
u9bMU3DAkXf1niQdgf73fAyahaPtkGg3z67FcDr/Vq3RTNfkJQeVUsrGBloSmw/Q
6jCq86kGhcr/1l86VvWcdnQXC0XOutVfcc0ocvdtdLnlLeb07CpIhRsIwzHtgv1R
4OkrFOmXs6tl2z7BBoTUF49qhEZ7p0yc2wegwBysHlcwEVbDuhpyJleZFgpDKKw4
gVaQ5Up40D4aD/sZsUbczIHFHZ1P30KSZvjDo1+kCyt010ZK32wCRkmefLO9H2Tv
ZL21oCQBjsf8Xo0mXkPzImmpUuY19ZtsIBjjeulwJ19ggoNRi68XlbH0gRK1+8PE
f+9cMrW6LUFkNxsK5OG+Desc9/7x4KYgp2nwVvVmM36gc3Kec44nErJZTTR0jkgE
C4KH/jukcHN1hexU6g+ttNGCDO3sqtQM/jECv1mBppp4IQtN/4NVQNk39mpRgQx8
3+JG1GXdudpgY7pjPl7GUJrQnqJcLoxuUr3QjX3G5h8vSeyXh1T1NXTNfQZ5ys+u
6moDY0eVvI9a2uI/G+Kk7xVek7TuGVu7Tc97UrTPHcc=
`pragma protect end_protected
