// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:49 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JMLO52sdQrZuggvtUG7TpgjafaGonzXeOfToAeAl4sFajy+D/6yEVDKTNg8DK61a
pps+Kc1v1VZ7TGvq9lS3YY5770dbKBfPq+rB3IHbKP31wddxMrIiURh5Os7BKN9J
/1JJTl5jVunRATJrl4JyiUdIv4g2kW+v9T4TFVWTKLc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1760)
4Clp1DGiULL7a21FAhFQ+im0NocsclT+ve//yeOgd7QNViR10GWUBUKIY+QRZmJj
qHS6yl7FXIVzMGBu5+VFdTsAhzCXbSI7IV//EukvWkTm3uuQ60Iq+4E5L0PWJ3SU
Jb2oQVuQ1Fqu2R88LQ3XBcEdwy+ntAGZj70ztuNwx73izsT+Y7ChU1XsUBGaji4L
ebVri0lCeShJ6HkHUuBGNUy+yyTq8z4EQsUHUEIknM6FJJFWkAWGlWlS7TTF+DNE
R+FpnGrkVRN3ESgQx6v26HKQalPm7+W0Prjqy3Yl8C3Oe8WVE0DDFW+VgXe97A+K
Dl7vWqtpl9eg5N4dKPKr2/Y3Z8j5yETkvUxNh/BUYv5HNUL6+RIgH2A5RqgFR8uG
A/XXgxWg9w+um257aHTefOmo0qEoFJ/rkO1w7lIqbqt8HImDOfUL/7DxOcVMZ1l5
m+8GtHhDMtAeN0gPvri8/JbUdEJP8QmUyAR6v8X4Prn+prvKJqhYimJX/PpMMgZC
nKF6OtPCN8kUROyvDdOi8H0q3q2mef+7YYbgSA7WGPxNBdti1LD07490aovq/Bpi
L5C9Ls7VkEA4sIMaXQGFHcLIjBdWHvKkUUyInWG10yqLUjhJ7Cek4voCuElUzkST
ZBuuX8VIWSa50sQbelnDjLvsCeCfzRtBCtnOHY9P5mRM73csX6UA4WlH6Q3mePgt
lyMqRjtbOT2iRfur08kmj+OuIezaPN7QlbduqYjxLEziNBDkiwI1dT5if8D/GXlw
6mJl/i2DuEEURrbWssiEJpXxB8MEdZXRoPo7guuLNCogdTSZY55ahjF24ayEY21Z
PhhrqpD+R8aOMZ3uCAQMCmQK9FeoKACoEzLUysIO1n7M6udF6Jm0tihBjs9cFmP3
vfOOTHUNDcSvCu/jpL+7dC47JQvhnWUOz/8mfVnckQ9sA7+/hmFsWAk1BUhvJO1/
WTlwhHbjmcbpIr5x5i4ODPOQ24XfN2zwLcnlwLRw3PYVd2vLchX/sEIDiTsbhcEk
QS5pe1DIiTNNPN1fBpJZVS6keszNJQYf2fKWlAwK7p3uIr0x9q6RyRHZ7OstBd/i
KL9Kl2Hm+rRNV7FBZb5Qwa+dLgL3MvYqUDwXkiIQFue9eG/i7tpmH9zlNqJDq/pI
nvYDLbSNTp2CuRYjbTxNv7TiJVUhKlEYYcNVgfadI+EO6J7ggKUol9NbkykQMoD6
E6cgjZNnwMlP9206J+Zf75hij6HK/wRhgVfg3yQAVRUkDCjsFclGTHzqjs3mqCB3
SM1MqbXBofPbRQzR6HW5yWEABOgiW1imX4vwJ0m4GIgQnZq59NOoBhCpH1Ib3DfF
tW15bm5llTzu5RSqb0v4GN0FIvMDQggoKlSs2vpm5vxcLqhJ2zutMl9fx72C1YdS
CgG0bYC9wz0uY8XUb4sbxEF0tU4HnZkkQ9aEq0Q6w7GPW6eDY39lu6gId6C1sJfZ
bh7KFMMjx39i1kJBJV2ipH778t/mavEP8z4e3kG1QqoQv9qJggvM7UEQkK/iGCxL
OgZuWpI2lFKbn7FPuspT/wXBbL/TEQA4nbZ8u0JjU4wLolGpLFifGDTR+D1rov19
/Ef9LayPa6zvsEGy89enB8I/mqY0SWbXjOR6JZKj+bGWYwYZ3Gyab9HnTdSelvMW
sNBc/rpx3sMq3ktPVCw+89GXOLMUfZWXVeVUrxWcSJfls9x7DoyHyrD0jwVKSdVX
rtpGhm2D3kYEE+dHtA9YipEKcH76oN2+NXyDp1CLLYcd3/axXLErV7tLSxQ5Z/KM
usMp0zLlH3XwQYT2NYVbc49vzSZqQDEjtUTdIs12xRnh7K1nkQ0z0F1Ab9R6+ykO
EeCgy5oCv2EmNZHaTTX8sGx7byaVpGL9xH6eFK47Fww+pMG8M/jRyzhx7JsPyehh
G/IGGIqbsmEpEqpx2Zpucd/VtYolItIC6uMZGnfH6kDdmDiJVZKg4X8NPizJc4gW
zq9+/hyZ72j1bjV82eVJnV8sPW+v3qAu88AlszSST/Q372n+SVpbEw6RNkYOriLU
CmOz23sAIyfLjgmwktCK3IOeg/cJ+3eJdBgON/+lW+DyM4KRt18dlK6JPZvu3Az8
E6chzrv4+tZo72n7D1wKpx7Nie6T78TTvWrbn/2bC8YM7EQe0vSJI9CdPE7mLCSo
b9GtAKndSV6MP4dGUFrjnLfnDAQTzKgxQZOJbhEukOAC6p7UYABuP6JmvcWbgocM
vHfzoLoiBbYf6VMv4QMWkBGBqTCnfn/Q8KLnZsxZ6hXV60SDdB78vBqnuVxqXY7G
cIdzeHWPc8VSg42b3sSVOsWW8NX9eNRXnu6VL8yfxwI=
`pragma protect end_protected
