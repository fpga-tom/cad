// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
h7lct6tYQQEikWd2JQ6llXGIdHomDdzu2VA7WUiCdJSd68HCWVcva61OyZ67SFUj
d66dgpLeqXqDUCITc0/zCb2HYVtt+wam31cgxw1Lpwutcm5aZBb4DcmilOhWqvsx
d3TSQUqNRZn6uQdxmZFIe4Wv6t2f2Zc+lUkLqsVST80=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13312)
jnvqZrA0Wpjt7iWiZ0odoOQQOHNrZDkOgIJ6XlNzCcBua05qk6cqBPA3coqCpAaj
zODUF50R9t4sIzsLGTQCK/vbGnvEpHb/qdsTW9oCBQo+RZamwBAbjoI4L8NyLrFM
zQ3rKIJN++cTaJIub0EX0P+4iZuFcdGT7ztshpsTlZWWlE2dJEeXsBjrmZmTmIDU
nzNT6W9zcXEBC2zR9Wve0FtS3EWXJIOZcL8U23RbEKAGaCD8pJpxfEKqgfH2kEw8
K26QWaTs5W08lmO0PIlfg6SFIYD4mgD5DS6C8FaxJgbuns32UN+lajBw/iZS9Uta
bi+ijjt5jNOIrKAmkwTYHkbfD+VhmvyYHRXliCp8MoaqiJjEV9pDMbcbw77Mh14C
m6Y76MjzulcmfHWY0cpXSK+0s2jTlzk5wc9PTbcVVda3ysKcr26w39soPFVfmOXj
HPorcvH/HOU6luI4bEN4VRHYcQKD3K3shJ450PDhARRkhyZnQif3E2Gpjmstagp9
txCzHz2IslkX3Uve3Gw9MqhvSyXBUeiWih+sF/UotNWzdkxi1VjjIGbhJUWnLK3r
RbVVUrCaWYFfXa3960DlIUZVXwdLllwleWPRcfvwVAZ5gXkmxD9PQ1uYHyt9Sn3q
RJFCO/Xh86/VYTYMDbjwNUVUm5U2XxtQpDwBbFpQoR+1xXXiRAFRbz+HOiKUxxWD
d/TIkkpaHKlblWzWWL8LfMlvI9hdFll6wwPRFytCegaTROIMdnCGF0R03ZOyw8zp
pKRLzwOlK6pyYX7zMJd8n+xRE6vhlMW/tflhu4SlMdTBy3++KzFmPqqrgCfc34c5
f0qnPZna66CANHhv2m8/fYAFYytMOlRQ1L7/9cN2TNcSahZzb0Td+a7ahX0jwtqt
UfpNAbmOpvbUZYP4L/sIEoOeZ9yIAobGijoYonRHOmqKVLMYPKd9I4RYvhH8vnbb
7v61pmo5sgh3KIabEzVO27Qqq1QF7LI/fWZj5gAMXBNjFu/JQIKo4Vdcx8xFoHtL
WlS2OO0S4XdFhYc/2v7bdbYedU17ZNtEDWK6BYg7TcmfE+WfxNeWfXygY0UVo3lM
/YcANjNAIuxqG1oIC0Z5QV2nokQ0kCXfpOX0e/yQ0gf2u8BJnTZnArt9OXkDR7ww
3vVDmAzdhTMkOa5SuenvXoDIBSlRbULuVmv0WpF/VD+exBxNUjNVu9OBlwBd123/
gEOwZ/jZSsrUkpwWYThAzpw8uOJ4JcX0X70mTmw6bZl4vJwLddotasHF7KrhpWt1
mgRAM65Wqj4cUEiC/M5G3BlwXW3gdsvgF03keXBnaxm4ju4xm4fEBTZU4e4swGSv
8gahG/erazVgDpKIR9abtOMRn8hLZusATLL6udG/KHCrKI1cyAbFoH4W1j5jOBWZ
XWU90AyW3C90lJpS3+jxnKUc1a5PjjoEq29zyaIkPX1vbg2fToyVqSlx+wx1R/7q
JUe7gF6fR8clCzfcjKhwev5CwD43VHibRnd2DVRrtwhUH0b2oY9GyG43nyXHv5PH
NEzEseqSOndy8jJ8UoF9GVmODVvxPuw4QkDGpjhhjc2zyu3qWpxQ+IjYrKyYeNxZ
K33eEdpgFxFuYMMnyVZ5wll66tgCbrg86tpDst5uDWkZyf5L/cuME4cCXmOAmVfc
0N4eDdcMH+SU496lbrNjxGYyYKjGsmMkxw6t1jTV0FBojPIxr+XcIgz77093q3EW
fNdGdQUjn0lcpwpnLyl4FiYCrbCuPzC4/SRglhjhixnH62ymZkZxShFVO5pwms30
cNW4Im/LQNOg+xOKp0ELRgvlxHYS4gDSVdQ+gfoFf3vNli7UXaKX6OPxkKGMi1Fa
Sz11HoD/kuCt/i8GClLP8mhalLAHhi6nj/IPShiWrvxhDu3vgR92TDrlJpggjGrk
tuFHHXlKTMz3gfqeBzOU9vTcTGDbzFT/DBauj3i3cRcjY92paq5dPuLAqfVDfwSL
6qeZgIagEIkHKrRp9UJ13KiRMZ+hDAkaaXURz4ndbX8m7Zpv8jLFp+H1r9XmXjLa
/paG0Vzc+yN31yezMNPaJLj1hoBSMHvzDnVeSKzC4xEBeB3dL86siuhkJPHy1EsA
Koc7c1QsRpkTDAko7L1ac9pSwMYLBgLs4v2Wu1P4IulpJ/oqvfjPVziSCTHMZXPC
5a6TfLbyC7SmcOdCeH+DFyvySJLsiKohpJrznz4ohC1ktjOQHTyw/9sGjbEnAD0F
eJR1LbWurhDldER2oxI15N1cvKt8Ouw9AlWaL8+gjki7IblLkR5ec4nnh6MMM3LH
0FTAH31o5dt4vyc0Yhl0ub/brsGe0NgOslT7BMM7WSRPuPN3wHKdFIFaG4EqUBYv
fXrXQSOIItVjxReHEeS1dIWA0gMNEVl4iTuGeg7vuU0jWrDiAaJL3KPEzjqMqDtO
Fir6dKFtYVFjvJ99Te7IIX0NVhGoQIBA0EkQx6yhw0iFnUheriL9PYsSb6R6fAtV
aFWPlkuDgNz3/DiluN5zzQN5QdO9hk2MducCUx3HPOFuKgwYnxOMiBCewgNqNstT
mTvGiCEg5e6iXp2S1ni+uOmC78Tjs21mIsiOmhpaAFnyDkj+ZOxVlSxueGN1l3kh
EMFnJSqv83z+7tY04ksi0lLRLii1GbkTf2XzncGvyFDhDDfJo4RByHxqNOp8ksBE
hGc8OIkdGdGcUlTAs8whR4Zly9WAYrbZ8gPJgW60PidAgLainzMGDKZiLkHIrPgM
O6QlbsLIjpA7jcA6vbMCH4oDmZL6kV2fXsA0kvsUTY4JlTqatHETzFs7SG6ns1xC
DeaqapqBYRjibPXiS+GzelnRW38/5+ZdipHQx/M00Ri/4w92oaRE1BmhuNyegtC6
PMrqmLn0n+Df1CXEfkngbzlHDTdZKvuPBBGxM/U93AQxrq1x8EAbO1tsUXutz+1g
S0I3SJd41/Chh6neTm9TLMTYCuYmGeGKebBrylI2+nZ02oNofwCH0TgsDRRP6vxv
hst1vEUZwR4ZnblGzJj8SHB6dWGhGQiOVMvUqmkonU8damTKoDH/m/H60173aB9l
vOo3HVCgYdAx52UUnedn1ZTHBcbeSCf9QpeU/ydFv0Ws9Qw2w3tHz2cl8kmkKesL
5XJvLkZznvcsa//GHKYbofLSuOqxsC8R1+IXG5KQJG62xBamKqfTUpoCJgSrqvpv
CYReZJOHIZyAKixcM+68hfpPymvlMgEh3GjI6cyRvEzp+E5ADQ77vLD6owp6jla/
1tRVQ5cD///3zfZ3jRZYwhJegk/71O8kx745yhHSOOumM8xFv1g4psOhC5yjVH1u
m8ZufY4ezGg+cNe4k+iHxmYpYvO3nTW0wwbyenX5DAmbUQd1IhwqUu0abOlJVJ9a
lKvQIOKGRmS/MjVT4mrjrjcH8cBY45Ls0OiDt13CpHh7aQHEiwznU3K/9aSNM/wg
g7lx2J3CdVacn8k/R6OlCNCAcikdJdbHUryFfNW3t9lD+CaEILvc29p3jSZN/UG7
AtalgK46vF1GvLpSxsnXetcRz7hyyftqE3L/sWnYvWdbivySWWm85QiRUWU/8pY1
8/Avm3xvIo+G8JVmUI9G2X94ySmLvYe838QFCAUt9EGrtmHsUpog1G3/s+LMmop6
cOydwki+K5T5QNczb2bXy00x6aEnpa4XL2gsqKmHXg7KzromAXB6JI1iw+n2Samt
ABWr9Rhs3MZe7sGET3vtoJ/hs853H/tQrLPM78a8s4VRVMofF+Yl/7uzPGRsRTVO
ABj2ge3JZsDGnD7Kw/hHCzwo+9/oRlvhR83UaJHCnaaLp9XRhkfVP+pxvP7kW9aZ
hBME6lCg+YaXHl7WGhDNAd7bsfNKlmVsq3lNdFH4B1KaUoKLYrvRiTczTXMQQX6B
D2dMdBVMaDxo1Qo1ja0o7zisOcV+DBdz4/cOGjx71NYK80fkdv7xh6zuL7lHFpo3
o+09sd/MbAVgitjZxSGLN2nL/+/Nmm2QwGtGwboFu+n9gDuVhruW8h1/s68z7sxA
rDtL6b+P4OMeE2/GtLTQJnZKj56OK3aimmKGfABaFi+PlQWCLo013WjpM09NAikZ
0sYZHCwwEhdh5r0xCahcWjF69zE+nKBXoQFCmEmFfl036rvx2PAx9GqI4LdjuZbL
fEa/6HQUA2ro5MTduWNtF/Mk/QvC7egNkE8iy60TKGoemHVGdi3TuBtRucHPyzNn
8G9RoQsDy2DDXjcYdBgSa7jTAjpT+KOu5umvfraY5rIkwUp5Esdz1YGYCMAZjrUT
96bFxxjXE2isWGYrEyGDqlfOAz7GFj6AIg/NzH3FRpAyL0edS9dtTQjxGRTuiAlA
hxM2YmmeLmVbT5Aw088V0sSVZ3gJkN9viqV3i8M31eLuTs75OQp/fyHCBwZSfGUF
784dfHJ9wsm3W36VxNDKR/0ddqj1A1roQAKtha/wNqceTsfIYKM+u9eeSO/wWUbw
/+Jk7AAXIaBcz/nX9NrEO3Zkcmyl2obJWf7mfjxD3B+Jn8fj4Wz+Zl0Vy++lJ3tG
EZdCLQ++SiM+qLLoJIWmSKsdOy3u1sSKuoosIX6FTd3LTlRhvHN4J2250cEYccqR
yTuPB76NynmCHp1oPx5iSVq3FpgArjKLXrt7izVC6JypOEo9A6tiAMElOMYO8Wzm
HdLlH/EmF0HqMOxeL3t3S/ZBKer25bfnMBVbD9RT8C+OdTyGDdvLy8IXwfZGdUNi
vzFRPjbeyMzUbY+kA9RqYBzhioYk400A8xKADu8f6Xo1WTcO3DMdbhg0IhhDAUX6
dDI2Jneoamwq2G2TrkLtRqZ4q2auAqg03y2kLnrKM2aZaU4Ft3QYUahE46bTEnrI
yl6YLcul0L9tDb3pTqFX5eeOWVuOXBPLnEKCNPx2ErdVEqAjEJug2dHudTsvhNPq
PTQ0rANBi4PUEoaQE0JZd+ryACTE7rQ8LS/l9gBt+x8UsBh9UEEn6SBLRvtWU6A5
Rszeht77Op9MqAG8AiD4zHScY0nG1mLMWuRn8GpHV0CmWwQ/fXGEcDFeQl6JznJ9
a8jHGbIM1XoNpoCpVI5Jc5pVgmo0nkexkpPL+ysAL9OH8F5OR7OlbexxrSCcuZ5G
Zay67t116EnZ5RFDCV8JKDfx+VpdLZNKLRnIg49AOU9HwtK8yeTeIiLAHfsv7jpW
+/3uZ8D1FaUpDBTSj06U+Hoqes7vXLVpXiLu0yWe5JFaurr2HOXcof3kmGOjkrsu
OBpaZKTIghT7U4qZpYabyi1Gb1Q5gQCKooHv+To1sdZJ2wCAz8oufXBr+eMqyHnZ
KP0P6iSnwhp2RX7EGf9MxPJfM7LntubxxLwMUGsLVe03ti2Rnnhr2DcmP2dTp9xb
Iwx4Rcpw9zJEsUKSyr0ETuy8QRTO74wunaN5rgdMtFp95fJw2oKTSxKs+kbhYSc9
LMk4+uQ7WOKmFfLN+H2jALKo5XB4dwCxBZSs9VShXfCkgjXMSNsu0odxxQ1nW9OJ
uvaShXJo/3vIds5u58rxS4JckQlZJtdbwLcQ9D05Sr5qPm3BtfVk/JsEZod3fffB
YG2GksrXHxDAGSRayACLdkSpso2kWz95IQK6kcvYkMEJM6SIkH9MK2+g8YiBfpFp
cKz5vXHwHytPG9Gph1Tegobw1d/0H4HMamGKw0QNdXxe5/gE0tdWqvlc31fOhEdo
KXLK1IBBbmFbwj2TIz9LL0qvlMoy4K56IgTOP7HSkF27X/C9zFtzV4xzyy4XfMlb
G4pBPzIvTxhUrvx9EQ3BU33zIIw1u343QVzk4J5mvo/MJv6Y1gwqVDb6iile+JH9
hlrUdAxqI1y+yWaSOtqUJMbZ7PJrcK9vXS5Cy+3oiYrgCjsBzFGopHeJYFBKxth3
Mla+QPcTd2eO59aGGQvO7bMvcMjt74lwocemtc12fGWFXN+Nbof7snAzGdRj16/w
YaGz+0HIAn0C7N3cPsMTLVkTWOygo+Hh3pIG8t0SXcNogkCNf+bSf3koLP3FmPuK
Bd5n2Ju9VRqFrBfyQUqv47KBEn5j4mByqEV90gg1Mk3cd5Kl38pMzcse5TbfKWGM
w/9Uzd7ch+1LPr/jpmCXCKj+jPzzaqHARr397zsqKcpFPZ2FQcuUab2QxhqbppIz
SaHs/rm0wCzBtFo8wW89dobHPYuyTX7yO9y4ZmmIppGi8Xtg3mLMJ6MBjIvAMcET
JtiofL8Rv14AKtRhP6lJkMx8n+e+GGMoch6AoHhnHKnjh4UqZFdrZh+4kL2Z3tMC
ag/NTWK9mbTDgYsLhY9BpSdQp5Jm/BZaDx+Yd604epOPEmykDIyosLgFtUsUeth3
Yg3vkGfgVH7on8Y9dd5nzJxRH/PTZ9BPFSCbaWSGiXW8w3f4PYBoi61tx8VuIA8h
Wc8vvKPKyAcu1Km5SBxCrVlAIlJvBjXDRMK3S4O6wQKxHZt/H49BhT+2P+hmCswa
yM+0tV4E0JlVAJq6tx4K+xTH86jr/edomUQzesFxWSbdGhwbeIem4bup62A9vow7
fsRs2idYMMuZwtlgQiFCsN4fe8+JOIujn82AnEIj8kL+cH8M1xfnouMxx03fRNzL
x0lVYIswD7XM1HpZmYsGoqSLdokPn//CdOv7D8otk6E7FMWl8xDn3EzCyqogcZeX
apgvG5b2lLx04yJC7diHfiDBtQPi2lsZhsunoOFTtEl9T/CgjdAsgF/vkX4PnC/O
pBjMN8BxqQCq7zVuDXGtNdFBdv8eLZzmAKN/Bv5G4U3rlCcJ/TuKkMfb5t34wR2u
vYcWqwvupSr+ntUFsvPvS8hV/Zms6A/VCj6umYys6PvW7iYGUojDGaasffmeRRiX
9D/LCxiZqvMQGEVBpBAvbCo6BKTDvButZriJNfposbTsFVPgtLSXtjdRoNB+QQtJ
qzWeXITqXUIaZt4shMuDVokA3qy0obetBLvcJ//DQqMLRvN6SVeZLbFgJALF7MtM
aO1r+HCfquJmKOGCaqh0vwMN+Nah8FHKk8thz4p1V65lxOn0ADpHM45Dbj2hHK0N
xaeNf9r/HA7o33c1UdsotiJJ7kqpMgI4sv/PkFmXt59I3e3M54HOyQMDurC8hRaX
Nbykwx+w12SRTYuWdxSbnCFIuWo/0P1q4baunL1MMsrVel5WdaQ4iCOYAeN8Qjgp
vay/4q7IXtwMQxmB+cn76/we12aITr41iM+cghzSsGVOlhBv4mv1ZzbkcCjlgf3a
QC/ZXUgURHv7Lvgv/7eazby0V0HwdNN6d9mxna0pVfrr7ZNKUXEQ5Wo9DMCLx/CL
iOFm3mX8QwsX7ymBDtuzRmRMjxc5s7tOgSKI88UwBIYz98yeRjgsEtQENZBksEL/
F1pQrkJvtH8m50L0BUNky+PFmje0JJ2QUQ1u7yOASQ5jrtG1OPwaxXzhRfzeP4EA
fm4zdyc6mGy8ilfKFdKieTZbiCNayuwBD5FYFWR5FwyBxFPT2pjtrTtfrpsTy/0K
n3q5Ud2vFS+vwmPrax17onXhpaIREnpjzzU3MI+X9nCpENd5YRmRFPaGPq+yuUx9
4OqsshGs1Eu7O5w8UzyS5nLR6oVnJryjlKQORTQGJf5vwJeWNKGtgiZk0LlNHR/0
uzfitketNKNHbAlNr7LX3AAmwsXCYIpsp3XELrujXGimwB81bdxcEDn8Pk8KEBRx
5LA3cY6m4PJV47buPHWbt1m4pRtUMM123XleF005sREOZ48cLlhZ//8v4+gihhY5
AG2TZUHx2OV7IBKZcudheK2euy4T/i7jLQcQT0cMFcsy1xJoGhbEvcT+ENREdA6g
DMTUw53MCEnKE2Pyy7tE+Rqi3sF8vZaMZE3XS8fYJArj5IWHh91S83HB6V/XED/v
ORor14pqJ/+LSrjKkVM8aNPmDX6vqGKPjClWQoS9x9dF7a5cHdrCHcAobjsUtSKz
42/1qFSHJ4b6fHzt6Hs9oj1pAtRutSO/GO677ehi6yV7SqB8n/3oBjUEGcRXwdZ2
A6ZP0WIMNAJU9zhjqTEFCnd10w4+myakb7EhGWyc1LwBtY9cAXWxOy6JqBkiPXKN
9+6tiCz37TCJRTnR/17ISXAsRLDFqUA4sal62fvbvuNe3uqlz0+BDlgrm5+bbhUW
4JDfvxrYrz9+XoV/Cr93g7m6Bhe0/9l0aOIq6W4+NInb6H8O1aRDA0nXwNy+Adq0
lKpRxwRdx9IYvr92UUyu780Khw+SpFyN2UTxipZRWqy0cyExfBTn0NhR1ShTsMeY
Wxw0kdTgpgaYefHtHjAb4iSXUS69x+gDywZW4p7J0x/BVjj9N5UZi4uhxtMtCMQw
C7aQJwJpucqY1PX7Yt1Gn5+IeUnqPVBbk4OVeNFcDvUGYi962Ax7m195XxgzKgoT
Tt1n08udTlR8GmmV84R9hsDn9JdJUt5hZIcD6fX7t+t7XQFSI/wawOIotzcbGKUl
6eH8SJGO6hHx4fl7Tq5wtphLIUWmWaK2/DdA/1nekJsUdjlwpi6DSt56aNBqlILp
v/l+JtithSsRkg0BQg6HVi5+edlfZFIxtYxmMKXI/eMAeq/710jTGwPiA+Zs5BiW
JmNe/uH+PfOLEgsGvQ8clCh4rCT7JBtvQPqd8Uyc7vZh/GO9uGfwLRhanBzU3p3o
owDipERZ9REAL0Wm8w49VnGPKF7wnUCVnJm5JOEwuzJ1SICHwnPFXDFQ58P8qLek
CDG20m2simX79pSE95TEZQb5cQkAewY53AYntVn5YnM0FByW4Fm65oZr8MGtbilX
dKbsIOaAFrVlt9byIevr/jY/sHDh3Y5pRXqzYh8yBoh80oUup8BECe1ZPUPizaMi
MVUYa3kq8mnG1wbOSy7YprbLiF9i3x/HJUGeVGEk0E3/1aJWllyvBbqzYP4nPJTW
rYmNmnlsdnCcW8cfqrYWCUzY7bal4f2YXX7pwHTeZ3yx/fmqlX2hwf/+x1HIU9Hv
QmXnEpar0Jw7pRHilzUKQ17HMyXHh9S9L/CZfUz75OoA/Hijog0d3D8aq2VtSMdC
2sThqudGHJHE2PbuI5+cGV6V8d1o6NrNds7mIo9ykHjG+e3Gt/G5Dmbnm8DOmnO4
5rYm+8IaY0hOAbh3+ziXY8YpmJsNff6EA0JEp9sDfjqADVmTaYncRyMBwS11XEgd
c0hAgl8x5zVswjKjyphCVgcPKX++rRi0slWpJjlQQhT7/WMwlaJFH2JnRpqJbDrA
Fi2wUkXaqQmO8P0DSiUYPL8TG/HuPv9shKz/bDUjJX7G+eOgof330NOpWLA+S9pX
DT230w74fAvBFvpYoSTYfeB2kFIPJe0nk5qL+1zIIjyxKCf/MmZ1P6aWXmao4B47
gSppakve/pqQkxeW9TcNdm9LBHMYw8XPmDKEoIthy8vhOOgmUuwzeT8HQRYYldJB
aRSLPw4xKVqnr/wrDvSkmdylpW9bHT8sFWA+RhSYYD02oVpSXAqUZNcFEgfR4swe
FHJ6YJ4sn1Rt+T52C9tJJ2tFqmLh/J811HjqnbAo7/c/wcarg239hhJuykAFA0EC
mQccMBrUk31l7o4gWBb7pCNGSfmd926QSOWB02WmPw+nHF5FKgiwa7inVKE5tpyJ
pqJnaAAvTuEYhTGEdyvOLKbKLAkKiD7Z60cK8YmNQxCToCyD18N3YCXgY9LdqYb4
uBy9ZNpkqmWEvofRp+3sImgocjsIZLAp+5LeW9lTbi0YJ41qfQMPFJ0UwM34iatL
/UxAMRpYXGDF1nvVGlt+ILnlHFsKl2XWRcyQiuEjcVg1avKJX0ShQGRTI9kkJGVT
TTfL9N1kM3BqC5TnDlaLAGLzBRzCx1RBOZiCzgPyw2kfhB0uNepbbMm9TAO615oN
lX7CUawnJoItv0gmfU17SPSGnTLb0AEoZBHz8DOnlrRTxuWiLEk83o2deR5p2LKQ
+tpfCQfRTKnwVGqXswqLDZyszOcfktnbSt+C+yRelsUukpBT4B/SSktpvxKtCgcO
z1X1Hp2HMGvmX8PdLkKewVwbEDIupdr1IQJY5jMmmHERGQcTBs1BhrrnEz7BUIUb
YmXY/UxaozDG1ZWtJKJCRY90XeWIgNjcBhxu4RhtYZX7PTy2h5WzKidRhqicnuGc
NyC/9g9K3rZsXyjcNmkVOxlbypBYnigk+/4ZzxjlM1S8n5U/r4+saStkiO1HrJdr
WtEBQgLcMcejM/bUXohYl7uY+O/JgoAXzxOtyIJtRzqRlYet/vwnLxmfG25xtZqD
kETt7s6+pxG+7/mvchD41fBAEMAiEP5dmgFVJqFTFSgQpcCxQJKMJKmC3Pjdt0Ps
/HgYnB8YKIN8z+hj5uZXTRDc91+D1DGxkcCcuNhno2Wp5Jeqy6Cc+ldqkMyLX5K8
mtAx6iHIREyb8LGfwBmjRfP5CVP0+tXkJbL5WsTCdAjOcwaVG9AMROBdDLjwkSaz
r8PKoQLtzz/4LvyWoqJVUCgXkf85xpCEFKuz1JOLKF2X6eee5FpKeJhOwkxj/mds
Wo1eEfZqeC2Q8/l3yetRowBEzcgGIjodU88gSTSj7zG6h9DNKCZnnqTWqH33EWjq
Xc+8vUw2hmEhVpCwvlqUgdj/tIPrep+xTKigqOs9HK1kf0dJcrPPBxzJONQpYPcB
kqah/GrLaGH3zicFx4tIQKmk+NdUIhONlW7P1ZdyNwb2g6st1WhstfQ3ggErvRY6
3dQgX/ZVcHpRZBuelanEYacOdUCLRmXeo0IgSeGN9ESd/kvhydbGl1EEl6CIq0DW
gqkV8o2wAaoLu/5UtEkOxLaWtmz6ku3+k034NzhXjMDZHujZc8CnXJD3LwqF8kWa
sVho1sqYbOiaPIXvsFijV0BJEmZlLIdkYSxcbyyIE0QjIPsBGBVQNm7O6OBX9lzS
hj87UEwLP8HJW3ruCbv7hzwpPEX3+PPBCX2RSf3MrF7q3/5ZscXtbQez8godbTO/
kltBzvuaoaX4lmPIgG0tjZzJjrfEQq86+2zZK8sDJINK/7FSolwoAkyLv2uzIzw0
NwMvPsjOqhee3LmTZiS49dLEulTqGZosAM19umymlTQCKimc03PXNuwy529Lfwa6
ed2Y/ZhNhyM49Ri4WzkU3QQsgJ3StEF6EQ8N6RM8e6i3bGs0SVgpoG8Ol5QAFNcv
KisBwcRn+nNDEJN+uwsmm3LpAtE8sv6EOJt2yQNPE3owueEmkDfHPWuARlPWCSsf
aV0AhJLyEEPZ7hkyr7UeufGD8UqBrg4etnhpoWaAHcHGLvbY6SH1Dhj9TtwKlFA3
rg5scTcj/NXwm4aNfa/+utF5r6mszlGXl5fVRU3OCoaMNLMtXLgJU/HOmM9NyqUs
56TWEpW7H+oyDfF9qVm+05z3cB2bJvm9VS1/pQjf7gk+K1gvC0ajeYiz0oMbC3jz
wH9ksrHBPVLpI5bVdFNFUFzq3CQkoF/bci6h323unvUnXuHE98BGEY7XeULVLchX
RPr17IEMZ6Sk9FjCglOlsb74h5fb03gXJUAqQg9WRs8qtDu5NSjjB5q171bk+gRY
zvnVw8kxb+lvTAxe+TOWmB1vFqRXlzPrOwU60S8xWELSIlwue7pWp41HJ1ADts+s
4lwbF6LFy4X/0weg8GHCxhrI4N2mSmjBOPrI8/mMewB1EOcNpDYGvx7uoeis6J97
fi7mkMljxWu21cZx01DAcnszp69cut268YFCk0+O/PnOoe1luC57KpMOB2I8HeoA
Gpu/AGBFJDIdgHVhj0sqR2G3vyTDMBNBKReUHD6CoROQbUJXFBy1hoTtsOPAHrxK
KGPfToEI9pmjoQBYgkHQHznTeq2ECibrIrqZV+A7+Ht0t6AMhBqN/T8RzKcihppk
wjWM1dZGYT8u4q2DCmCSQ8dPEGvZlyszYH2rlE1jNBKF0ITjy4d2I0tjgEM0+omQ
CIVdKwYaNx2P+isR0ye4iWajprx4ZLphfiYH3ovR361wgoHjgINKhXRPm1y7dBL2
XT+vLTvg+ibRtOj06rxVxIZcJ4OBd/nzwyz9f1Hvpfmqa/e8E5zmV6R0AGkrQmq9
U4GIyGiWPWmQQ5U089Ev0KIZ0i48BhhwRxLCZWrZnnhgGuyShVTMFtvOTF0LYiPa
C20oPA2846Zfnmv5Vww9ENFvOiROM9y4ZiHuj9Eb366WmjBKjQx3jrPeIu+zy3Lz
irybOJOsKWUBgE/JBfQtLssAxxbfSgEgmEMt+GgIIMd+WPmrZrs4LaCwgvgjGn22
IzmfaNaxQaF5m/554hlmcEYydqUJfhfoPxHcshTsr/5hHFloT/6eiFcUWHx2zPfM
NqBEtc2SMIeiafMEXeR9Tu6/m59gUqDqEOHQswNDPRHLR/5G+ncMjLxXuTkozLe+
sW6itsQ7V4eoDBO3nF0EX2QFZCxdU/EPobrQPgczmRJ1O9w8VsPX9MHL54dXv0I5
4k5CT+x9burLCnWFAqAsxEnPhNMXfv2gZjYQ5IovzaYDAVlrUTSLuNQVECAq+tBU
D8x+FvhXpq6B16UuNujesKJ0UDYm6IAmUhD0WsuIkpWG4J/EYFsJNbIpibBQbcSu
uqUpx9+QXLtg+trIBQ1AVjJ6G43/5ZF4/X+LznCThY2A1Z5S0U497U5IGlbZ4hyN
0cmXQW9g1ApsmdKXnnLgO8YQu8AfQ3RSW/mmX0wiB4A8vJYwrFpxHglc3R858mui
FV9lEytbKJfG8V71Pb3huJSf61uQ57C1fbcjYYlOy3JAwbWBqgN+A3/+dfm4S0tk
SFdSZn8LawejPWQbDdfcBAYDzaCHe3QLA9C0Fd7lVozuTDTOD4RlExHQudDrMdfI
AHNFQvN/VO1N1JN16xNTab+BZ33VnHG/8pzXkA1VHfaVH992+stMSG050l5dS05m
FgpcrwVvKjh2ThfYgbYA5I+L8Y1nw0DUplwgL8X1ZdZWRS6L3HLX3jgqtW3RRvLs
WMNcNRsZvVagBuJmM9dsQRiQz7mp9lHGV5wiI8cKaQ1Pmg9ZwMlgDtQA+DOMcWoL
uX7QKLQg+DVqZ2k0oZoEBeRhCVkZBBs8NLPsnM85e8nqg8PusA+KsQnvPJmzmIk7
kam36P8sRIMpDc/66Q1NYysNiuuZmA3bkqsLsPfH4VcYA7aPJuhmJx6jiEIYBKgn
NZI74IQbnklVw0opz9gzQIjBchbT4dT7HLtZ+atnrdeGRAz6fZSP3KWtgjRVocbX
JANXYAm+ypcINxUcTY6C2kS+UrIvpFcU/Pu5mAZJLIUPtJOe42XE9paPrVu6B+tD
ipTb9PNa0qcg5pWprNCGjGsHPoB1LGsXVLpFkJ9QZDm97bip+r/G3E5ryHjemy3s
/T87qoQtpxrEBMq3HHxoPXjmVZaUJzykUHruCbo4JJ9zovg+ZUGFmR56N7MHDr7e
d5cLcKgncynlCTmE1xRDDkv81J2BfXcz+ljHZRyJnA2UkO/7gLwK83AE3FRohycI
621Ht49bbdH4jbukWFbZlEsiQG7jB/v8vEVNGzCXebUR6qC0aRdtnbMh0Pe8xksM
Ww3dG5YK8x4vatqiub4Viu97PKvRIGEADFRyZgFeVALl5iPCkXfu1xTgadKp/VlH
nAAvjUPjdICqhDLS08xYd/Y+PMppzSb7IFfhNl5yj87xpN4DWCAVu2k5+ftmylJP
z/Sekjnl7M03PzW3sIJHO7N0RF9qI0K3hIzD3E2/15Q4Qh5sWKxroBDtYcdw4Ucv
E+u/MD19DnVMIev1wL4xWMmOg/OLnels8QjQQMnfUleTuSPBIVdNgrheMjhRqTb+
kfJun367PgQETM36It5VFuGXbyUI5MboTjQhXr/HZgmeMMestUQaQd2SzMRLLV54
XACkiPEZsSgWKlcnAZHVwTjLpZoyyOH6LBGtCZU51YUyaIu8maqB+exStfrSjDlN
M6x1AZSBnKuk29F9xA/qpzIGzK+zesZtueTTiRT8jlMzuEdORCWApYXKrnWnUvj8
H8Z2+13/NRj8COO6mZWAX0FR8cJoOJyYs8X2Ij7PaGIXJyHPdvvA5RfgW3yLV4Lp
vyBisKPMwcnGb0Xy2rtJ3f+NRXKZkl1di5unRKXt7BlE2VJbvktAqnSvGs8Rt95p
Q89G0aYR91fGWyhSw2lRsVK6Epf3pcnNYO3gRVWAr26naRu7MlJ6hapBC/5uHuP0
4QR07n6UVcWVr0l/ihPPuVoLzeZhrLcrw3schUkz3D4k8Rf9T6sfjQvwyEMmmmtw
HGPWNHttjE51uvpwD/5gvqleXg9ZbxvJj41ncXLtSXuCaJDk8FvpKdlsdfvkNV28
mzjWKawKDnFJB8xBRiMGiPN6v6Lrk5+ffAf/AHwFm2oT/1hjHQRQB6GhUcd6KTEG
RAu4ibxC/cFJtoik144c3F8a6kHL+HP4TwTXI4XkQrysJkUv4NhWRoV079h6PH7Y
kp5F/ZJl7Zdk3alOweHuNJ1XpuerlI3hOiTDg2BMZ+Av5MsNY2g68c2tuaKZZc0c
2O2G9jPk7qeyCoupkPQoAmTtPFC0FLSQk/lci+ylMvYMHSst86ulQtUHCRx6EHoN
W30wRfGLyFBOyiFnLZuLzbpWJyxN/YnaJECYvahcgu/k415pgZNyIxfLSEVGUQHh
D8vzeKQw4jD78kgLS4K719X8ZbV2LYcvKWPk4OiAtpqSUAem3NmZfBSiHhfDEJuz
ftQcRInOY6RuefMu9zUeOeIXTKGJAryAXaLQQQBBdhGkFdHsK4YL3G00g9Vk2sZ4
Fw8yxT1MzzRGFGV6fiq3IyYv9QIqiwR5+jkeHghhu04I3bUMeELmHlwsaKR5V628
1jSCOjX/MGJqkh1P42YxL2dk51++kr57Epe5hsD9EWI1WGfCzj4ebnBCm/04uWIR
gyeVFXQ/njxeE33xu0wnXe7hxSTrOPIrZsGvMPosuTEkQshjYywjPQRhMXxfM5Di
KpIBfrPpaULcV6rzBb4qpvnu3WMRed+XmkR3HmCI3sSTT3tVPlhaxXgxgwKUMiIL
yGSW5gV92JY7QGjlPxPUUwv0Yu5JcVt5jH1dsGMASgCsCygt5mcBIp4QEGpSYzn1
ro8sAI6ybpHcPsTBhE6RpORPsMWmSbFe+haCCP4ffyR4OuMcSdi4iaPqoLjjhXmg
EkSUl2qLAOP5LNRFmJGJVWxnybWeQVOzNdnApcieZYc9LSXpgT/yQWOERwBb8UdE
G3Uzoleo4nQGuZgnuNYZFbxm+VvDc3l0mXpyL4f/9qjipJSmFIHZ8E0yOOO/EWxb
MaM6xRktdB4kzvXsRNWU1sjjwr+INEfFg7rJBsr6TlwdutVXQp+eZW+jqOvbeQ9X
aczmiX6ahGBHl2LlGr8v346T2lIXIC3eiHkt/MIISt7Hycyu1ABdj/g5/I+6i1l9
4/9X2nUBMzLn+YrgY+Q0lOBGp6ScJT0fsVV1NsXH3gYBVtnN2hZuFnUhK2VX8s6C
H3cEsCRinQP6a6xTwR5DBMuNWgSHouJEZcK2mloUUR6rTSf5tPYgeIrnSf4VnPTX
cgZQeeUWXCYQm7Cuc6A13UtjuqyS69PgTu+oUO1bmNZ2/PlDseu65Qk7/GTGZ4Vg
rDj9YVGJHi94NH468tFjc+gBa4I8XcHjOju+r8ZlOVAeK5rgTZKaQ7zPhLo1TIl2
H2pQJ1qGk1xoV45QwcRA5HXiVWOniUDOZLSsh81sKFIERlk1F+DZpf0vJ13Qr5XE
rjl/WTtD3JoBpwFmveTy4Vcj3mh3qJZS0vfFHIRCuqwDE91nohJIP/j2iOmtFav3
2f9M3JJfBxK37yGFIPmYyzliV7Ogm7WZdiyIQf7AwU2xRObq+7HkAw6wNgnehXfx
UGyFVpvB9KrN/DGRepi3hPUgBD3HonY3wICpnWToMncR692ggHKkmoV+ioR6r51k
stfM5PR0p2+XZWzDY5se1kIfECLYTROTbm8GZXe6vk1lApT0D880T3rxYUg3iaw8
vA5RFC3d0L5ZkLvXpvEovGnXCunG5ixiIDe5ETKB6buXW19+dej0hbppwpn+FJZw
5hHn70WoaBl+2d7DRDcdPd+aSb7sCf1HWjag9Vg4XFkj703I2q2pa7bQL7x/G708
4zLIAV/WPONymuuSiBefw6V9NCjEFpBtdWcfG+pNSsA9h75crkULyNMSY3BoQPqj
QqPVAUt9rwICKD28HOF8+VnsKXf1UOS/vIyCFBo2sOoR/dqewalR3QiMCfiAhf27
sO2zrdwHQ0RaQZpRrm05TAREVWdJj6abjDh88nywIY1EWLSLAYOK3o3aD2L36Bb9
3jF4dteZiAxot3lia9iYX4yrH3zN9QKAjNZjsjWt42EG7ZAbEIbIC2yhfasQ7VmQ
f2i/uu0FXVfAuLJorpkRnGkTp26XqozXQTY9TlCeNb9GM8g0d0+cUfGLzIw6uw4j
A2W6zat2O3UJ7owpmgktUQ3X/qJ8iETpFVl5PmZKSh7wjX4UfX4c37AG+6cbJcNy
vn1iSr2zMrRHAiIiZKgWImlh8LRvH5vY6I0m1KS9CBdp8dbQNaqu4UZaOlBbP/lH
zK+RfNxneBwrmPJwE4rxTKGDDyjAY/pSI9GuAcYaHKxKOgXh4GFf/BlD/PvgEGNa
9YOfAhup7vagEbommZ8oz5B7EtpmsLJQNI7ZJO6P+VUFmcbpk91u0AN3mYfeKejm
RaXbeRmMSMKXY1+KBIvZlWhnINO7Gd+pFBgoShMJgbwDerJ6o79N75RUUmLkzW6h
uobng+flGHHOOvhi2vZnFZ8vWxYqVuo2VTFGz6M1jBZ4oj9dsnwOEdQf6Cjpmyt8
YD1MvNlzlnImIQvpzcJZotLxKYtD5FawHs/PigBsqg9e3T15WnkW+gZR/suE6fQw
pDCm8uzfFbUOlb+UbYaLyi9+MTP+8ygtNXvW+fk+80cb+Mu4i+cAYEXLWsUsIPKq
H1PL5F7rRVV2HfK4GkoUNLnefGM4fBWIWpVRvNdwzZF5jiM5gX3QtWiRIGXfVWnG
8fhmsoWSKvgYyLcgAMJNbcYKRDJIvu9CNWL40FzyvDX8gNFGTQYWzVFO5M4WTU6a
YUGNwQ/zMm8EOnW3t49JQyxs/7qIgSNNKxdcSFlF14/ib/nFaTdxuW274bZkq39W
FDR4mOOrLIcMDj3KDNqP+yE+ZxcraVk+rQJksum4gXjPc9WZkqV8eKNnUcaBiz2M
U9G8n81onS+1zSaVAMBcPNFVuBmDCfkhmJiSD1R27TuLG+rcwuiuSY8JwFJ13D3o
GZherYjY7TBASHVkjYXwO6tO0Vxcu92x/sAcclyRtiDxdNtbF5bujEzUi+d7tSyh
qBwcjo+JfFQlT0PgjwlSXtLtEDBQU2PjVKDs3+kxTLD8+GipRwDJ2xhCGRs0jy++
q2DIeXDsgVkNxIcsEs3XghXNTZX6qnneQ0Cso4RZzahYyQuWXmE9A+oVfmiCs21E
7uhz3VYQM13vdJvtRdBuH1Nf4HhxoV1eMtxELtAwjx6we8KTWWwHjE+XMrJ2w7xy
L/yGCuScI2AuENkzQ14HGr1vjzX6r8Z8vIPliG3gKkwTbDOS68ZXeEXqvVRdSSW3
BnLRU5P99KS3azWbxGCG0QkRV7CF/3KCgUg2rkEnPNcSkyPYbIE8H5cCaXzAMg3c
JOBhnU42YNB1JGT/FNr8TOkIidESJ3yJS6t1dTj3ZgNdKFufousqc4mziyB/BpE9
+kLisnAn5DsfIcAubos6rkVTueZybEMg58smdW/R/ut9Wp2hhicNQM/JPHTSWUQd
BmMGvvjEgWExtlc4JzkD1g==
`pragma protect end_protected
