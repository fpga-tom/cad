// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
o7CxLANH9K+BixaQ5qybHkLMjr0DO7Uc3XstwyxPPwdSyw/rhytx9K4C0EcmgJzZ
g4Oc9l8x9FqwYxDg9Rf0r1Lc7ahGf14Zu2ixJoIZX6YSg07pENYdjo6vKJVCZJH8
Nz/APwVLY6NwQwvHa5CmcxDvOHS+gOZUVB8rn7gaiks=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57024)
NKelG/v/Y0E4txE0xW6C3MSnL5mhs7VjPCpoGiw0wymSVvdE9ALE5mhejg8N5MB/
VADjcbHJUQESOMVOdgJ7s6nGrO40fYHO9GS+8c/OcRxU/A+HnB6ZNUHI2Hfth23N
8xHN+/fxIyYfgI+QOJEuq3siMM9VO4X5fla80kJ+F8E70BS2sHIIk9xPxDVRF6kl
qt99HJcZoStqTeTvx4gtdU7zmn5d6kTLsUoA/1mDQudu7fyQdybSthjp5q2N91oI
v5pguLrV3pmYowF7z2tZAYtslg4p+hSQo7ymB1LP2ID8oBQnxOMuonFDQnjQXFb7
h1+VlPOW+BH5zepVyUy0Mv+1oAivUHowAqXHn6gUDk4bEVCJRbgCl4eqzDtjWRju
+8XeW2z2bwTl+lm1SF6Z6vDBYY724WxOYZANwQhcXIveapBJQ2KrGxke7g89IXNJ
W2+1y+vBrkbBIqn/x8psqrMVjPYGseKONbed6zQMQW2VXSmYOU8THUAoH0+cOVXC
pDQeaa/SWLSeG6eFeRfEFM4iICpKIm3ZBZwxbVY8GApvMCla2oDSc3wJqzoBRhFd
W4+RPAAKTyjR9jbJ1LIeqpPkIOm9oO6mAOdRi4wLquoc20TtC8fLYiWpcBb/1Wfm
V/UoLRt4jj8sdqQNPSnAXj1J5FxsqDdqcMBf35JbwUZKLe6E4MpGtgGatL4LNnw6
hfBTToAKKpsliF0im1OSh5Z5H0l++NDT8nJCGPKwzznLYhvAPptg9sRAb5TF8hmJ
GN7IT6p/ujIW/ZDaNvCQHEDMg9y9X6A6VmnX1WiN8JzuF15yau3ZXRahaE1lLx/r
mpHjUQ9t4E7rjUl353WoNdxboc7fj9hkOuBJq0T+UTOchNJCG5QHVqDkRTx/eVr2
SZwByo0pAuqpOgrIbJ37xLQoxsUL73nnQS5vv4KNCcX2YKk9b0rK5OJqveBOAL/o
LnhyDknhJunW8LF9d6laXy9uM1GuVaGUYlsa5PtBgDoH4SS/LWTTOsJKBablOoNX
dxXs8Rs8WthnID6gM3m7Wu4S+nlMf3OFcrWf0IoO9l744ibx/iKSXSA20OQNY8gw
jt/TOb2wfQbx9VHfiVIIVs2SQano8Tkr4izTM8egdP/A3Ftuf4hi76zD8S9ZnIk/
a6QsFS3Ljv4yx1Bfy0SqvIvyHqmGdWJxHmEt70Sh59s4hx7NOnGRn6iSmvQ5jL2t
FQN8OLgScUwBHxHFZNC2jur+4f6IqUpsrsVBjrhm8xPGTH94sSpW/qxUkVyQP8KP
dGelD0fN9nwODGd6E13lGLP7PZ0D839w8GXTv/9Ttp7/lLTVmxSsgPbJGeKyWn1U
Xr27VBLf7QPovCatbIiMeHLT6RlQNy6p+tUeZ+6let4+AD9uRKFCXMl+NUoJKtup
KN9fe9JZqKfT4pbdZ7hgvF6Sgj1MzvlYYEdXYV8jE2ou3IhOKVyPICTJXzfqlRSh
OouLNcxITSfjqPfACD7AQ2zrQJdI3QHFpoUMx2lx1nXRMXvbSdOLSbE8uP+TioUu
DAvBlbZw+e/cr7GRxRBspNLAqxOEfvRgNBz3D/uZqOBpWS+wUzBVTzWFPVhHPQV2
mIKgq1qxA+BKVUkfC2TSIbSz5upcWKkb5SANVPNE16QWKVvIplURwexVWcadLN8p
1GP1PcaA2dZAl0HoA0li1cfGeszcYTfE5ZjEjaLUc7Ub1HpJxKJWMhEW3rg/FlXX
JeG5bZWh8rU49YGp4/zNJE1+Kn0hukvyWwYP3kl+JFjuGSB6qNk/wqOlwqB0y2wa
BJto5cEr3jieWvqj4g63dwj0j2vuH6L38cAQKK90yWk7LWSBdr7ssKixMqbFQ9dY
GQMeeDk9qi1UEA5STATPZTLLpYbp0CNIo9TV903L5uiieVwd0bx+AcFjtP4nu6dv
MaAZ2mh3e3YkmAUL+L3RGvSFGONehVpAjz7zv6qf2X0MRhQfz83ROHrL8q2/hKdm
Mphow81oofK1Nz6r9KKZwOFJLECT/0jOX9XS33+aaYeGUorFku5otTYB1FOWFSdx
tuDDohY544Pr+c4DXkhKV3KJgP1E84awl0hCxPfJvgqQG2IOFEEvD8+gN6cDfI+Z
fzvSNlx11h44i4iH8nnPohnHpFegL7ulLEunmUMFEPBoe7E+GL74ckdehAF+u9HZ
zEJaUdhxwELfbCjLLDFd1xmVWA2FvBHGOo9dSswMaec/iLlEFK7Mybuqa0HSP2up
Pw6YjaT7VDQYQT3ATh5dvdgLFDru23d4X4T+FXeuBSiru9qJWBTO0DUDyzVg9mZe
82lwQMHm5MPO2/62Z8N68QzQ0/VMivimAie/clCpTFipJGU1XrkEAmLm2t1KZGlo
5SdoHpanSkVlLZ+RHQhsOuwmFkB4aSmCT8GVvR/fvIsGgxSjyO4MOfvnM2NfL3ui
VsdZiHyfsVZh2BghtwhSbTSIiJ9imedTokrfoW1jAfd5oI9RNgLXtW2e5MnjYE58
AY2BlEtP4XSEnI6vQxY/XyRG6AFGgqse1uO/uuEPASsKg9bK5ngW78fU5tul8kzR
2YvneeXW3pxp2Hl9mKGsD8ZXYbnNC5VpWYGRAA0pCDsi1dBf92aQQKlm+h0Wrgo6
cs5ahnxvr8N9x2/FvyyoYxbsOXR8KPSrFFUOw9iwvQl009UTcJ6hv65QSY2gA4iC
4uM3fiQOcoPYIGUljYKOO3taXRfIDfE+o9VLtF7qgD1b7y3o9diKuXfcXEF3dTE0
lE8WiSx7HQt+5NJLJ2uZmPTaRgUz81O9EGfSQWzrPwDlGix5fpa/En6K5sgQF6+U
gpJ2SGNIsjiBu3kvNYj8tY7xcMcAA1d35u/5M2Ayb5s21Aak7inTPsmhtzDHwc2A
zKD4puWbnuXuleLZ4oSBMSEWyfCeAR17k4g1DgQGmf8gGE6EWjKWyNBKcyQGhZWe
jjo9Rj3MXRpLaZQWKRbQZButuVM6ZElOPPLLZ/TBW1FbOWExwZ53Ewj6y4m6lgbC
lkHHiJ1vuIri5ZjuC0EClSTxw6PeCImVDLI3pwlTjhCBd60XYqMXX6jQWoZkCrD/
wFpoRU2EXp5/lRuaO6RSln13OOsmT8mO4RE5HhD9cuJQJSS7OY5b0ZyhexojuKYI
DLiudJZyIS1LOqy3X4UntHJjOyUn+KguPLWGn/jtPXTqio0C45/EIzKO6R4OuJbu
1W1w5OKLTfRzTOAcqJevo4DHhayj4KDY1hBdvFZ7eCHU4I+awiFptcugbNhowcDM
G5G30ik42V5zxY7s9a59J8ixWa5Yf5p9wBOt7bH9879Z7ZmDEVMlKtfZ9+LdtE31
JSvhUtRqPfHG5x3/VNn2z5GNAWlt7OQ3DUnEVe/jKIwsQveEDdEhFegtgskU6kNu
Gj3v86Rw4kDl+0CBCMPe54AMzNG0VuJmQ0tbKr12TcYzr6prRwOcq20vqgS5TjMs
jRiFaoSGGXIUobbLlKlMD06MW7BiGZs9qoNJfOs75xpS6gznJQYGLBUIrtQzSDCf
NGHa6BgyIet6oXgo88FU1Guiu/MovK+WDejTd+Br6qzeDyaH2au6q/qlgiZBNUbI
HJl+mvOOSkMo+QfC7x+cP4ZIsIAJJd1sp+B0d9dEQOfU6WRkLfnreRjkLQzmeLl6
luNJlq4np7rD7kQTgiOCJ/bLRnAFPCkIWxBVRtbBYCRWTrKVaeBm351Rb03EbhTG
TbpflYfCgxmnjtLUHL8MPOY/I2bNf76Ce4gU1h3KLUmlIXLBjDsdA8AvalRjmMlx
CZfqV28QsBzjAO0HYQTDGAnyb/XUJS4z0V5cov5czS+hg4iTanD6Lh8Pk/D1RQlU
3pyW3TlGr/+qWRaIEOpcTofafUiqVLacieuBtFC2+qK74VtbtNpJh6Xc3x1VSgy6
AtR9D4I24cjGIk34Dr9/SS7du1fDls5kBtcZCr9XJMdY65r/oGDTW/NDvkc/tKUs
CWdzurcIvcXXTbdzDAfjgD0xmMOxWtGavYnhiS5hztXR/WdITzpeyT1ayWIu9WOV
MuT95LOQuhKCuTZcN+BYw2fnmQI7NkFcHXkpmuZgBwtfkXH/9ah3k23ZAiiHQkNA
vFHJmgE34bI47rx5yrLLaO3bdyuaQmQHDxQAK7ajRMMKIXTmbiHzIHFnUCsiAlgE
7KyQ9xqyxW9St9odGSnD1mgP0wuwxc2PaF9902OTR551TmL37sMsSndxN6WoEhYZ
0JbfF5nIbr+RdFgWyxtEjEqX27FrbHlKxFhc0OGVNT8Diyubm5JEqYlTE2iDxszJ
QGoV6d7JTdaRt37VnVi8zTSTcCjvXMUK9SHX83uqXU0KDL0/z6GMMsEMCOnUmofS
XUd+0Lr/tnAmg1diHA3wYbsWEw7L+NSb9i3NSzHelrXNyvZTeXa5SMkaUru4cRpD
/lQ1bHXPrxd90ALDAIXr7A61Kn1+4XVLqrksz0MkX1IssRasn5uIU45lt7CJasWO
3edj0tFBRUiu6mAKQ2Y8BbTtdZfe2EvtV/Jdv8Iq8ygprICBtD94rQz6Q9GKdqry
C8kCmN6S4dBwVO9ElbAUti5YcPpQeiARqVgt6k07rjqcixPxNXjyiHU68O7qfhHi
z761i9nVAP++Eo10eVsi7V9wd+P1Ao1RVS9UkywNwFODRYE8uDwEj/qO4NdRS6St
CzcqVlA/s4hYun31XPTWQUKaC4PU7jzhxu/PAUFw9Mmsl+Picg+wv/Pp+MnNwpQ5
0EDz8cBgFzO8cEU0trFLeINtNPUxkptT0GslLpID3E6zrwDkWHfVE4e3dyzMk/tn
7AVGr2jZRFZdk1L3UZ7QqJ23+1bls7vWuoDzlRcwprg2iwXv0uxeVXFiYNwb6tEZ
e7z5ilvBPweopJjGP2DSwW8+V2J3FqaapTnawUaa0qfWxP6vYORJ/glkaax8eWFZ
wxrM3dQ+AB8wm1g7cQKRd6xH/6kXNFJKHRLJHAR9rPw1rdReGCMHci3XmHdzoPR7
xcYI15hwtrXJ08DCWHK77gNY5/93k6t8qJnFkwO/3bqTpNv8Wn9AdlFCCWObEkyV
mphMP+gapigNOsAuTi/7VFkCtmARJ7Q+MzC7Qixle/qyz3pV96iYCRLIUaCSYXz8
wcilA5j1KnV64G7KMnL9ONS5x4AR4zB4jotZId7dlgvQl1BsxOfE3l9HtnWyThnJ
l58L9fkAg1977iQPtiFgesTLkl+MCEm6l1hdLrNmlkEo9dFgkr+9CJJoUZMaJOHC
c1CF4O/XtlXlhkUNLEDCfPmTpCR9pOJOHpOJB1z5ihebVL/9nnZkHGOCWCSquzzr
dNmuP3ALhqa0fLpIczmMXlksHBgKNmmteIHwz4al6Y49cx4DBrvjPoXRxM7Et8Sq
bEEbGeFqF1C/xg7fJ55h3ACe87hCsLHfIHSIrNbe4qdQs75ANPrL5RXtbFIyWNqK
P3g/7+K2nz+Pz3uSueqTz4kmYrbH3DUGKF1mkMwJGxOAZWoveiggQDPbX2XzZ910
FLb29+tXnqobH8ImCfb+e+Q+Bcam95zaS9g7xv9X4WXA5SRaNN4h2oMyl3rAWA5D
mIxqC29PpVljfeQVNqWao8/VgdMfgHPMd2oPVkh49JHpkis788INhgoS3hq5dNYq
6MM06JQhWGMGdvBdP9ZqdmC4HEx9vvp04HqXX8XL2EIFJxkfFqqOb47QMF8EXWbb
6mNNnRp+kgXl3SGZ0tKQ34A25mjFn0T1I3eDpPlol6VeUmU5vgA3GHfVI4AUP2Ft
/So1/nf0NCZJ2mGC6raU0aIzw5GGMbVdoeHz1vLG/Y+xsvtLYY2GbQdDDIBQYGsT
qy0lMWcRyYRmjkGaRV/IvKJ3m60K3uJDezlRCvvHgJDTDP3+g8cYcYCye4bZrnsQ
8WdrZJOW/1J259+HbPePAaofbk++MBzeklpqYQoiII4NPLGY9sm86fAwqIRqEGcD
ByXao/5r6tZPbOOwBkeBsP4gkQrO3BFDuSKs0pftAd/1JecJnM/A//oJemC2Q8Ng
fDZ1vYf0Bd1phg/BZN7PQMnpMpOMTWb21PtQvT2Zjb/b1SKJa/jrxLiuRaz9N2oq
jGA04fxBWOSu94anHPmrFZIbWR28XiqjVoD+J7iLnSvR+7V0phbuOn1dGkr9qsYb
QKaAOdDr8gPS5Tjp1yeNN/q5n6kaOxB8K2bMDH+hrLzwWz78+oCcwcNQbZ05kRNs
UKPHEDnbopxjB5Mudd70Qo45MW7uUjzwEcJ4Pmd9AMC/BSL0WU8X9mzM4SK+9pHZ
dLCwINfSUw1/OBUCHdN6CCv9GjHlYz3auZgWY5ogp34su2K/WXZWF1s8++BpXVd/
EStmGUFfZ9CgV6Z/2Ocq06lUSfIvlcZZk77fKTqjiMqZzdNg7sX6/vDNpb27O0Un
rQJdn2GR7SRPmc4t2nOG7iuoYwPRaS4y7Z3IHqMD04BGVBJipNVJktdfmwO6NS4n
qgWF8xTu1RF50q99ILUVyndhwCdc5bL7sDo1km1RWXaREyN6MZHulch2DfzLxfj1
5q/CW5IziJgGniypyo2RfyPTES1RPBvl3kCim83aI08zkuHI1AmxY5tl9IsbsGJR
CF4ySlMlCexqZ9lOcOCeyvKQJZbuD/8KP+gw+d8uCBhGiavRlYOFXxkVBg3m46Rh
Pb9tTtdxCOeYrPrhwVWdBBXSygl+dmRfVMM9YeEFQV8vPpxrAeOV6M8y6onTZfdV
taiN5bNYhqwGNEBZo5Wf6+Ttx38VzfHSiYG18d5hxdxWNZiAYaYvy/JHveRK4KTt
8vGtvG5t9kUQbWDFIekCLvqEdMvD/Aj8t5p6RLwcXLpckUkKA5N9fk4RBNa6jKlv
LcRx+QUL3sgHU97UHVVhLVJVgWSvYN7rmo5DmT7KtTS2A1u47g+v9GxKelrz5dx9
u9EnE/00rTgG19OzY7M4Mc+ILLDgsHz6NaHazTRh6ftQt51ObDXNA5c5R2yVCjjO
xzTEbvMPGi3pssiv5YTfOQ9eK5lhf0goTnXGvK9QRMfmAnoXkfrI4szHRdNhK8cl
Jdsy7XDt1MMnIV0aeY2KxDXQy/9ZvEmCtRDVp/tTHgE51j8pP3dFKNmsVJJeW1E0
X75WuKprxTNULyfN1QPB4v8uXCCQCoSC3NUE+Bz6n4pnJvAnTUFp7tl1TtI8a7YO
pm8t4BRa01YQOh4YkwD4vgTyunqGViiNAVKPK48SgGDdC+u8hZSlBvMigDOOCGGp
sgyr9Xsh1pdA5YPEOwBUu6asUqeImMrUysQSCLIqBTGwwe6wKKdnS1FyC0EIpPFI
tp0A7YnnJLFilXxFxZXJD10N9KNgew7AdmgnHOrhhk1O3GbZC5Kxzgl5H46bWClR
1XSKTQkcO+hl7ccpkEDJD/WPm0VRbSN+n+5AI4bQtGeKFBRYGYOkp6CrYMdHvJap
JYD+DOGsDzyQ5sMdvJ3ljZx/K9lrk3bqJ1Mv8+BbiXwY9qNajGoWmOwMbTNJ1dMz
fQDEv1fueOEA6FIVx8tockRTMCUsnSa+CtFCPOXA65cgtt5beeU4lfBc4gURbXKK
I4awgSD2EDJGksn2xr7dOrUaFsH6KxYvLVaTcSBUCm+KurZQyArmWCRjJhzbT+Y2
3muEA8uBG2Vc3aDs9K2TyM7zOmhJqcfw0JxPOg+AmB4x6hvq4Fy6mHKfXIuru3R9
K7h2ORq538mtgUaUcJbmTd+FKRfl14Fdmv7SXv0aI0NdwsvbGaxpDBlYZqL3g5vZ
RsQLxmpuomyp/tGtUzWUcJuXtSdtY30Y+79PsvKX9HyjkLBtxYKY0eJJvgOE0h3a
6ZDeO0Vw0aQAcUIXBCok51BdqNjpO93bAQpcgrgC/02AIKKxxRcOGsbVZjeScSu9
RAuWn9TfdVx0GxIE+2wRgai+DJ5SK/kFWQYT7HerHeuCVM8iig49/6JPN3aBxIp3
ZAIwhXUGaPjhX+vTtqOSy0Frd8ivJyYwCLxk2oc0lS11uafkxX4YbyiN6IOJyjsy
aAjdJ9Q4unOB+7rkktALDIN/EKn4hCOTx56un90uqaMq/HNAR8Kq4+LTL5b9xuzD
sVKGbDroJolzgdcJzrK6IlWw0SPCu/ghzPsUhaszPY8/iFT0ez9bsrICQ/brjoAf
6UMRPmgTGxnatWcovIG5QLbTn2X/k3Qs3R8UU54cjBK5XlWGdBGhWUcPTkuOdByD
CsMDe/hCM+0PnqVI1pIZDg9FuKevYi51wkbRKiVnOO/PFoAyU1Wpmta9jU+eTGVd
tLw2+xVP9tomVMLrCymB+XqBP2cL04ecemRd0spXElh1kRNn/bJZm5/TqH+rc0c6
/7a6XQBjNDCEmPosej3dLtRlNAXWAOkYRj2Vz/ovLF2I2tBErZaXN6+3Nj4eLcgE
L7AvYfxD1dlcPno+KZIg6oDlj/s8STsYjVaOXVCXQi8XfM8uhyF4e7A/ypQ+663u
O5c6Iv3pIDg3apE6LkZuCfJXYZ+nQ5U/GSSq00wLOzWLIuvlAINJGNEF0WH+wYoH
cekATvs4JPR2RmqObf17aG76SUU0uDHL8UNRlCrRL3/eK03+q6lHvd8pc0fUKxNO
fezITOPCTC3JKKxVaJorDgjJUpsMYeATvbP2W/sCrYautrgC79lBX9Qh/ewUPtL1
S+NMbkbPIeEGkS7GHBbEF5S9h9zW4UVM87Gec1kexEu8ak0I0LsF1bwPTj1Bg5H5
wr+FAcrRAD8Vxc374iQKxSwrRP/6nvgpL0oi0OHMafIb6RtQNzweojLOnc1UYh8L
pqP4o1njTxkhYHWkcxv1mkli2IsvRsO27CQybaExqYIxhnEG+76f718CXNTnoQ4d
DsxvW56TSHwITZ/wyKjS9gb4gDZNOu2415XGQshF2Ktt9cH2jP4ucrFdyz3rReC/
sdPU9w0K0kAP0/OvPL4UxnNoATTKfVE4V5BNnm7fgtRMhCqx0JgiIBAep+N7Bb2V
pW0YMI11gb8DGDdXhkMhSdn29I8eiPatz9HRvVMfog4aCTk8JS6iso2iIiyCiRkR
r0J+nqtRQyCaVmEB2fAc1NXoioz84V2lW3ZMUxIPJonRosccNnVW3ekBhrMx2V7m
G8g76zfgBztiso0wY7+bAf0ZBM6z2SzQrwglYKOdWf9uEl3XBLvaBbszG1ccOVBz
uNMJNyICimOrAEpGGfVuO4XgZTjtwn8Uqu3FmTRB/CbyBsTCw0+Ene009SRcEZRd
Nw8rnsjUsvKSOMmR1WT7GxQthM5rC3CERly1vPnZ8HroES+KmfC6/qQ4qPA0RfDt
FPoZYZEAbs6xVQKGU3y1Aaq3YsTjIcAhxwQhYVNweljtsUY4eMg+HuqJ3SpwtSMp
PhoK4EJRGNpIvsfBzdNd3RjLerWSfIWEtXVy7zOHE2wnMDgsrGb44r8n/F/KLU3y
5qFv1zwE3AA8kKpMAuDEAiyLOsjUnLn8VvvyKXa9kgUzzanuPfqrVDKfdwqhtjet
h0beSUBjwnJ0j4S27tNRV0QO1wwqvNZ8SejXOMDMjVLCoOAmg6iipmJ145pa7/nC
sFz5GIQemfVeqWG1is1WILIAl5TBi3v8M8i7b+KqfFuuIpzXoMlkrgxJrhiWRdAf
27y8TSlaz6e/Yiu3inbSmX2S4XyReYZGb65VrNiDC0iH+OCPlV+8klVdyqsb5rfN
iGJE4/WmCToVJxiCTQTIs4PKtjLHJajN4tuSP1DMNBLksXaIUv70yKcfhz3L9iH+
UCrrTT13NMnmpzUf+BSvOjZ+dhajR/IVBQDSf/rz3aGRWStlfa8ZFWmycbTDZHJL
3mrc5oB97wMcl+pPAtK0ltUItvMFJbXPNppe9PnICP3S/s81Cik4X5/lD+yDlAVy
qwxlmrCBYz/hRsicYVA62Nre3mcA3EbVfzDopP/X+E73bqYJqLvw38yo7qZPU6UV
EvS1/QbB0CbDUnsPn0PxkbUn6pEQ0rNwtijxxlAiQmKIHtQPxROx4G4kWBrD55AS
xvB7okI1pmsnhzAFde77u8eDumubadzw5zXBcQsdREQWbsjWX72jq5gk/s4WuWCy
lpr2mmGJvuRPg/kdSrvWAka5i8Zm4AMRIuaWMLSIdZX/6AVteDD2eQBgNxbU5DYC
c1cXaCU9L0mO5hiahAlfKgTYgzb/tftdYj+e3UK6dQOz+ZPifMYqi0hoJkNtr5kr
2SYoCgv421GgTbTkARZfwuSCs3f+DjHrKNTxS9G8oyfCpMKaO3+bgtkZDAYFh8bT
RE/raPZ/j3KS7i5x6U4TfxSR6aL0jxu54BFFtlAveduo45p62eSitdYTXDTrdVQf
WaD04EJJN9cRrua2ne9ukSM5Pi7grEtpQSaw2VSwhQhYECt01s8RWw39cjFClVy1
b2xW9MaLNU+gEKM739IvY18kqqkobKpSlNK1Xyb8p+Mur873VkKqharUmGys0P0M
ZBepvgt7dFWx8uu3ldbaaIOSUa4E6agGNi2YjPUuTdd1FukTYQZF0o2hr3nkUh7D
yczNnJNGireEdic98gSCKVmVd5HMfd8lyC8v3MClnxsGHjhpVJe0Fr/+hy5ThkBO
1RiHJkmfI4mRTzbingFlpKppQuexcZTagwD/fq/suT7dNmHaDUPCd9S1pZeNUNF+
EUG2qcF03W2I6T+GFYyBa5bvRgjEDrbjvyLv7xszDaODN6O4pahkrNcntiJYVgVV
yi+qH3zkedJpGtrPAU4Q8P0XtVI5aFPj9HTM87pFfsnQZKrZyzbLS7lZmIDqhnKw
af/d6FsQR7O3j6BM1umkXtd/hE26x4J26+LPaWcRESgnCVp3zF0zpSrNr+VAAGvK
CsEhVJOZO4bFTYnSZF5zeKDZljnQyedtmLN8XDShOhv32SN0v6T00MohogrERgnQ
bhnWhcCEaufcUHd5uFybyXiMu73ahtvRob6uxvJC4VQLStgOvmvgfXh6ZUIWzLGZ
+sZApL9Cb+0CvGLkkcHPZV/cYc5v2xrem/8bF/GVmzZ3EC/RgjeSpgKv2qvFPnCr
sGmLcTjB8Jt1Dkql04IoTD07xclCtCGQsKZQVcAbj1iU1CuL4jltO6bkbUEt/A+8
R1CHNxZ4FdJGD0QGyGFxQ5Zr2ReUNQ4qTypxpnpbL0wv7n5vIURm4oGoGjo0mMeH
8x0AcRC4ByA4yW2ewl3/sKeuG+LkclH1r8pjK3op7Tho8ut9oOQPEkIMAsY/eROS
ptOne+IR+keIfXkYr2wettPuDCU94JtygTPKRl6h038cBvhtZF9rDmQ6ztc4o2Pm
gcOOos4nBjuPUohPh+yh958bcBb+R+qgdvAb6CCTUJc+7hd0U0InMbEUD4SqJcee
RTcI1B3z3xHcF7hQFl63nsONNHl66lfSZNGAzMrSKVLE4L2sJ0Vt0k5pb2NoQv2i
YBBzNT67YFYoS8jq/oyKtBToRi6QoNueGAAWw0pvkxtJGYdAmDuucgKbCqAly1k8
FnA6HSzUjROOVyEDaaqr2W0n30dd8MRpAKc96rtx6GFaVVPUd6K8Q6g2V4eAuP3B
sI8LzG8aF6moW8dGiXDvEPEFaPKyKiuVzly92VSVUXZ6Yydyg7wRCViwCRKeg2wg
ZN38xq05C90W0BBf3yAc730Jr70twlH3GSPRVI4y0bV0rsJZ5AFgCRhQ8PXRWGaX
hrgYO5W08JtkkUO1/Zdw66vbEDzV/2NqQSnsqOk/H+Nntm8Kzcv3FmFdaVBmPDj4
llPfuYZGqST5Lei1qT1ygIMihMqoA7wdOQuLnoIYSlwo8QJ27sZQaLj8muOraDEn
cEab7wMMLWKvOKWD+VJ3Gd8V2owkJ6onmdkVQFpjBKK6aZeAj/HcwyBlWxp+0jcy
w5O5xjsmCCAQfvASMDVgTi5p6WPVP+R0d97YxbbFoq1qZq1zHFVX2RJUrrAbQIKh
rzLqyg60Tvn9y7VRoeTOtCxqGBX8ogqybCmCR906AWkFf/Seu6NIjGMAEk4H3DM9
7LLZ7S9LRzVAb4D3jbbVz7s+NLhdBrJ3eBepXI6es3g+TjQeEakzip/G72cOtoX/
dmKFCdsLVWkjFWcVvS7ncdEocqfVfQwVp7ib+J8PkmmdDxJS6Z5Orp0M4YUuGpYh
60+NJXF/rI3dm1fN8L/Pg9vUZ4Vmyw3L0UfD95QMinOrENSHw+D2Iw053DcpLivi
Jzs0rzm6ny5SuJY2vDz1+1T9ma1KznGBGQDqFytNvhi1GqQzbIaVxn/+rTLNUPLZ
ryJGxXNkwgwUEWQOlniYn51mkmnkI+6KYdTmBe+1IIfWU3hxVPyGrgEEsJP0O7S1
bNaGnbp1QmBBeAfY7/rWZD8UO42JS0GaOd4v9nIVHOhyv2YZyxJ/wusjsaE5UTk8
I9frATiAjlKnHwHe74WsCWIbo4CSo3k35lt4BZx4b97ZXhVarDMAmXUEhPwFQaJH
8WqCOQJx0MZGFIWeyX24RR5mZtPYLGhGgnIeiZcLoAqpHKkivn/XlEFPuVNz+i4F
UmQ9yJpySGkXCU7UHcwHJr25uLDBMEavnl6TqN31VFg1UHQSDa37KVPJb0uarc8R
8Y0Z5hY9fnJR7fImirMg77Y2fd5Mp88aGzTdvs93K6frf7Ya1bNPLtRjL9Oe/ix/
sliOeuSpnhOKe+v+4loj2XWQDIz5gmX3BpmzuRvTt37I7e0bidQhq1bGIkJUbYX0
MJqTkw8zM+Ixklx7utBXu7Aw+gatMCPmP+3mb7cAQZB7NIk38lqZtmzGNgwbAAUX
yaesKdYWnMWORFSzHrOmow3/f/4yH4b8PO+o89+61joq06wuInApV/0Eryw7uuNP
/qTcXO+4iaQ6EoRax0lNC4ssw+WHUJWef/vLtPM/u7FIv6o/8X1H4BBSEj7p+u9n
SWeIh3SDhbkAyWmmfghC+CUJ/B+SpmpJPo62M6eOg4U8Q3rskJNk5i9dHUF+QIFq
C8REOxzulmP4OKCFQvUmz50MnQR9zqc5qglSl9aYoxFYGmqX7nIcNhdmGq8Wonwh
0Uz8pFA4QYkImkwnU2sXZs3OzoxbNwpvkAXURUGdr6/QAASlqvMIyE4pFyx/rW0p
EGZ9Wm3VHQ1RPHR0M1xi9NzHLHQUCOGO4BHRLakxLQfQ+Xk+Giq4r26VJ/EMXVvm
jBDIr6drYb966burRMlVhdofA1G6f/wrK0eJrJloAzh8Lpuh4KQCtSzsu+EKyW1f
2HtQIiy7p6e2+I6HOavpEWIhGUVg0TISoyf5Lp3/hzLiuvWbT4KqYiVI3ni35R2y
Dyp/hb8411N/HMZbzm/oNIEzywMzd2siAEo9ELip2aMvB6yhJ4cL8ZEVZg+03DVe
SKDP5D3k81mzH4CcVgt06K8n1z8Lnblnuvbq5vrbsOeFlXKy85Q5OopgY9DCwjw3
BrP7b7OKakqJjYrCfMXI5lzTikRLyCGzehYw07fzSubBkOJYrRGTKMRqdozFA0FK
xIaYHSRkGA8YYy9oEL5T0KPDgaKH31gZBshP1N1r9MeJ7Dc6PRNinmsDaFmuURm9
kMb3Km9b+7t3c75CJ0v4U/b9KUie7NjwBLaCrsSvNgAVrMRwAGf8rnxaGUuNX/fr
JbIraFHwU+CSfhZYUu8YRe1T9AaRk0LEylaqD5dq+6hGM6XqEKeKwCOY/WF6wqBH
f5vzq6F/PoAgdqsx++h8p77L2arxKuUMXFFZAUotsCgEtF40DHBnFhDa2m17V9ZR
8sULMKYEVGT9DMSiA6y8eIDa/86UZ6Ql8hOhYjTx5i3tnRodmSCLZ7pKphIt+dZq
PGmucSx0B6Fpo1lWKux6JiodHeHPiRMWm7/EfXmE87YZ5W+gGAHn2hVIwVZOZJHs
VJeJ0Vj2nAvsMQSN8ZsEesF2H1KWvriEo7jX/TmMh89F0nMDIvtiUOAryvI+VtWy
3rsOAePLbOSB7Z/2ieSJwWOFAFFppm3mgD3u+Js76PIeKa91vRaXCYpkf80QzSFN
YA40OoslIZshRzFGOYmbsg0jUeMXQ+pEkYnRsdmzljzbIBj4aC9g1d60aSEn/z6r
MAP+xP16oDw0OD7t9YCrrdKr66MSSHHNbszGGG5MeBCPEg/MT1c2Te10j/+WG+pA
8DfN8bNmMO0cyBHpx6cTqq4pGio6ZHQ4Il1lS32ffI3DxHIrowmTl9QsaXktPotg
rFlJ97eoqoYNnp5qMn31k9uNNNhiNyM8LV+3OzPewCaLSgrOvcHPw0s4xHBgyLIe
P1UJJPCa9osXfAYRYh0nDTcyq8X4EJoT7cRm7Y7Dqzrdlq10lLue7taAYnLqbuc4
1oG/FzazT/hgH9glCHaqAG1JaU5kKWEYb02Cwe6Iyf21P01j+Ev6lCFLpyXGdZF1
hIdIIGvWyvP7haF2v7yego/kGAUhIRN5zmdH+qVwmq9ozuPK0Lpz3gy4QaYiLNNc
fkY9VC0E4dzDLDXSkV8KuyrancqLny0oCJbJoAkXpcxUW6oTuPGRA8lTelCZl3oh
FkZHbBSdhkPFFeRjGqk1wkJnTKfu820E1xnKRQUlRMh44sgj5am/ukQnBcGlgF64
FLWgs/4zIzCP/IcBD2pIg837SsqerxXKaF1c61tODjBuCZkD3ERuTcXh4Gv+7IMP
q2dSak9Zk4RXQjqvBU5B47Rt6PZyLZIoA5A4FoVLbxpufKffmYMjN13NB9XpqF4j
kJsjgusZjmfDHhxuZI4PJG6coqxcyG1Q2jbFEYq32cq6p7CPTwMCPgS1u7ll1v4e
nzn4yoBlZU0zWdIcOdRuTICt8NnNd9YInhDz397Ct6eZnpIxo/R4vUwoFH6k8ade
m18AKwQ2+jejEYVY7PjBLk4TxCVBxMIt2vsEmFWKIL+PvvB3vp3JV8XA29cFqzKY
cJp6wIf9d4ZoDtO106tpCR3wAdmqeFFvgdk4IRsiKpJyfQTb/wrWD0jsL3k3ulTc
dCaD6ZlOKNLmqmPr3yn5kDXGPhnbU/3TTgReWeIEoDY4k7ZWXbF2gJ1a47Ql2M4k
XwC1NPFmKs1p/AzhND0TCzSpSJz0JbuWCX/o1hewufNULUJiS+7BBVM0MycF7ZP+
GPRMG9nLGFWKUYJLvTH1tByGbtWpX9McSt5imrQxN2NZXaik5pEaLxRhldPZ8cs2
/pOb0QyDL0LSscO5N9fQFYUGL3lxQiOpq6Siddg+hyn/lgANYSVFWrNhdyvcFSKx
f0iwCGGUjxC5CRDJQHf0V9FbEaZUa8MaGvi0BzQyG3s2b2k9bSBCKgkueqelQskJ
e/pW24+eF4olqBol83qi7f4IPQ3G9UTP8uD1bmllSoqM2UdBMj1rXV4kvsbYMuHE
m+WuV6Y8yrvp2JY0WnHk62fB0za32pfWKhasv04hshxe4iIXfRc04GKvmNwrh2V3
xXERgzj4/+1rKzP6iOH8EadIkzRnK0K0wdzgZzsOM0iZor9dH9CoUPnI2V3/36Sm
HaHp5yC/qf3KnLvNW9tB44nMOYoY2uKyl5sb1u3Pm6u395dcraX1GYk0GFAO+wOs
u14lgRIqmoZcLxR8RwHf35UxdQSXvnAVV73RYx9NSJLOVGdd+w0CBVd8dn21Fdky
CAw2h0JD8EpKR3oOs+XtloIb3RV25QlddAnqd8Cza4lljzx/k/opT5/Kqcv8CM8V
2KfBjrvNzkx7FcnZoA2NjQYkMpThWiW/BY6hE6r0Ab/9JlPZBGXfuS45O+RCPqhO
y89ib8z8LfEhSvogh9JonObeQ09ZOWp+Z8pHiVDzCMJ94oIAXnVimIy9H/v74seB
m1uTIrXqh6+kb0J9uiwIV5NaNEVf1sMvwjd8VrGWUy2EuCBIjwCZoMEC5fCtmWfr
04aKDtSXHCwtQzZFti1apv5yDV4kdbHIYKMbmI1OUPiWHNv/RjLkoaotSWb0PTwq
X4np+x6iZuC0oPYNy4hno7cbt7TRV74CWYrkZu76EhHnxa0l+mTNXayCUItUhF9l
SoZp1Y7bGohcPV5yJfAt+LLOm1QEG6PH8zFexu0/GPy18vADQWTMV5fcKSX7kgWK
0K+FklFB1zVYhnU4OCRS9ZjWaA1pV7iflSuKUXAeFwKXHrJoWwl6Ygk+LdXRd935
rTS2oz8GH7TrDK5Y0e5sVrLGSqR6HwAwO/QQfv8Ea4C4eULrcjxuWlJWRFUscdbs
JRR+wkLj8RNaGQT8cZFjU9w7ndtQ2ENoZNfRfUK+M9aEX5ZTWiut/KrGDFiTxD+u
6eCtMzhgztu1Uh9bz2+HIRe42he4O3wp9v+e8y5xl3VFcz9+GoW7N99fdeVKF8MK
IIF5GFE73biCc+Cm4MhLWN/5ykk9hD3avyiSIQAdsdlqOtzQyZcp39zBQoWHPpOP
MpInegWlYKOvOK2m5WVVNcRP/ZYhhcZ2MmnWHtzH/Lk+Njft4vvMO9Tx4OmGYGUt
rpj9C71nfKlM4lvF0Ob8vB/fKPHcWv8b8i3YRHwwEM0WhlBANb4xRTA4UzBV2yBY
JZT9alu1SCh8qhy/Zo9KHMm7RVIyEmR8INvFySJ+yzZ/81JeoKCErlMSx5rwEZMH
N2K8Daq3of1drDXJP3svRBMzRQ6AyI2lR5VrMyoNHkbTE54ryheWZabeOsKMgO6h
tsUfz5W1PQod+A+TQa5/OFzDiIA8WF3/3bhVOulx4EIs0AvV2uIg12aYBQVRQcyx
uc9oYkg9xdTlY1TbnVQdHGoLBj3nxIvZCnd34uEjHZ5P5qItcsw6kAVqiqJVUzGA
lmJYLk/kkEcICVGygZ9RoMJ0VjHUWIJzxM+PJ1V+QgTeJXpBRSGo6Sbas/38iPMn
ymgrZpaT4L+AYIcyIc2hBFAWOtAaa5Kc/sU/XjvsxflsaX3pGFK0JSrpbSOBrkoI
OwS4+uY8l16eOcmRbgVeTuI6+uUKuh7ACZJRGVPWextqsaYxlQLOUkQznqixHwYC
7DmSCyXl7sP+rXd4zfJdoXp1GcBdyQopVuRRMenUHf7H/dEtSm8eA9t36Xbx3jsF
bBntEPSj6Oi4HSVUphOBRznOtN92NKkeVIJXkiyU9X0UX60bCwRv9KtEEBOe0wU/
lx5mILuCflil61AofPeOAz9v5pQwLSr874rUE69IzJoyj+2UUu+rz7p7TWK/rsD/
W0RLoPnI8I6vx+HRcEpraBuEWtBhEKjeMzddkNSxHLOBSkoJicqEniStmuKmyrQt
qXIpzsXlljJnX92yCcEfaRZ83tGQAWNQz7Fr/ML6NUs+GHawtAQejH3wCTQaSwkp
9LM9jgt2O22YxXfqJlMVwUEQyyQTczIEY9fRLrki0EXgeYdFTzOgj1+FpBtstxrX
hbOwaEWRElViS9KbxV1aMJNkVRA0wzRH61bmeOfOeou/cO9rjrqQ9dhBfc1x24us
L/eVFikRt/LrWiGAIwfOwzEVKgwvRtWkUMPDJcHYMkQiUFVuOKGGk6I37v5hL1h+
fjmkH2CMaYAeNT2/lysciheS+d9yUQGSKyi7iNVNqobg3tES5wUDP8AmC9KyY9ZY
dSChsfvDreqglxdSKMYs9W+udHPSOQ/TPQaLPE98jImAjYFVnNtlsoaIZHTpJzWo
SRS5LQMF8CRyJAd4u0lXfzLTaI1OgWwzTydYD0UvpgOZc8uyuR0jESC+5+7wkSdU
SZHh045Ayp2MudG9V+8wq0wi+2NlvhNGiwZOxJpUTlStbhKUT8VG1viyaRfU6AOQ
YS9KF+bwybdeP6e8ieRv1mVNf9Yu3J0mgiSAFcNX+tEAdfr2FwRPVz/7OWHUdZSX
oVRW0KklZunFCtEPRbaSx7Aj17cXNaZQOuxLwMJZ1fHnI2rFTY6Kf8l3+dCZzJVL
4N3obFCtKBd7QBQGP+h9vEvqAQw3nyBga0Ih0D1oFmFSA1Hhb/gqUoM6LShrIrNW
6QvVFrYWzkT17W3MrPu2Co2PUNObQQ7/+9cEpgeLiXpbe2ElNCFhllZrN2UW1BmC
N5nlDXt4PboZ66VA9dnoNxT7TbiWQVIaoOlTEOKA2zgywzb7vDcy2VADTTrujTFT
SzCLgEKR4ARvDn2gk8xxijuhfBnoUWdeIQI+cW6XM/7TzvOEnA5dfUgggsTcg+Sq
STmB9jfc8E+CPIQvOSXfHmtOX2n8uLn2R3HlnN+pk937Dnihb/U1VMQIPByUeHmO
mnIjSzvUloy2XPTW1K4hOPRu9LbfLfnNHP+ypfW2K764sXYKxtE1aDAzyCHomqU8
K97gt9woA0Fh1ESwmTJNYJOU+swaabeoVBxpniC/l5Ftk92iatCz79Kqwg1X7HP4
/6Xts3YziCZz3TkAHPRKgLg4Q7V1eYYTF0tv9m8+YtoJzTpTjRm+Y5NKojpmPWdj
MtbAL8yRKUnwEwPvIhVv6p1Ha6+QSQNgRz3BzRb15vhOSUrhZxBF2kEWiTHtooDv
tUFOU/GyITzXdHrB13peiHMIM5f8ci7/RhIsMY2QOTi7o8qblN3eJko0AFYv6KdK
UyvJDHEX7g+bYjUyWRWcxOnz6SHvhdLUI8oadFupJD+RbDshoGDYf0rmHhndRdVS
pMaNsgDOUlu5CTTzkfp0nToAn3dTKEHX2hk10Qw0r7kmNKeFq7EkyWxoM17STOVq
ogtk6/pMsSM0UD1xBegPEZKwj9ldIYiNScFcJbf42O3XGQc1MBtUW3V4usNzp530
ERg/Yjy38ir4MaUUGpG9V6nl8kwGvZTL02KbZLqHlNw7vN6r8iiSfA4e1rAuP1FR
8qz/nZ3K0o2P1LnhqqrDbjRB7eoqj+8sMAw6CHMyaDQi4memhZwaqZ4truh7BWBV
88eyxa3avQ812RcOh4lH3kiL1batR6jFp6IYLxTsEiyvC7/mOZAc/Hdvj9nA5NiI
ffjUUl9EaCaw4Qpd3X4TkabZD9Bu0ePP4TojG2X7a5r9H/fs1bNa8sko56CRKSJW
J3Pq5Q3i8XyXlUtkDOrAxdGmejRyJEeky/hVguTuZx7jYXXrvsjTgUPVRLi7BNaQ
EpIJED/6NEkbi/BPYiBEZV++0934xv8SAPyXcVaepYeGl7Lw3QgYFK6VYOgPWUvF
kxPFNcdQ1WIao05HJnemNhNkBvTxp4eoSh8MISP1Xs//SiR1n3FXPAGUGMU7vqPh
jjrIccK+kbHvkmHMOzS+h2E7fujL8gX5x4T7FpCjlVpNMFJo2qafNj5jPuv+FV+2
RO926g+jCZaz8+vLVvQIjGY4SrtYW+XYECnMY2chlrBf+JDxQCOm7On8IapxO4qM
U9jnlFeGF8H1ziawGcsW9htE/1haAZn0cmLLXbAT5Y9fx6kUKxYjTYbSCiWVdvzb
4FCrC/p9cqDuJVooSwQS7ldhFDL3DJOp29NLSECBp5cBHKu3K5Uil5Cx9dT5JdR/
osRw+rXPPm+G8EWaaWoL/lHtpatVP38uWtRryMbCfJBY/W1hu3vkmPvdQP7/6xgO
QMg75JExjp3eVQdtDEq0atCprrVn3mBYC+U9Ki/5G1VY2JKOeKoKdD/MnZrFzL+U
0JoZ1Isect6qJyrsgPeTSUGaH42IMsebLrvTmoiTLCOIyYPoR52uve92KzK/RM0X
z0mIVymwq1RGsbtubgHmHEOExBcG00z+rqdHMkReEWUngdTLKiMLESwdr87/tRww
E/BgGF9FEDuxz1+jYxYyMbynor2HfnyQUdhrSOPppYv4vU/6K+KN6yKxXBpNmf67
JYaus3Vbxo8Hoi08hHtmPHrdJYi2Amvp3pAebSYJK/3mhG0l0muv+aZpKz1oG3CG
A6Mv3CyrvGGiX3nxUV+EdhSH/tHFISI+lOqwe2cpmCHDh++lvS7dMDYWkhn/oKew
PdAYaUYmWa2gC/ctNj4ISNGSdoWKey6HRyccwOU0wrkm97Av6jowc6H2zN10gk45
N06ooG9Ps5VyXJMgfvXmMRgs1UhS25t/rip60rYIscRTORfHt7apzx5QhUy77g5d
Zhc7ilMJbSACCTv2mKCLFgB2yp/4wBmcQpfeccjRisWFM3nAb7oLqo/ipbHIii8s
L3vjxc+HrnYh9q/rJlgUP3prRS99BOXAc04GNm7P2AVtx+Ifk8nTHHXsDMe7YchH
jNpxf3SAo+qTvfIMd3ott13TzLD9+QdO9bUoIWaUTant6u+JiG4VAMFHYq8HG0eS
i1sMlM57/c3pRnzpoE3kNyZ2EjRoilmBAQ8K5JMUSOJ2mZeX7lJtHiUNnAAlOlVP
hv7+vZK+mLDFPtdhMLBrecI9etlVDaaen6w6ISlsqukEJz7UG07xj7bqvoTkJr3O
kHHRbfzENRQ9lXgpQmyTvKabOh7f46wgfIldbTnjuTMYGDAjxNSIqx5GhIS9cJk4
9TIi23m/s57QD0YeV/BOuYzfWD7zaYwYkTK2O56NwC3mRBjy/BC452Cx7iikbin9
BYPCAvco9DVZZ+z+kvQkI6g/4yjfBXOknDruETThENuVuN+3ypyAtOBsoL/j0HZI
BNqOy7KZj4An4W4QtYRRGdiXBqHGQuOFyNdvHbaeCwTOBV4Nv7xerdW5LXjGAJBM
siRM6BY1bc/Y68CDV41x0uNjRpmBQW3ihq4nuz3YaCBBNGojO9IchSQP0I/i584Z
hFuql9otar5+/DvDT39iVJWztv/Txj8NuymMW6tTasslOMUv5HcT6rYpDAqVapr2
OtJeuOw1BavnHh53LjKkmMHMmbpjUeyX+WTD+TKJDBIduRU78lOOhsthPriOUeEM
eh/lUKKyjiS2MQMl5bPbXLm6W4vSEKxSVRtCjPdNcy7mTh1xoaePyDf6jXUJVwFL
J8D7hO7Piet+aCaU0YRwfW4yF+7U9gGFmmevdUV7D3C1+rvK2XWv+lwVqWvmi/dQ
Pfpc7+ZbiBXcW97Ia+aA4F0BUW+Dr2w/mAXH8diTVURpFmYM7T5GQufPQcQrGQ4O
Cax81WF0xCOA1gq/3QZFBn8KkKHQt5yZeJaGe6eZj7gyngGWirq5iM6gXYTXWkCZ
XH7GLTKPuq+rLYGNxLSkKGDDdrFQSQC9WFgf7KuQffQE0WOMADNeZqt9PM9nhQCr
J3xMJyI/Jq3y/kC1vsKj9Af8a1Ul52Wq/sGVxLg681V05ZnNbPO2NMt2ma04CRPx
IWaAy+yxOVQTIFlWbc/pn/yZIJ9wE2vL9gHXcm2Yheh5Mk1wV975RKProIfXJO4S
AfNquQn7gaSRiKS3GydowfFv47MxP8WkWAp2Gvv0SxvD92pnAARSx/6gKX0JyhCj
+UynCY45ZOdgNzLX/Wkry+Ro9yRedf9ebDP8xCVxuejdppfaiFb63L7gybCai6v8
xqOFJgC4Gg7u3KPW3DlxAL58KDEGyhHuSXU54Fi1OrKxyPYslRNtnFqjhNUUsYaH
4LA5KT5vqbn+6TsTvCDGZ9OezWWrburp2guN6HMl/uKut55DaNGy/kPptiLJh0Oo
nb8rSvY2cag3nWLcfcEl+OPsYUzOhWhdjE/fSgZiUdbJ84tEUQT4EHDbo2PWrXHF
f8OF3GTXfeKy585C4WUjoF1ByHr33DlSeU16oXj4t6qpwRyujWUXBjsF1QHagpo4
g3zYetOpDnp9Sg0byWHyBHSeUifSQ3mInB4ExrPCk+yCM4W0ceH18J0Vn9Ii5geM
oeLj5irmYExUunotabl+0usFPbUlrHtoneLEWJCOBAhM6fW7eK6o4ql4ZqH+M4pq
msACKjHnx4BYOQlZzr92Zj8yqDL9SS7klti744FcYlurr0AbI4Lsezfa9+94N0D6
XNgGHlBscUqIDnKM2cu1RfZQ7RVrWOUidDAQyHDZrL4+HVfBS1Uw+bsjNCL+W69v
KtlNZsXBRWkK9u3GahB8Hv3znnJPRtykqWceN/fHClFRUyP1QOkSmPf8Gm8o+KKD
s+nAMKDPznB4jpqF6kDOGklCp+UeTn7QAsxdHG9CF+gK2qmNN7G5HhaY0FVVwd2/
hRzM1Fz2UoKHIAc6zNcQD1aOPNARV2xLYQwAmJYrTcZ15CS6RhJ6UsmuKyTkybkQ
Tm1zkBvJLC3Q8CLHSim5By92vF4kYs9lALVieAKxDUsHBr3IBr81xkD6oTQd64DE
QfylOrAE7Fb9GyLUzTD/SE53Wd6svI1n+LIQB4ID45UsOGV78Ynjv/Uu94nGT18u
ZW5PUm97jrMQXXEOHwn04bPvNZ9C3OwBm3OEw6IeVLfweVQ9x0YVBdcdgau4oqYD
divdK15TeAZCm9TdcMyPMC2lEnqMLtRnUNoVciIk5FlF9R5Fy0yYzP0RTgBmqMfk
bres176tnS1Ic7Ro1FlYG56C3hlqCwnSpEp2VEoflBVAGrUdThS3f1HBDuLnNGHV
5KxPIu7Ouaej79M/6JKG+6myF/xz79IcLVtjQQ1QA2lrLWQVgE6XKNvFgWxDBdn3
c6RJaMJbEeiF0UuUWaN9gXkt9U0R+dQ5u8rUo2SO44bxFBzGcFA2yVzOe6OJ3WJb
aEYHkMZCUvqTkInfoYYj5P3V7S9rVLTAJfZKC6OF4W2VwnlCmIc2ase6EtFn0/wp
d9N+NMb1+at+1vaaySJNR7L0mFL4ON8yYUsnqt8eR1IviS5ZJdtF0fwgfDmUeUCU
dTUcYKNd4X3HU6rrzY9VgALeOs83nknyHz4nHxLDxv/24OBeDeF6W4iBSnAQrbOf
N5t4pzqdpeNEHXJ9vfokEJ2pc7hEWbO/bzRzgrM7SXfGEKKcPtgIdB97d8R7gexv
EJPA3wZteRrYkQUt6SfaPOGb+ltmTTujmuPNEoCTpToHBEIFblsXnQn3gyPjdY1Y
yKH3rZ+yw71sAhpGlNXFd0aTW0pFOgl+gRYHdn9yvlK72rHDfOLwVU1YHPo3UYNS
/RPLHZqBIvhxht4f9Wmg9dm7Chu6B1ipZphUlN2gv4C1eWpRl5mK+0vHWPhxxBTp
gEiz34mGQruHzG7X0uYgWaG+p+t68/VcBBr65ZR33S7y3zwqr0plMJaaTB640grC
2KaoR4p9+6cZ2ZSu4p5WgQw685m8HM3J19at2Uw0BSYlzT7eaSs1DGk+sMn1Nx67
83ATQmOU2tMIvSlaEfuXjiFz9ySneQQJJ0AXVa4j7Be69CN2vogWkSOwhZXO2BXL
9e8GDCgw26oEj51NcKsFjzKBs91WNIpuO5SiP2tGKGsQTCmI5Ro4KR0CIjr3RL2H
Djeh8m8FRBJGaKkb2RVyRwNrorJAaLCx6SemZ5q8NKEl1aqbpjBuiIXlNImhdSZm
zGr1+KxugKoD9kNQrjrv+RhNA486lt9QbqRj1Ajx92UPgUoafe8xkuy5XoT+iepJ
x4gDPzM4/7FYCau3GDGukaJ6+fW1cyBXGJLvvrS7prkcy/5I1H6YYpG9oClAxVhF
deagUdl0NvW2tGH1+zavF1JCWhsivrOWRrz0mtBb8VhyRr+8tV2lHzQeE6wc8+H7
5t7ZhLCguW31MTDVf2fFbrMgfzZzzdULjq8+JVkUCOlR07s7EIiFSGPuaCpgWB/s
YVn1IbWtSLbx2B9u/V7FINPHLyknpLzeAQHJsDBhpUfmK+QAUmlv07wU085Odms+
CPRPewZWNV10Sfewe9WT3dsx6iQJEIMMnDCCG7j3UFoYl+Cvu1SmrGohrclKl+6e
khuihHw/g37egjCjRITxAGN7rcmuas18IdAgCQJK1YedB8gvQl9ewjU+ASkdXFo1
FLe6oaSYuhESbVUZHtiMGqzQUjwmvSkPrDw8IBqw0PdGr1dmfQT9v1mb6BtceLAN
RU3wHYzE34GCzxqYGdB4kZ0I/h908Z7mGEXzndnfY988i3RR11lbRSzhwBpstrUI
rGo1jSQ3HZgA0V13eNoxkbZyg7J6+KxIOqH3ChO+Gahns9toXY0aof4OOEa2lpZQ
m2KweazsAx0vKRT37z6mlKveUKQx7HtfEcqmVIOJJEf6HhYqBzoIBRm+kMrCyHSC
1zD9iAjSdPdRl+ch+Js5L2PWUXCzMaoxpcGjeBczN5GHnZxfA5urUysr1to7NyCd
cMiAh0dlW+RzrIFHJgtD5+UGFu//SUaZ4Vkj5pZCo6mr9CecRMndBfrLAo3Ffe/t
7Fq1uVRJ+e69coo0mJk7crJD5o7l7xIFXhdcQ2FG7S0qmE8vMdpLkuTWq3XTz3g6
mjmclpAj9GkgCv3Q6i0AUOY1nWTm4Ei3P6hKQ+mioePjDKStuJOjyu0xs28e4xcD
dnY464vDxib3nyAb5ElozKZDHov0TzF6u3BBs0AQTtZrQA7p2/+jZpcMY5+SCD0u
JWIrnL9baLwWDsEFpQskyp0CooJq7u+gUWFEChDcYll+TNqwNs71MtJgS7ZOebJf
xijSSVmhM0+p0bJUmaOILCZu+IlWKYS/PsyZdp79tJjofNaUQFsIg/cIH1WjGqFC
IZzXKBdIPEfn+qP6h0HFpBEe164YTtZG761qpskV3R0cTcdnHb8hNpPm7q1l4tfG
pN+t7JgYH8z9f0eBcR2YizpNJspr6LriSgMjATVi0DkOH7SZ/oYhP/rRtd/Hy3V6
xln95MHaVqdXQKKTB2A8/A75YtjKTTyldlT03qm5UMpb6FJosBpbIsB0nMoeGDyc
mrp5YfXgiFKoX4NxLw8C5YzKgFIRKc0sIB310VbN+jWShSPShJGu4jRrKWvb4+VE
SxCi9flMQiS3jijzCIhcWweBEEmdBsmZUtwm/Hy5i31Yl2qryJwMtuY/KKEE+8qK
hM+xMtbwrwCdkhJ0l5Mzqm1/SKzj74r3KpBQr/0rVcH2DE6Z6Jy8VYPuF/7y1yTT
Dk5Lvz1Pm4XkIIpqkIfPnFSWhPn+nN0gXZhVuxkfRFU1EmIZ4vQ6kH7UbzGJphsx
5DZVFKnd41eDPneW7n+0RGXEei2S1/t7IMxUztrZ5zY4kNxQysw4zVrlWvius2Lb
bEXhQkm3mdqSiqe+PyOSyr4RkrvNyGtJj+e5dPzMr0J7ANpAoD2E1yVRalxXQM8X
k8pXYd5ZjMrgkwkrfFDUtPscPaMZscp2ijHhZwAwk0OxdQajX7nB7qFCNpZjgFUl
Riw2guwLnrStSDQQxcULz4vRYiMWJgc6a2A10lvXDDPuoUaQYsXj3Wn3npHhfprR
rgrXzsWeTKU3gEKYcbKYV/HajYzw42iR75LaqW2jsEzOnXpW54C5t8CTQZh9GZKj
5Uf9drMda9r6WUG8B11EuP4KOXgKRe8LAwwh4fZH4rUQ+chQggtn7336Juav+2eT
Z0D43MBj09RyE/c+S45M026T8PnXjxvJ1A+0Vu7pSoDeVvZhJO03/Vi3RtSRV5Vl
bvrSjT5OSRJ1DMqMNstpwY7ENQ0AsFaD2S3420bsPDnBUdF93eXbAmc0p+pTK4VU
q0Kq4/NfHucNBkxx+SSKl0TEaLSwCaumZjHBEyt3uJVgXoESokktHrTxSgJTYjE5
W3DRpvUdvHj0FSqz7aEryu6qtE8y8S9DgZYOJTOO8eLiYBW6IXalg6cUlGXcUKa1
KDOZi5JlnlKW6xIjGp7i0FGPVWDUUe3ggFdaD64F61ph/10DikvtuVT/t88JEjnq
fG3jpDSUqQ9KNHAPkPyzGoaNE490gW8x8lQ5H2KO7dNWEPSr9dTFt40Yp8N6l2LD
8wHm/1dy5VeuYmT42FfD94NSuvprcHtJW7yWkcHCBjegaeXoUsIPngy4UeCAX6T5
EkF5vPkh7wPdr7oB/VLQugN0zC17dadomQaTvn+xq8N2zpAviDIv8BPQ1vBlg2vC
MTObprHw40+5Mcr5pbuF5HvIfVENjnVY5oQox2B+jIzbDq+CHh2EK50+XHBtSBFn
y3OCnJ989MZo3gWURfC7s475dEpoxrjAhdV0hVsvgHs4jaUjPSvFsnBDAsM4Itxb
bsEFtLFbGgcX/1fkAjrpw/A/xK8c0oa7mgwWPNVk4vkjgsxDSU2+evXkhDrOYite
q2rkvwzYEKBZ1ATnsQeZ5RHhv0Hi9tC0ZRU4OnO+g++pc1b8E+ONA4qFix1wncas
uxv6WSsSh1TWndVDVkvtKBUiyi5Eioh8LMfHh0/hM4r4pFz3VI+OxA3j+qfIt5WT
DMC9/2clUjni33cws5gndgsyH8aUtF2Bsj42Km66H5CnCH+2RyQXiht0MG24XjUg
pABsriommnDmVIySOvAmxHFK/9Z6DKAPDyRWX+nfxSHeJeukumgH9WiOfp4SNy9E
Kxo70BvWppTXLcr3fqqy+MeymY3bgEFydIeNfk1xBxhVWt+f79JjnerRnFodUpPF
Zy9qcjuK2BFlnLe3TeojfrP+c/Ngyl4gqMuIP4cSkzciHd31xYtDuEM8sW9VQ6KF
6Mishy6PIWXfYyNJPL7Y/XMZAqqfBA+nXgwJznO/kKEMJidOKLcMD08mC5Y5YO84
Qe9ag0lfchQgUw9YQbCN4UYkGdqwAUENz7rGtrRzAppX/cqd7u+fHVR/vCDKLvpF
GL1By7aFlIGGJjNv2iJJfJ5fSEX+3b1CRtzx5R4uzJpvZAR4AauTC3mgQCeNZifj
5kBXoXRyOdAODy1j4ZD9YGzf2Z91DQ57ZD6Nnd3zLfQpHwucC29/OUAzA55z8OPH
DGeJvkJouXSEqKRnP/uNVujJo2TnqdZ4tWC5oFsnRdzIJhwyNRbdCnc5lxKEjlEV
evhGJ2gNitZ4Hipnik380sqkaInC2IO508tq6vvrj+4d1rUqeYL1TInA5dNhzkWe
iyLJ+R2fbTGtBwMlP5MZSCL0UlRjlbFDh6P5g7A7mwSfsValEPbN9MMon+tniiwi
aZMhzZQiCPUvc1D4upMI9SSOgA4vJ/jnzyk94/NPDIYXcieqlxDuRkTSOHCAtAGP
vvdAJRomIuNhK2rJPNhJAOH4KiyACx8T2x1bq57nTHQR3/uwnStlRQ3PvASp63I5
z5TRP9bmDydRHTzwb4zpxvskPlGHnVFnqBdAJYSWYERd51dlcNA82xq/CbIKTjAJ
ABP8B/lDchCFpew5aVjd1gDaKI8x17fCvQBIYgOrWd6JMkq3K+RCzec+11cmz6dH
g2UqvNJ5EEj/lrsBWav9GYnxvKFCB5WIAliHM6tgoZIXC6qY0cAqg4E1XezIkxM4
Q50Xj1WVpn8csTtAhCoyVDQnOe4RKXy6ahesJZgny9tHFhzo9DMNPVPiwtfeVN0j
zvwdqnDjI8wHBr7j9jNxUN3Vo792gwgE5yHsVpjavqzu7TMJFUtB+mwRcf3cY/Qd
jYmodIeI5hsat9hmRp67L0Zs/snOMzoN8oGfZTLUtfbw0b5UcVXK28yqDTNPLXlB
Qz2J7TnbXGMZ96v3B8FYS3bSrolyZMGtI2pcMUI3PFSkd0/09FPiRTvbhC9nlbhl
w19tb+CMjTMB+UgqQCrdgMM7Tvb3+i4FkqJjaMTyWzvO51t4eeyypWM3j+py5udc
6wuNp2lcUADcjUctTSBcI4havYAswJ4NkeOxd0Yglsol4idVEZDoPpQHFG6WqxOd
6DhYIIkSbjArV9bl4oQW5Dmu/VsZGUjTVZhgjcNHri0PgqJTBYUVq7Fgiot7EQND
czUHCE23sgY3m8/PT+rbbuT8Xuh/JPkx6RrOxp9rbscC2yc2Pz7Cl0VohYjqFLRo
nhriCx8xhikCg3uZYgr8l+SQ4IvjBhb70k6uK9xL2KEn8m0SnJuCpl4gzHlyDvCF
SdOBkIKjsbewh09l9OkoIGkclQCdQQr2AU1p2GuL/7DRT+JfuYRvJefm6DzHvSxP
Ca4bfckbV+dUwHGz1z1ga9U3GPJrO6D6cwOByQ27NrAf7wJuBsnSm/ePmkV2fnTO
IoEOgac0ypjkXszCx1NPqi2IV2VFixav4ZbPMmQE6OECd3BZ/u0xiJ3tD8LO41XY
oje9IKv0aYAFqvxd0KkABH+j5BcnotNGb4HZA2+Qv8SypmqhSi8UM3m17Enq9TUa
Zbxgoiq/wYT9KTPx3TTTWnLNnD+iAG7rzqEHrc30at4zOkbg7BPfX42rHCq+NJBv
ooCqxoSu8TmTzdHi6+KCGvU82hnqQKDhgO4Jer7YjtkJEY36TGEKk5tfZKUWEG4+
PEhGlrDOYzhuiWFykiVXSh+n73M4Shusvr/K2OdvXCg/UBhfVyJA1iQuE5BjiVOq
LRN8vfaFMdAR5FSjK9VegOh5MIH2w0WXxW6fGyeIE8aUkxI60Q+Xgau/zWiA6cRF
A2bufeBZ19xfh31IV/uURCFY0AI8M5HRoBqNPpI52GcbfIwVz+LdJbw4KDDQti3a
guUjiAEH2yOjfBNmDI9yvI/PP0iJu/XW74wB9X9lw0+km+u/WHbF9c+GkuLkWljy
NcvEg8+otQbGxmjXX+qFkBjjteXCRmyn6qG7hc7j9Ub7qWmH3mGnZOnJmEMWq9M+
KySB5HFCi+GQWNSALSTLNXihPC0SKnggybMCyzjTO7ayjefqxB3fTQ+m+rU8QdMJ
DZ76fQsqVG49y4DX15jDWuXmxvq9/Is3Zj8Su0CIq97I9Kj5Zy2qyCrmzMtdS1Ay
Ntu51tkCQ39rKNPjRLXh7cVwtpG30sErjojq8ph0EbfclCZYvlvT9gAW5ZcAYiCu
k/ckejR6KOQG9hWuAoSREAYtLXSoE4jqeCkquoty8BCRBxaO4bAz/Q4HlDiQSTM0
5FoksVSpFuzjilusKhUJacSFR03hdlp6gVZQHH9nwjgylL/BvPpw59Lsnt/k2wcj
TOErkRAY6SYvAdnNSxCdnKt//GyYWmvEokFA9knzJ5jjHX9HBGw0FAAlyxLSJGgP
rngsMXaVfL8ivyyw9msxXAHDr/e5OZWmK2wkRUCaZGVKFZ6RcR295dGM6uc3HDWN
tXDzGc+SXQvCBkZvupuL4FVbKT8hHQPmOp7dhKOACWTEm1F+e1NXxRrliV7A0+z/
OYcN7OZ/fqV/DSfGHtGBR82dYEkMG63lCnnP1N4cbOd+VW8U/Z9N5AKo8TPCLQG/
XVDXESNYeCfLJiFUnF5+BFBp4bPVGvWjzRNjVnOr9H4mONeHov9pIeIdCIlVTcF/
oXWB6OZezcOak/7x4bR7qgFJrSwia4tmk/EPHd4A0CwBxpg5vsvkerUD4KNHXZ7D
hCry4i+e/XC2rj+ajDdxdH6+9A77D8YsWay7FvxXVzpwCPXy5R8sB8pEiHQnuY79
TF9kbC43AdI8HewSlsXiD8tvtxtMQhngKZG7oSIQKJZhD1bXI7Pwf2XADuYdHLOx
upIXOYEa69DrdPtDys8S8CWAkXfy7Egf+T8ffZ70PI1g3dJHZYawts4Qu0OcUw64
UZKxlpX3TgTGu3j1pv5ugKsDSXBOWf8O8n7NZc56M/NbgiELVD6hdi5tqt7BUthR
obojxY6oD0UQft80pd4PBDcGpgEhhiFfV2nNlBf99KAa43fjisQLr9cvk66oJBVI
QuwKhF1tNJrfkzJOZfbeAEEmg1GmWZ3ztWbMorX7GgtFMHt8aVdEA+uGKzqm2rgE
EKenl5URrNJ1McjhWNk4DM4q11H+j53XL7dqPN1BoEcwbexNuzqy/e/XRODXCmil
NOnFJtIX1/nRizfRw3vgZqg1LTSdjHVhzFncnkmN7dsNYR5r43voR1X2njKCGp8l
Jrr1dX73bsoCdEwrWoPNgr6Zhc8UeWCSZaYWdD8wAW00qAWEZdFnVMZPC4FG+vlP
KJS6qTeBDNOJwKwkp+u1PSxzK1oHJY+hTDxjZ8GKEXlEl7/1qklBXOuzLsjH8P8c
iGobLuQ9+x1cmhUSdxfzwz64FDznyoW59Qz4yrhKPgBs6y8ZqnLIyybWn3Ny0CEg
W6oG2xE9pgt9TzsH9XnsCnpohrX47WTpnctMcKtfJdXsPgcBkM22L5nHs7DC3qEJ
+mJoOghGamQoCstCrZ/0f6CPeqD/sbT42YlwGZ6tf8UBtodNi6IN0Oeh96St2arZ
XpNPweiqiDjSl49uW3t4ukt0HhY0eQAQg9wX9jtxBKX+p+LK2XBvd2MzvlEIENTy
27Di1Ji8OA3tSYu1XHPdthvEyxryWWH+ZpMvcGqVuBgHniMPYpZweO71k8xZ4Ek5
3Bemv3yLwYsnp6q5DIG29P4mzZFu8Ky2Z4IrZ3q5wtXcSE4ft8qbn52bkU7a+xWd
yYNhu/GXEVCind1BNdvoNIgxy3m/RhAA3uI4538s8XDkH2z/Q8SaK5LFIkVMDqmB
GYnBfQVj9szByuzDphOq60c8ytx7ULIlTRZLPfYwAFEZ7ZUIwEDiyoYXdy4qHWDe
y8jB+5uVKAK75MonrMgb3QHkvtL1XyvpvCUorv8uJ9lgyEHN9uCscae+a3z+QNnw
uECXT2yT0yEOPYjQqRlIbMRNQU7xGE04M9qkJ0PvcqpjH0xvgbM6JJ64RV+fQsf0
4yP4iyq//VPdUfS/V4kJlYQ9I5X9DknqZmjEaTkCPVBkYZhDlAitQLFrFid8ax78
hcbJ5JOjYA3gXBODdzIGctaQVYY3ky1ntOXPfcXRhGfPWAKjUe/3FYc40vFdls4f
aKMsRbXd7g1D2kOvjUMh81pqp5DUu9wAgoEUVwVQizWCdsySdyhbux9PGeW8UUN+
xS8Y9nONKFNHY3hgQQjECz6X61ttJ9HKes5JJ8JVtyrtzwHlqSY8ug062A7Gtl2m
sS+PWJX+ALUB/ksCRH+7SvBKRetTmvfgx4ldVxUkoJtHWDEVphCsCfx0w+YOhE/A
mQhhaa+ADDAG1ki+u1EzzJpN5s9lLsI/2X/T4H2sWhF7+MXrF2NS7NWSX6KoPmjT
OGc08w7xWvMStNF2OYdHvOlJpqaiCRe61wV/XWmlZSqQVypu7AL8UMsrSzTJRShp
JVxf9RhIV6kyEILmSq/lPtjRUX2JeDGUUYOOPxZg4hoh5Du+TXwpOM05xJ5e7Wud
CyTEcHu364SsTh2x0EbAwZlS/ZRBt1F0rmah7evCCpa3Jgu73Xbx+l+RqhIMUYlq
WwHw2kqFY2FS8L2spqpLHYzyMB7pFNkxX2uOQOq5F02etgHGIXhxzYFRiVDLziMQ
km61xgnKW2oKwy9ZTI9D1fyFN19UPQRXoiZg1bEzlK0M5lGvIgruFRLYM6AqJYhW
JHyUslxfxs7KYtvHNxY2IXb2pPL0rXEQFMk7hFmEkykggsEH5cPqvvojt+UVYHRV
tyL5Z8om030KFB7bFlPJaZximr4eOheo+W9GwEy+g+TevfeMCQzJqWe4ck5eoFus
2d9OmzJXAhcvMuPJ4FW1jTOGr8o7h2G6PYTSjw3M/pQZczhcnBn3VJpFeBTuUy54
9tPsF8c2rQgzDO5kN77d5c4USTAd2qVdVpM9YmYbUnK/f0kti/P3yGSH6ccUd6d2
V0ed9O4lI2SmK//FVC244LPog7aO++Xn57KP5GSWjjK1/HA2whPOXwqt1cZpVpXv
E49jJXtAk3d76fIGuhvNijAqDMAmVdUSBI9JHc4jHvDKOPf2srkbUar1QKXHMHoD
cKhJ1Q5nLrNeR//OLF7pGO3T0DHeGgLCuE1zq/sdV+Rs+sMzhomKWpog3Pnc7gTe
bHYy9cM40pJ2vMo/Ph9eQbSoUxdveA5N4ZSpQu2Zvje7mkvsETfLfaPQGCzfAr2+
AxXJitjvnMMN7a2g/gwTiLVxdN+Lt4fKHMIakUW/r8Bgjvz5s0DYCRkqy8HLpqZX
VBbdZ7nhrbILUQ4z7M+lisrLDFXU05aveYrSCqy+eCJdLhy+Q6DonE+zRdOyRF90
PrTvKgwTa/AZsOc+c9O9sbLvsLBgHb0CQ0nA+LFC6mz9Y0wl0gRPtvQItNWr7BYb
l665yPMkD/GgTYkb7G6ts52bge78nL3UC4yhuOKd1AY2+twpO/TpwJYAX1OYXEv6
zG9SEuYMKNuB1Hc4uU9yX/Y8xKR+UMzY23SfCBg7F30lz3060aMIZf5lNQ1GLJ5B
M8IakvWqUUnhzR7PZzffMFRz4RIg56lqoVDA2vEhXuUNA3uLX6lL/9/jvtgTYPZj
8RjgYls8vaQo944ws3wFTGND1uq8bRuBThLSy9iSSFRQciE+YYo4hm3Ui0ctZ7KX
Etn6mjMbgc2IWguUpXwIr0sE1vicB1+5JotnQhIhFszcpM2R5DKP0WqAcaSbRIg3
Nnhtjv+4McMIwMUsdQV9A0jWyi0vmprtSbVo1fPtxiuO8HNLyG6JRmmfM/gG41Dt
//lyJwawVbu9a+26Y/ydYS/PqsUdvDcCLZZRY5q7yszc9QkzzUhqybylwfHqQpRq
IiEXvZzEHkbums4ZhODKmF9Tr+dAMpEFXilgm2KRdjit8NLeHFm9JlJ+SrcJjZCD
aQd/PDbBnp28K3PlmChsOXVVDQjdQqiOUSWUWP35BpM+kccBow1vF0kwmp2JR848
RNNwO/6DH0URx8Dif6MPe+v65blv+i/l+B1nLbGesk5JNrsUe+YO8gGBZiRfW6M9
LrGlbTtIdZ0FMJfc8wBGntA7S8TdesJcwSJgmQIQFv+zL+bTcf0Hi+cBjMW5NsbL
QcnkrbWNQtXqEaWMkG9v6fSV74Rpm1K/B8Amj+M0EVqb+Ym3rEojcFsTor9lev1K
jfvCmb5jlLupTOHG2NSg+XbR9doUEWENhg97OCvmzSSbx027hUMACjr3k4xGAfEn
Huy1nu40sMPr7DFCcGZmBuOhH6889WtxMc7VKRsnZyVRCQLpatSAsxJ4q5hHxBI5
0M2yZ7E97SB66nI0UBSglBmLBrxQAjXra7BPaynEeKmGA2/A8pt3peQvGE3eMUS0
y3u9xgtTz4d7eqv5IS2gB8SwXDZb6g99fQkYREICvwxwftBE7tOJfHAhMg0YBE4p
NEA4lVNb0hd5XjvBWEOdpzeMCS7FeUBOhVnuI7Sxczfk1IDBs8cOMMwURJ915OQN
XtNiB9B5BDh4Adek42SSoGG/6GebOkzcsG93zZOYvl5LNn62lcKtgzzif164KFNK
jJVV+I51qnLfLYT3gymSZrKauFO0JzWv1J3H2ZxMuj+UyNGzn3RhMr5yrta4P7rp
pW9/3o0aoXZANkhuv4PCbwRzeg3FzERP01Z8rYmDIFez+c45psQ8zXw2MIBIRDKC
yD8xvTCuoNj4KL0TS5K5ZnpdXaQL+6p2GNP1rr/tRJthh8h3d8mCB/6B0u5G+zY+
3N1hnfplkYuWjrZo7FjkiqjGLOqk0ve3bSUwLsTafKQgg7c5s519RHX6Tn/V3y+D
a4CzV7ITdvXKWwBY/zu0bQFUWPIas44AiGcULxVYeZTVINtajSeu0Opd2/iHfsBS
+/jm5gWNzIMnQIHnCnhnk0idtiJPHbBzMfAeuxWR2wKs0u83Owe9QqNysxdqwlcu
O3vzFmQZ3rDQBrgsn0it2RoHuAnfM9ensIi+jFBrYVMW3G3g+3cyc8V1NXCQpmyv
IWNCS8K/WSJoZ17/pbT6wPLm9kRgruXfjaBq3mxkpuXEpUfTq6Wtw5VdokAJvePq
EPYsJy56r8HntUCk3nZ4jqx60ywsuWEj3lAtH/HDqDRNjaBtzYF96grz8RbIfsvI
ReCggY6MjncLc9NffZUexS7p92NMyrgLUMoa1WS9IRiVniG70d/Mr2uNwML2MsLm
Wv9Metk8JLmlZ1IF/inicbF6mJX1mgbi3gqaECErL23GbzEnUsUwBqrdeZlMTaRD
jz0OT8kWhZwZUBtUSkUWNxlUZ5tjQ0SCDCwYc0EziYXzHQL9mydDeJ8Osgpj4t1f
ElFBmXDuFwlBncrK6anPXm5YwefkEQ+pPH1N7qd8XyZwOuN9WA0pQ8h1fzFZSxr4
XMnjoLk0BTzDHx0r6Bh3TUs/oeqkrKRIcOBy1RCDVkiCQcMhQV1DNPRnhSkiVt5z
91fTP+opQ+IEXgdgrixJtTpCku2SdRX43VXJz+Sswjp+uACJnZGzbzi2g7EV2tJz
zFSfetXu48ON5od5wWIIS8EhjdYfLISqV/Tym4gKixj4Dthx7MWuehdUGno+tDoA
vDmrIr6Dumhs5Ytex+4iN/9SSJNexgP7x96lR8LCXi3Diu9PBmmIJmSoWRZWZDzn
CNYmcxawGSGAbi9TeS8iiAu1q7Ca48VlYpzGxkEzSJ0AFNreRl+MgSqPBNLAG5vR
6GWC4IrZpNI8f8HI4vtkT3b6jS8KNGXDiVhlWqoGO//0eetezF3gXP1key7kSOR3
rtEEw71GzHBy3cP/tMgIzGsgILFLaRL4aeLOFINADs9LQJ1+FGKufllxh0/pfq6j
ntNTc7FTps1mUgzTL4lvB/4rWmyGU9a6d/R+HS0FhhhSFE6kX7K9pC0DbESR/4an
1NPPk2y+/pHfRhlTYF4kGCHxECIWM68Iuq67Y4q8GRbmdjCeibE+iDE0gvMU7sEe
QkWs78FHuW+DnmXbX/DjNbt5kh0nXPE18sQ/s7hqTlVG/WUKc2+mjlkTnnvO5m4P
RiTXBJJ0aFEt1oPTohlC46Aw1uKE2NQp5LLl5v514mZQuu8Kig4/YAMHwH+bcFnj
6hMbrQOjMowjtMbQ09BGeLovvgYRPqfFIJZ8/InKE/NXCywX6ZGfcLAAdhMi9vYR
oxcRTHrH3zWtNqdGn6Kgurdv719nKZIIM2CdN1YGsOR7d2wkJrtM+HcmwUWfbaFF
ytQ6I7yBxTaTBavLsJydGGvuf4w2K+agQOYOMSaGN2ljtQ+t7o20+FJo3Jb8eugO
90mlIYPfbf5g4H4XUPDUuW6L9foolNyHKbT4YW75KSRaWfbBES4fk8+HesVuzwyc
54FI9xcR+8leFykoXTTsv40BKH9JsbXh5dkNIN0viB5hqLRFYv8Aj+jSvzVfs6lC
kfXNMzk23Xehv2FG5S/c5w3smfE5eXfXSFSfXLBM5mKzlXUmIkfhAnsba9YBFifR
kc45lKmV8n+KogfO0869Y1JGK2gPze2JK7cr7yYlw2j1VArCDjF6jSydUFZA2Dtw
ntLAskxrpmG14dKc0YPskBvAC4q+dnMG3WMW6edawLnQHpQvmVe6BbdVG6qcYLua
vqq3Kiv260iRNSXXNaX55w+hX08Qu8KzBeq0ZGv836dthsPqzpx0tBD2dy1gm0la
aKszwCW04S5aSSG25wImXC12GuES81n11Giyp698FWaosxKsYk1LIBvR3+kVxuyp
KN4yOYpI621FPNSizYmPQ1g1yPbmGdFPUcGQTnmUptly9HM2K+CSHtvPWqoICKUu
yCPeeHdJqJqjs8ezztNQb2OX8rnHnNmxZNZHdF5BVgM2hH4diw4JOIHdMnh7UOpV
pc9V/6aOc0f2om3sHOf62E/wn5AET7ukc4HxuXY/JllYTBu8JBTHnnx9aRu/boph
wLlFcLfTQ+HZHfRW4nKa6L3RnMl0GzBwY1r0YkA/BIUwNJMauVfnlZuvcKJNnkvT
35C/OeNrQ2Kii3CYwSBLhuuoWfxUUgNhaUIejByfoo5Tns2gFOEHrcFw4fU2sjPg
yvNpy+qTn3uaQx7Qf7y/qjL48kWxJtzZAOIMnuX3ym903EzUCHXzJeJ6HxyKqEGl
vuCYqTMJeQOYyZBIH3IUaSlrY5I2f1aBaTPGVJql746+npqwlnrkpxd17FB3DHAG
unWx4/tqMWQtiDNfg9q0kJaq5Wvu/+xANEP3IlkJiNdZ7q3U4hUHSzcNu95Adc4k
4evN1ak6a+bXkOAMKpYEc16wXFhkq3UbK77DhhDjYakYV8cDu4Xzh7RdLm1wvgS9
sN1EZuEPjK4aAx/YSlsVYhBGZ/KVBEAkJd+LlwZ3o8DPlbOLrFldvg8JmOYn7KXd
NRUDNex7v6nRLBmsFWOLxMxW7TsfrTSJ/iM/Dy6dSyF0XOqnOKIWpcF6wzCyE1qL
5WgMUIW4t9iHcyeVE4dLsz2B/gGpdRpr0+i2HJ2ObX5JT1l/ZIq85Y/AjbkRRamG
OnIZTW95W6nimFN0E8vPZi4W+iUm/xpNdSUojAeVD/v6NHGXpIKJ6PdTCZdigaq4
KbsDeeoq9PvNwpq8WgZCBs0Il6SGXb1bQqfDb07FwC6Nbn/ZdMsHhydiI1wwwnNS
4nbJW2+KhhXYIxjRR9HT5j48TOKzKF+3yxEuiMbqrYq9nmGRPtRswN0XtQ1H7N0H
epO/HsXwp8AG8JWjy6zZG01ad4jyEjc7DnRuhp+tsLAyl7DOG1L8Cq+xlcGStn+d
5zJ2KRQ6e26uTHQK7XDqwkkTuHLCjzNb4QCggbvR6EEk5wRZRnWAT0aFYi+kE1CX
F9A+EzvOqni0mJFsIDyMQ6+MKq5tPhUcOIrMsykfES/Fpb2vWdiAv2vgIMjlSn54
tE/v13Y4LnGaU3lveiDgl0bE8sFwiZNRwH33Zy0dvWBxXtIr/75eZ8cVad1yz9OO
6/uTi/quGK64It5aREJJ0L1Rwz1/+agoIVZ0xnfR4o9lIkqyBaiSnHMI73lUc9KC
W4f0jXJo9gT5ybokSDA1lb9GKExbrU5PD7VAv4UVSyNbvOov+y/AYbbOMdJ/W+Fw
52kLSMwCzZYL0tAOIQi5nII0es62JsBa5OchbLarINJkjx8QBuxCXaQbYAKg28Rn
F2fVgRtaG+eIcWnoKVsgSpVulO1of8TSGTW5MGZZ+6zqYFdeuz2pIozd1XzaNUrX
Wyub+Yro6tyPeL9QzjqzaV3aNOBsfTUBQT3Fqdd5pWV53pqYUrepMnO+KKNoThK7
Rpb3LsiGK3iV8ziwbzWCjmyUMqzcOpNAqrihGFO9331Z4gaFamBuJZGNvb6mDcaq
lhWc6QkSXXtc4JEhcKS3p5Pk1dMhJ7WgmuqqdRBsaaKnSnsUCy73BOAl34aIRE7M
8p2ThJ+q5x40mGXaoYUrifOBwpctGskHtCxXjUS3Lg6ia4TuUkmWnScToPewpIod
T9ogrO2/3t8lrYrjr1uD7pKyAuO0yGYPgBuiKAPGXzOkP6N7AvTNgn0XJtN0VZhI
V/3LJ0AXe5cq11h8qnjO71GVFsc773BKJOUw16rAzaZVAOZ5FzsZ6b5PaqYd9Gmx
yFaJbM1XKjs0eY2nzaqhpN/peaG+avGB/4MxZuxl1AcIU1IMR40FflQUzKysF9ad
mJUTf8WOmALvb7llJxCYeULhP11XlexOsDx1mt8BXeDfiSvq7yVFfcqzJhcAG1xe
n99cIRmpKpYAdWRSCiV15WkPuR58w4zYIA30KbI/etIGNOjh1HQEneylg6QipRLJ
W0Ed3c9SKqRkeNMUP2m705BySIgirrJix7oxUfc6IfbXpjkybqoA/WPWdtja0GAb
+bGH5zHXnUniP23114vwGzFrC/m5QsVY8ORa6GoMRslWrqL51falc2dnzM2aRVcx
XgNA+F9MFE8WJ0hIWf54NDKMqXj4b8uD8UY3vHnIILNnB9uUCZcOMAQJpql3Safl
0UL+UrNpJNJ9x9bTy6DIeIJ+9vBSxLmgk/M91FRhqp/eHNVD+5G2P45xzaoxyed6
Nd74VXL74FwMV14/w6QgZhGeYRJQXcJhbOISelXLy5TQLIPulqpMilsnga6ZwthA
Q/tNX/OQSgfck/uysY+Da/NwVyc2n+SmW1Gi+M6uv8ZYCaclhhBMkAbz79PhVDUm
Yun5nD2xjWFTWKonCEst8jGgn/zVF661FXaKYIqxBUqv2vMrztZPYzNCUi4+xiax
iYPudPk+z+pCLR0W8L19lBL6rWxp1e8L9GWfF2G3KaOm8FxU+wBA7XhNppIe2Ptg
8efIqPU9kcwg7UDIl4QmEmW8XL4Za9EQCMYVqo025BSLCZwVl7lPjFg0n6vjDGGi
gRrX5Ke6Fvib5UvpKallRkjh53EbXdYSdxjhCoe0V7FN1Oxhu6i1x8wH0KXRFbWh
6Ks0NftX0v1H6jSMBuSq2CvxbtSJvd0Lh8tZ8BGA9aLHNNUqtF94mnsy7xo1/Zv/
wQ+qSfPsziB0RQWYGnTGXkFg1QrnARj4OrO+FkoUYlvA2uxQyu3aNjwOzH8MyH17
X8UKERDdh77xfTGnJgkX8vqwFdUb56+7EbtkvfoxkD2uELrVnVSNzDsEXUyU9QlX
FrfY/9Jb2ypJzS+eRinc3SNT8Jfyx5KPKM9K4oLk9AQpjqESh1sIk5sfBE2lOLe6
ZRunHLlUACTUHRRONKjqDlqBXnVnDu/l/viwrvxy2esTj/AqatBT2a4ojGIlptJM
QQBZ3IYkmb3VQyPNbq1XwGqrrKOj3UMTzxPBYtzmJXB0FPZaHmme1o1QROur3g16
jairVAM5EI9++tWFbJHEYeKnDCvMGxLMknEa7gv9VH/ciNxCQRxdMu6c2aYpR4iq
VIdLMw/prmT3FOpqajeF0/GjmnzReY8xB0HuhznW/DH0yASE19KAFh8mWe5fLi98
UhYOPuUS0vrZyYvk+0ViBCo35sZvoGVs25iXSkihFbwYKggYF0blRp3aD6qyg2fM
hYoWKLJSSODq3mLQ9IWxG5WXVigzq/W6FAp4qyfNAMN0bb0iJwrYQ/l4SYlahaLQ
C3RzJzaw9+hwRHzwJydfV664le6MXFNWlIzfgkAAXjnSlEDdngL2IRoBvaJTfmw1
TWv+QM2kVNAX5aSsaQNoBwmFg4xbYJdMqlVJ6XfM5G45lbxfTWyVoI3YDwE2EUma
8b5q05CaFcArovYHUKgbv+oRfYOqFWc0BHOEnmxGGsoVQj8juZaEvLEfwp2jKrOM
1jbG7HooR1iXyeGjhReprbmefEYzxwyhBz5saBZj/eXLbNrZJ7c0H0uFIrPGYzpF
cyhHD11t2ME+A7Awlvko1dW3K//D0kjxxd26NH5CsIcqmFtMkr/LBWIjrhVeP/ZB
0aiKUFGWopp7lCCp2wKT1GY790p9mKImSFQrpA+Q7bjMXq9LXFBhFND8cGtfOD67
7vHIHhS1ggeJYGSIh4Jtt4/mXZ7PKyXyFQvR6L5tMBCMa0SxmVGn0YnABR5TKlu1
tShcTybdavdEqFXk66/191YlZIfNXWCy8ctaE2iGqhxuGT0ic3bqlQhHPvjO31Da
f8rGnH9LNcCKyNQNmj8lfSTRgx0hn78UcOC0E8kdUzQ14SA/Xy3afmRP/m4FfPCc
ZUuLfAcy0OvMKQUqLSaLeDg5o2SRIAYUwIITNxsfg7gEiy5YCYhgzVQaLPjx2iGg
B/CL3cencJA3Qmq1J5Co+pjGE3YAfHGmAzTTNXuXGOt26N6GrYaKA3MeYGsv2XiO
rHYSsnfGmLOW9cQ610M/scdLkDqMnqqeJPiefpVmh4YZVG0lXpDIpscvG7wVo11e
ZteMo1QVyRnDmpc5ggSHYsYf35+p75wZKD/eWdG5Oe9nrlSHkY5Yaz6hsXnjYLQ4
s1AvoVMAeF4fU1KztS9x2wBuv3s95uuyKBrypQmV41OpS/4oaBcJ3MOnZWDyYGTU
0qusSyNGrdDmDTgOb8V34N7kljwd/aRDUyyptwCetAYlX0z7btV+Eggud1v/tZnS
oQmXlHVDLJShE0MC8ctBee1IpWZIMb96l6VwqHifrPQlnz201MshefUQJh4RenIp
RUy/sE1SwXRjKFTgPHsvoKGDJF18paU63gQdv/6y9beyPsyw7lsHjtX16c2dy8y8
yzbwjXpExh8p8RphB3wjUWaWOb+8ur6ujxTgjjl1jYwX1UAs1uoITAkT+5LPRjFG
FmO5mi09ijcEttO6U02GTY5RIfeNU+LlJQALEhLbO/poczdhj+sVW8GHLzZH+Iop
jnfSd43+RKQBVehjdsWon0O+ZXBvp4tlas96go7OS6//e0icD2PDZ3++gBTX0ur/
bzBOMUCqbVCPY4LTEGgOri42AuxA/5GA71/JKTwaqDzy8jNsuyf3SXJ1dIy4tghk
ILcvxKURPXg5a9HciJDvihNm/mXSwWHiBP9xxQl0Uypqsk/FX2yC/JrrSnMeiC5n
0f9WI0h1zzGdI4ggXsq8vxQVix1YJxplTvnBPuZzCdqWt887/oKwCFCSlB9o8weH
JW2gROw9f2AM5gNZNZtkoga5Xi9XlNNj9wZkssffbFkCDkR05XDvVABLVOvBswJO
jetjPuQaxCmnQlNBBkkei8IY6PCpyKp9w9Gc7dLo5Kuk10GZhVEtIRiDfLYJTyE5
tqN1od0Xn++nMzff8sKK25jRzbYehkOBe1LqgidglEfr5II7wdIrgL9ReAjY462r
cNoGVxE0jpNDkIU/875bgxLqZxUnCtjO0eRgxh5SLhPj2IcaVbUp8vNzmnSqs973
nm5AQRykjgutISDZ4T3r+eRGsvAfZR6J1/RNwYNIvIa9XdCEOLyKG5d2W8MTV2Ps
gwpi2FjPIZKL0GnzmjcnoQrLjllpPBtn1jcnwB7d3jSMvraZ76cUuOnw9eIW2lnk
/QiwrXBuLKMk5gAg7AOg+6MKlV0LjnMXxnbfEEI09o7/iZmhckMbWW/dYW1dJ9X6
hpXiZsC/0SG90usjX/EEE/JxzybhoMpFcfIjiLJAQj9N7vNllmek8hzfp1hdvbsJ
aEaMxSW4svmkf++FVQnT/sq39eiNuTt2OoMXw0huS8qkye0WfNJ1rGVHfkx3MyN9
a2fc0CKetAPSVumJeBskzMZnfAiQ5dHaC3xa7obY9bHQRihIcNm3WoQYGNBA2Ulj
zFL+PxCNx6QDkCv4sxn6y1HnKSEfbcgI9CKWXDz3QF97ipBoTYoJhDkqKbfm9i5F
8Pz83VHxPZmET7yuG/capkUweMi9FbKDGM7eBzKjSFll9ARk2NNaX7fHh7Yg7Fhs
zGBqex1H1CFF9VtDEC6S6pRqPZ81iGKk4nLr3WknCJGm7oSTxyfCklwz2v4Do+Ph
6mWUxqrlmsdlgIOycho3J8630pvZM0tDgC5ZzTfXQBkWt3KiIDoJLd/0REl/ou8N
as1RPnXbKajME8aNH/IAuaZej8BmKfJI4Bfz4IndGh+aVVCfGs9sHm1pNr0YimCw
8cMHV9zMfRenDldLbqoNJ7abXH7TjVdQXB+Ljclha0rcmDqYkU6txVqINQkbL3rF
CB6CZAfLWZWkE1GKKd+Kw6RnXlddiE62ok+e1CuIeSeaA4VxFHXphwZ8Q/oHJ9d5
neYOdDyzuJn/y/3uhf+MuP7FdsicJe7YrQA4HEI3EyUwwKulQhcl39rzoyCy7lMa
ti2f2q+XpghL0a0xHbrNzrI3Jm72NRYka1ae1t+Q4YGAABqf/N447bXCE9+m2GQJ
3eKxzcCcbNxxDx/Z+xOnp92Ut/AyCWisPW6w83deaAVhc8EJ9FrnPCKTGXFtlhdO
04fXC/j5tXjDsT+3LAiYJMFs9MT1g9AdxQd+cE6sTeH5xM+Oh6az4hMkMJw924Dz
mf0IbqUmJK+5Jn3Kb8FxFFVdYYQoH7/kUxSQ5TCLAm0s2a1KzGKeDFfppZuPwA0b
RfefVm7kCsjn620nGl3CVRjFAeEB2oroIXd0artyUToHIfUSeI1ELaxenS4fD0dJ
Z9C3qp5YLaiCCuMHCti/+Uou7dXsORaeVhgvavNszF0mm0eUaSOS9w6ZKEhCCEw0
57/90Mt6APBaoyehbSIASFxbPYNpYrEGwaVAzszqnItXwc8vxNQrzuugrU32tSHg
FjiZ6gp0PPoSrUImpxgtfTPbc6mw8ka6HDp5sF+aTVroTl4IaqL0bdCBTOI/Z6qO
DuWX/Dls0SFgDdlWyg7G7D4IHFFhXh1CZ02hr5GfwZbWXZOQX1VdkMew8o+amBMi
Zw54gdPkjN/R25iT5LLeH763XfZwBAUWyI9+WqltgO9v/1nfLFcL4ZNnv5zOHGtK
PFRM0jSZgBRSgywRF/7Jcmx3p7RCTPBP12bb/kXlpFuED1eHv6i+TklgfFV5PeRr
sLDgToi8czVHfMb8NTOtNy30eLQZNElPsYK2QV+sh4ZAuqe64W7EzjJ1vObXdQfS
ZN35bfAxwtfpF04PYrG5V1yymSnYl684wemoGUFcuxXup4yJzb5jxdMk7hhSAlpr
ldUT+9AL4PPXPCW55fF0kVTheaAv+/FzRZY46s8/1xriRKWVbd/Y9YWuAqAFwfhl
X7kpNU4iOiI20HsHzkE3I6ucm6H1K+fsD/txvhcvL4oXsv7npARSJdUaXHQZ6UxU
K4jHxyj8+NQwz5nudEXfIAr8Kdl1KBYQY/OKkyNs6BTOotRQ8w2SQpkMD1D+f4uq
BsJ0UXHGaL5uj/NnHx8nPe/8R4To/ydiLPIPOtEzXsYhWi3lSImJKtVWJ5vvTux1
EXVti8yb/W4JrHH3DAp65v1FwkMjDJzUtPfi0yf0vTWGj6RnOGFXtCsfdfNQw7e+
R/DWFgzNQTs2M78mFa5l36A+yRvTY+FS9kQYNpCSGz0hhDpZk8MrtMWViGV29yMa
rjknY4PWMxBCVwP0EClZzIKA/9y0oUjj4h9uMtEiphc+iKBIaZHw1daYuSMdbcAk
dE26q51dORPvzTb9Lwx+LMlqcMTPOCMcIUc/YK7lrabThrvcFPsZhuP1mTWxN3Pc
akLdfr6mA5lZxFWykKpyhV2MV58hsUTIahpEgfVkq9vpDwpG6iCZmLgO0IT2Xzf2
3a0ydg6v+XYioEDDw7NWfxjxHB5Is4b8kQ0TtKAw904xiX9FuRfo5B+SGe9OkfVb
SK0MnEnk+B8i5vw1jzXOfCcheqEfdGu26Sov2GKDdgz+SUju9HCE7/Es/wcRPPay
p9EEc0PKyYUdOXp3WP3gRkHL284GaF5yyLrDO46bQ03MoigFwMrSlAuLGZDgoE7v
Zm2suW7znfuOW3xRgRMW1JohaD29o9jH29wbBj0l48wu3HlTrhyoXsC1gtkcHmjq
nzgbaER59mdYmPqq/h5+D6S8p9j7U3ycnKqgJyE1eUc6nb/Fz8xeSjo/dowK/LDh
RvJMcxmWxtXBvQa45c65ohTh1OgXtb+rWsWH2QnJUPfBUhDc2Agg8GP06umwvxSH
a23pQM16swzpiZuSqWLg4aGFj2fQ7QStZ8vEVN/QZnV2cJ2cKCRjgjzQzd8GSTYU
Lf+RopfG8UutnPStT6tgtHJeRl+RUZRMSCHOWnBOPaZC980+d+15z59C5snZk+Hf
aKq5yPV5nm/j+8upQEo/x0ah8GajDhrctcj/wyKsMmj9WHXP/v4kL0PMMQMqcuPG
JkGH6yaAR4CgwbwoJf+UzeMrQhCKCioyfqkEF25HepiKXp+47uTuC3ec+bLkGE+P
y1LnR9c4EDTqOuQ5yHCQeDIPNK/zofJLvw0XiIOpRgAjHumsKRnMbDDltXkyjq7C
9IG4B2WIwg2Ec+79mpM34ec5wem7rHURy1iXP3OeIBnQlqKUDkJ25+lEayFt1FyS
YGUFX9cs9tamNKDYVMog6Uu8azg3Rlt5U493r9P6xlHQdUSaxJ/vsyGvVOlqoZ6S
TpflM+Zc1Fx7stuzBuGEuRFt0eKf1BRyRndtDP6VOSe7gke0qmfFwKXwb9jAhr7b
wIWxf67J4CfcM420DhMCFjp8PY3DKtYG4qPlDeiYZyU2ZJ27CZOpnq2HBGJ6aRls
8+Ja4f7uIpoGinGkdLQTuRIGfTlUc3aOJGDbmIRd6x/28dlTGZ6EQkwv48x34724
jbxE2mYB3qyayU0dwA4S+w4UkfKzSEzxetXbs32PrNXDhSU74SPqJnhu87Y2KMGc
3sE3ftOya2pocmNeDznJYbgFI/6UrrkRGggQcG8t48HxNSY8bOBx7DDEpMSQccz8
sK3jESUMJgDxAB3KCopdTaziM/g+cOw7faPwQru3J88hyXaqDx9MZS5lF48wAjIF
gdNrGkFGT2D/x3xW2vv6OqKifbzogYIZYhsWfsPnfnspfBH9FsTJaIHZm+SprFJm
tZJfTnq625uaHa29vxItqSzi5ZSfrbYm/Hv8TMQMWxJ/w6aaKVWIdVwAsnbKCrwG
8n2b1ThLoe8sM8INYk5JiGtJqCKeN/33ERPueZ8jjcNVhzxzpKtvuKNbM4Ccv74e
c/oa9FWNPFujY2t6FrfjQoN+o9iBYIxv8jRd4744ISQcBFXO3gV5rD7r6IXCb4Aw
auz6A6OgapSr6/rRhzcDK+zQiprgPu7wxy2znK9R6X+l9BHr6kWvk9eT4m0zbPsz
gjUM0CQGPn5oyH7jGGJnySdFz2fmiFBm2HzrImHcHP8i33WHAsQOwkCuDMyJpNxF
jdEa/cGzJ/NuAIWPNB6b2jZBiXuutmUAkMuIn+MrPAeQEWv6zQ3DVgFgnuL+adnP
0OPQaXAq9S3DTu5JqG3Zb+Un37fsFemRffLriX4u8u0icKM/q0YPQt6kKsabAWVG
rM5mI7SXkQFY2uIa2KBcsDcKxNrkhmyTApcHcf4+eyHnHPrLAGa0T5hUxpUzk8jo
X91FYRTh1LwTIk0w2Cd0K1mbgHZqrNt4DnpBGSuMmUy0lN99Rg9HG4AJuioun/nw
hSWyQrfeGEHYk9f4jilHvVljRyM8viPswsfDCEC9n6yz4PR3AM3H5gvc7eXhDRCd
VuqYpQSV+Xlde69Z65tlpK3u7FT+mVF78HB3owM5Q07JS2pGKKKoA7uiYUw2B4jS
0GfhB1vu0hk91YVjLIo3HBibrQ71jkdPKpU8CrgxxyOzEVrv6BUpFLk+Y4O7QyI9
FYQ5/whvRmlOlbaYzi5YlhXLuF5DgDeWK4/ciczqnZTJZMKtV7zQVhotjupC8KQE
VYTnUIbmGHPa7HErob0cl18gar56x9abm36cKlRSbdDnY16ndam2lErNOmbN1+Qt
XNSQMu6sZClmvmXoeqX1+Edf+0/ihmcQTJVoGToQwku1qGre4l3CLuoRt+EUtcLu
57uwQiLAnV8Ax5v/x6NW+V5HsadH4aYvflV8WzcYE0HvUFByTbOaof9CSN9pKAQW
NZNR42giGRKpQDrwzmXhpH0mm4Q05okM2z2xD5iOL9Kjgh7Q9WVpr2v3OvD4s3Qt
nnP+N+PhO97O+ozlRJhb4G6xEjlCBB6gPrf6XFDE/KaPvsGVPPBXlateEuFkLV5f
4UATdZ+nfx263fibmx8+skDLQzDD/tKvLj8eB+I/Uttzjkch6z04Zxl43PubMwTa
lndyZinNm1bHRuHASr2iKmRljO/r+KQ0O7DVVBVRs64Ol+1MPKTsXiKBYS7woS5C
54Q24/Y2qKsdj2jKSY5xek1/CCvpb2Nc2OfnaY42Oq5mY83OTJWyLesFTmV5+zjG
JudU6kU3L1FTwBJ5EuiiTn3i+BGZXuPBT2mKYrClmVXo0dsmotXduH/DtgTkc7WW
9cAjqFDmDCTSanr9n4WKEhLZe2W9bwp1lF9pfVBF7EQIv+4VMhuRQRhHCdV2aHMO
Qayvr0OWFnJfQZCz01wnGfyGBPUuUTLfVg13ZuoRO2ovU9vJnEzWYg+f64JqDNFo
jdT+3cFvAmwyUwYQo28pfKrlZ2RyDrTx63tV/sNcbpAadFz3RPYj+Z6yoMkK9oAP
nrGtMjOBfWxkkVNsn9Pjr8GYbaDY/dLczyccrP76OSoHx7LhX5Te8BSFRtS1crvS
Uy+13oHcHac3g8NyfA+illiy1dX+XOYR5GgqI9gryeVSFluKLRl1/hKCMWjfR992
jO6DHUFe8+SHagDoG8UFV22wmhOIyDN4lPo2fBwZT//dQl33IoQiYYCjmIzbpHNJ
IOhnLDsh1spyZo4QyLzUa02rtb0VTqU6CAgBhmQ/SoDWL0vDak8SyQ7sG8BflnhU
/ZblaPSlarnaQfOqzhWFllD5+xIUnU94D9u1OKPe/jK1PVANH1CAijrV32m5Ihw0
JxbGFTdKdUo5YBt5wp5UFeEhQGduxzvPrTjwZ2fzaN80+u5T7W8f6vyQWTCVNCUZ
dhBi7w3qSp8aU5xAg68H66r2dZuREJtKvATsFDeUYmYGuyu3E2kGE0vrbCzovB16
eVy0+0gCfHLVR096tnXuLufyp6z6WrxMDYWyHvwiYmWxMewl0HIQSXpe3mswSaHy
X8FWUf4Ih3cN0+y8ZA/oabEngaqjvFEDWRBcT9kEU9/tTgRoUn/nEm774kS6sXPF
wbt0bPFyeqS7OqOKHYR+XuyscYHp1WljhzXT0nOuJM7n0/WsR9Bd1N+x0y40cqeZ
2jYHo3170BtYlj/ltajzGvHz/Df5q0Skj7kUSc5sV5bR5XR92xlcoyvCq7ExesPk
0WptOetp8uy0WKtiRh8VmrPuYSH2XiX23hrnsEEI/mdaH+VhGYki0lYeZc65HjvR
CAVTaOrSABGXA0ZZ5sjUJ5o77sI/KoRn2tB51+NX5CE/aH+0xN82XXAKVULn0nsu
mUP07Wf1uDLI7m6xBEiyVZDG+mMu+M1AF3ZPNTROccGULMBbuGt+VVLACuiIzoNr
OcCmRGe1LMzfjO+5k6PY4PDM+Qp0fvnHbaTjOwjFA5w7m5ZQOF84RhAFnEc8E7By
f1v6AH3oy4ohXfZa2k2w+rEofqZBjrS/bu2rSg3Lgo0fqWpsFD197MqbCP7Ssq/j
tz9lBEbXBJ3H2CD+/pbKa2fdl0Bi92IzX7Xon6LOE5+tsR7xe6K4Uso6EpDTTI2v
NSTVUkM7MBSiEitn0W6L0wemnctO3LotQJGK1dKrtvp8zMGLHb2KT9SCXJUmmRtc
nE7jGhO2rEjTCg1heELxUWDEq9nhgw2DI/VO+bZf/KCQwpKYBWqGrxGoTaPWs2Tt
p1xV81jmHcjIejEPEWZaRw1hPTMtBP8rUtBuoMyaZpy4fKvD9Ah/PeExW6S2SRzj
+tpzWS6vgpIfuJjbG1JZaz2cwSnSkCJG5ejUv9Lk489kEg7HkNV+GBrigojBK0Io
GRMvK8xpThktioLYdkGiNXbb5px6d06494qgpk4wBkBlHaD7htZM40HAa/fGJSZ2
uwG7DtyguFLDmy27nJL3s3wL7UPGRKZzyqsWuQoBOJ5Y+FZn9DycIIqCODgv7cbN
QRusNvEuK5R1luN5msL8j10TGPJUQIAB7NStPeO0C3IR1nCFiJXDIhEB4VGJdx7I
FxePkf0jkdx8fdKQMriGHaGLYFvYinEYfwwi2E81zY+f7oPqApzNOpB48noD1g4g
TnqxD4bTEpZ0CXkFUhoSNbbMWw6uhAz1crmvDIcIF5HhtERPRSFL7gn1R61XHybz
8kq1qGuCZLDzqzF2qhsIRMiekQxEnHHUYMXq2Sl/WuKxLd9L69QGyrH+tKQdt2ff
f8iYtI/3L7bdj7WuIzuEFO6x17YPv6fBVYI2S6DSuWLYZvsUDX0rrqr8MSsMIr5V
J6GQqZJBTKLfNQnRzTIZ3ZiAtDulrCXQjHbkznv3olmH48FFChgv09OCSLTumZXy
6s8GS0EhObPMgA4nTG9WxEwXnICgsB0Na3PtkGi1vojCfrE1db7t5ybl37C1ZSg6
6dDingc9rmpSI9j6tlSfWQE9ayi9Dvo3o5onTlxwTdFvnDj8hseZhFJXlqDr6Oe1
lYmMFjS/8cEDkyS/Mta/aFAoQ/PyleiGVtJpDWRaxtkgoUM7RaR1GmbpLUS1RsMr
oh+40xe7MFSJokgYBuIhUUSWblP5bQRDUeskif2qvMZng7OOGCuy7MWZ5EMe2CEg
Ug5vg1seUYhyfp1z3juy9QYr8zJ0cnZNOenklwi3FKe1tzu4UNbnyqh8qZ4ERg6h
bKnAZWoECx3id6cTHR4cKdvkGVrGYJVINHF8Ao8q9gQM4b+3QChOCfXAvwneFW9w
n9PK46vyHrdBB+aOJ2iXB2j3e2zz9251RfRxYk1X69h9W60/UAXk+4kTU2CALy59
xpIuni0ztFV+wth2pmjGaz82IWkJaxv71NZVeBv8GTdMb8qNFcq1QWi+pFFKpU2t
6m6t/SMXqijs1wGfEFIGPYZ7UiEUAvejcAYISKrXeVL5k/NMT3ccl0n6Rg8UXSzR
dEmpGbw/f2igt9LKGL6OjDvW6qMR5tV2RUD6a3+KGu5Dl1uWq75efBJhHMzwUvKs
eSAVptISsuAD/YydkJRG5YQtMbgSSINbrn2vWvd26tWdy2QJAPQLBQVW4OSViB/o
yX+aB2r7Bd2qtQB/RmbEEWVYsF9NZOMGp/B1a4yOKOgArWQUDJNwlNLh1oB2lL2/
vimLcKBu1pjcOnPs1pzpak4ZL0QkOvKAEqSXBS0OW5gx5vOrSD6CHT8yUcLtD98w
yJyMTPcDxW3oYNV9gwYlOkeSTwbpYvTjJSy3OoEaZj2g2rfT20ChFJP/d8635nUd
y3pAe5++stTp/JIby5dACp1/VvnxrNLz/mH4ukvhm0WyHy73OAXbCLysFkWIV6tP
918oo2B00EQAd6OPV0jOMVsvS+w/+1s78B1my9pW4peZXEN1v2MII0AuMvMp7vfw
5pevpcPAyX6pISHA34k9vAyOSvpSCvRWDNJbH4jY4a4Jwj7O4UuiIH8bqkGWVGS4
giOw2Sm++E3vUnQ81iM4UX6vkV4CNZsik4Xt1p7M353FLLsljkk3uRlLlkQbeMZg
Smge3d63N2Yo4A8UG7db2lkukQ9pBdQs/0I2cvGK1+zBMQhjviWYq4ebpmQg0IuM
3SsZso7NP4J9IcJIi1re73n8Pp2LVBCEGvw7ULl4QbR0I/ZoXlmpaQOrITw9yzu6
ucF3rr2gClsq55oixE17opef1B7LVp/RMkaOtpdK40vFbigP3mZqKcpiLheJC03r
BeCBN3qjxffgZx3WzJUeGmPAlfgrRd20BU4JPbMsL3pCuaCQZboUExaMoSeu1FVC
uT4b5F8V/cQSES5danTdJ4gNsJIJ9xUukWbG8fgJKnavjAHDFREmVRDtff+gdFer
YHpT6Kb+GnyeUlAhj6YxAxAEpn5W2JnzY1l2jL2SnC7kkW8C8mx+5o5B+O3YGMcT
HXJYN2MM14d2gXHBWTjvY0xfkaVtwlTVwoezUnisCClv8AbozhawfnZef0gkYS8j
ZP/PY9OKkayCTKVE+2MX/z28BphL4KsHuoGkxL8PE5c3E4YylO7Y9STkLqY52KZE
Sze/eTS+gijyoOEVWt/p1098Clik7GQ+GRJ0NFkH2KOg5qVPuy1mHJZN5AFsR6BX
an5033ViKspP/X4vJt3FXZsxF7r2Outu0HT4Wx99PtjNQUCd6jkJIA8AhD+v3Tz/
rg9rDx8w/dJVlOekhLQ8yHL/N7HJeucVtcaLlMzntujFlxlDhZWr4wPowAsoXnks
de1R2LoIJfPgtAMFvXgeiMMW8Fb19JRmgvCtHCBhRpV+E1mvbRBnS5f3i9JbJmGt
M9JbwzvgZD/GTZNoT0HKoBQ8hERMG6YZYrLwwo+L/1iCIXUHDJTkD6OSyZJ2ZiBb
OclLcUP+C+TSy5JEq0OKWfkcodMG6+wGGdTvvB/iNFzn6d6QIbybYcQ4qFA4SNsk
2a3DTueRREuHyXNWFqTb301zmSU1GE07FwsynrqyH2VABy3F6vwzLy2WpDr9j/ZY
zLT1724tcdO1uwlFB+knqT/sS/EgIdZvxWGBcAxX7LHAQJiGsirW4jo5Rpkxy+oh
i3nKsfCJymNPosczcKjTQXtcFs9+jJ5+afU1F6q6lTej7cA4R3iQZrWML+4VEsbV
iSlQAmoJi5yc41JpmtdQi87i8/N127kk9LaKdSOB3p8fQaaGTCuiriqR0Q8hCF7Z
My+hvC57ufItfNnOeuE/T7aKaWfWfO8DFh28WNbP3en8q9HXrvu+4rGt1sVInzeu
ZgG67FcuL2AxijUTPyaIDohx74MBkucHBXLuoX9P3VEtlwkBxfcQuyyFHfEvpHCD
iYRUGJCq6O48fRQGI5qw/7F3qvtWO7Ij/hZ0keuQyMkZudjX26/NveFm8OlSFzX/
Qj9Qe5q0vZzBDHPDU91sVTCh3NaMtJWNyu28dD+GGXNujEZ0a4z6Ag81BSGT4IFX
EtriLLWgeCUnha/IRCTRB7IRwtWcPwFnsmyLQpUGZhQXxI0tGR24OuOkPdxfVKk4
V2zC/a8us5IelESUv18XDQiB7CjHHzA2NsLKIET4QEZp0/uP3G8kw1q6IMLTfvhL
OYoxWcvF4xnQchQkacaVLg+Hhjv+mjyrfOxePUczgRflkJvkkPiyHI9NqL48e3jC
QlxQcRIC13bdAQE4AsawZB4zUfrVYxop8ShhTiwtOe4OfbfLJghEnRqS3o2GGzs8
OyDjfeeYj2sthmnlF0qodRj/L4Pfy4w3hsliWS9T3pOuFvacEGiyIEicIrfBgI00
Aj0HoL2LXxYKcW+70vHZxr/chvq/yCf8LwA4tu3jt78ruFnhodeIlAhtGd5QPvBU
Ckv2zJHObz4Vua9esVDoPvjFHRyPu331Ru1vgUdJeq9G4xvQ3woz1gqcTDgTa6MV
DZAv/wPucRNFtH/sg8wZLX7ZoHXdmvTmT+B7gta3rGKRz9Z+0JeWfxIGB4wb/S/v
3+358uIDNmh4NJifoAxmgd88/OwOS932MyZ0b59tZPyVav1GPx3gOqBOXPsggU9p
VDAOQz2hKChbUUmegIA/mJK3l3P1tVM4zowVVeq/eqYCKRGyAdWLDASfYM5GB9F9
L/CQ88SNe5iNK48DypnITpnegi1G8d3oz06RuPiZKgCjIGWwm2QnANHIsNb4XvDq
GoRAGhfy63J+ecLlQBhPcjCWEaFrQAoIM8LkKIKPmaoqDpqXVts0vmmdGduISasn
5uz2lgciWetvgQW44RXGLU90c26b5wBv3ZRWIQ/Nc2Xd7JiSKbdxZMkWK3RZE00g
iAcx9MLwtVcij098IMLjI1E6oOeIY0aYlwS2EdRisyJ+hsYQGutDv9UXAGKxg1zT
A98L1angUR+NmNfBWq5etiTr5fkDXmUvaseGvPPCXQLjCHM8nC+/m0uG17pt4WIY
3IPQFUH4dBSOpd47WyWZzXWFgHyKKJ9xQtiJkBJGV3NLx9AUHusI4OibP+oNCqDn
cF8+wkBI6YvIrnQXNOJZ4dQdp8fGtfmMDs/4bHikijFUk4poi+GHBTz5Pakc5iRs
TcXlrSkNpxLNvmM/xWXuZOloYR70KiFbV7fLEspyNCCZxtMH5SYeWjPcUBxgT4CX
GDbbbcNtxKE/1jOCKPHDGpl6L3HE4tyexJVyBFJ6UvZg0CJLS7bABOxsBc5sgGTf
+cN3MRC2CG/zmv+0sQ4+0ju3CEvOR8GKLIu3LxZI2JitDTLgNs8ZGkRb0i/QRkUU
lVxccKoktgpw0m2+eUIiQgT8JE+v/QTYwlcOVGPbq7mSmA/LEKUaYtvzU4xikeuw
FKNP1OMzE+13zivTCnN3UP8g+ZkMu7K96yO7f4PAv9hAxJf3ZJDsxKEc8u0YPop/
iODUVL3iNRSpBrMHdy4l4asD4JuyjGTe8/ApJJSALFODgCdbX8w0GzhZIOMeYgPq
FaHuCbCETmii46ZqL1RMHGNoQKWXxZdFNQvOWnzqqpCVSNMOXYJZYOGA+ZCWZl41
RI4XpYxBfUhhpXdNibLoKmruNjxkL756y3gqU9065V1oiUT48Kw8ttUTQ+hJJ60Y
czGTxj8zbp7/f2gSEAvOnY6B4bUAOs2MiLzGuM8rS8z2ke7Ms3VVkYjYOGANhyuX
pjgtu6ccHkzSr5sFGkxvt4DaVrhxh70EawKuWFDeND82tE3npRguOXIzQt0vWKuf
wP21y1lNvDzBU8si9yGeN8o0EFBh2jDyVgZ0a3vWKZ0EFe8uTGmVQ9ddcQbemca0
ftwQ4NC81gaP+rqnz7s4HvIkeRbB187MTXzZXgTpK1FGIcd/MjThMlN6nO/Hg754
KHzIRozctED/Y17rly/yh38zl9M52NcjmVhRq0NjcBJak2TImexZCd61vSiQwDi4
OMhsgzwcGiLpHp12lOvRk3Zys6WHBJ3d08HGppZ2vie3AMo0/VAIwsY8zD1VQq3a
E7f8LnvuLsKwkEfrG/vIUDRQIKWr0EmNiq7pYa9K0OWS+TOwNryJm3t/+A2pN/l/
T5Wj18k3IA/4VLpU46g3GNMM97HS7hfhkpQcZD2fTI5FRcQBqCpDbv6KOGkcgqbG
yrQO7PdPm29G7WkRm57tVzrX1kHgsctF/bNZXqTmon958JFzNORgVZDVxt/dfLQb
CnZ3XXWN9lKGEW0ZFsp6cnLYn9o9eGuQ24HW6h406mAu+mlp/P+2BT6XQJ6PmMia
z4/kMn7N/r1ysOWliGedTCNm6TXy7JfOHTlwNuEnRk3reTuLc6BBU6mPRiuLH6Rv
80dYYC46obNDkbNtkg7gSOGIRPRBb7jdGtMcE2eUW7WqD1kJSUMc6diXoPMHcRDP
mUisAkBjXGxu3HavNPaj0d6I+QV+6UzCkObXyNMto/BlwenMZy6jVmPNG02AOtvO
YbIBTGxWQauE28jOsCNFJa+E2NMeTEPBPvJCwSbP9lSbOD+hCI0salYxFazUJqur
jvSej8uyoW4C1OFpM8sxbI/7clNyHajhHTr5ymc/OHXKdQnPR971nM2yWwkec5jN
2ZY0h1yOR8mT5VVacndJ4otJnvyNzMo2QL1GAMkXbDSYLHLrPM2O1cOLFLwOAcW6
WDUH1GLFGJ+4ViIx4Kb9m4GQQ5rqQS/RIrxFvVr0W3i+Rv7c1cmmRPcNIZVpdsyl
jhD2NUELJVrfjNt+Q+xeQaytxaVw8zAAwUN5sG9ytIpml+toU/KUU44hqv3/MjlF
sMK32NoBpQ4VwGeOQYl1jooL7GsAftlx1ytnvZ13BmZJ6eF7avm5dUR7x6uQmk0L
vgZ8TuhvMVLx0/GeyjiM92VBEI+glnRzXMCccwCh1la92F5sKY7N+jJL3oE6IXbh
2TY0XdpvApSg8jbRgY92bxWCMpt0KQFM+ga2MsOwJNzsCnkcBbXILrD0bZ/qsxxa
BKtbtrPpjQ5fgbqW2Mf12QIXqoIQdywVjQX1VBHKjKEknzz8Qj1D0C2/qIOOb9q1
eUNVtC2gIPFY7g6rS2zR1E5eqZ42I351cXOwdoC+YVcJ9B/tZTuvRRvX9+Bvfia9
FJnua4AOj8F0VrEgSKIL98lto/mdT/yWaHtvnoIDOX/uHiqr5fSdMtZEacq8bDiL
2f8K6l4S6FGxlBBAiLz9SN3BBg3eRNhaOgD/g657k7Lo10FpOSopYUAQhPKcneWv
7DaS1pDyKxBUBOu/m+C1b2GHWbjr6QMIVvRBvwVZB/ipB0rJ6UW8yxVVU2CgZh5d
NrYZqNgH9kPtY7xk7/JL/XPpLkhJTFONvm2KOnVJmtkkEexnPRBep3jrhqw+9YGo
PApZPI4ySlK54CDWm3737aFrAlGI8VXvcJLAp4cOdEwKIAVcUgCMDyAYbOnOOq6U
vm4AudBE8hGmeHL3RQYrpn8O3fgbFbLuV3XEwwVQTIg0oCJHP3V/atOuyB24/JNt
NF8YLmWA6nKryea/xZYV+oxvtxWQQFIfIKqSLjZnMQjiKqHQZl6pe0nJkOEyqce4
wNvrEQt8RcimEsDoYXDdOL1BAGWHrsKS/4n4dzNy7Qefox2KFAjjKAzZ8v0GMTXC
fPJ8zBg9Yqml9W/gUx3wHIzdAhNBMNY1cY5xXs16aQm8hCuMl1iahfaDBRJE5lwr
kB1t8o3IfrHM+2jEhOeidbVKF8DtmYo9itnaV/bZGHRMXErg6RXkM0ineW1173TC
SwumU958DAMHiyEDhIpLeupZu8ou9OoRuTgd6NIkxpt0zTip1r4aXp+JKnjaLTHV
MhMIJ3941xoqRRvjhWsyNk4BI2xosWiDhZ8NrUR1LHrAhj/KGBjm8pwS20AAycwD
U9+WUru6/LgbVIKqmHcpMyfWSK86QhegJtheZYyusMb+h398W7iVsQl+FqmR+MmV
Wxotx3na58w6vXk0XwY2EHLrBAiKZV/2btxHGtOH944bH7vbJZSodTt8a80/6rY5
jiXInQEv9KClZTN95QNrbcHKQYHHwtJxWcPIEPO8LjzdV4bRkrlQ2oxd7qheGRg4
/5zVF/l+i8V6VSiEAkwcdMu7Vkun1ewcxAOKZIk13Xf7qNVlhBs54oiCtqV4XueU
mzPq765mbk/lsFTkN+9r51I8Cm2oXe3QofeblssgIJ6TQ5jdk9gIHYY21bOV1ZeZ
OZsxaM1evNDavX+5iOoHN3AnMvMZTH5GH4ynjvOSLscidb2HL6bHVd4ckorGoA/f
ifjGV1jl9go1udLQDgWEcbFVODcYpnAUxg6QpMMGdR1ZcI8Mw1kXDF+ScTc63bx4
+mi3mPfc4c8ugzZBDij03mXaXV6XRNH2a9auQJZSdYdfegwFJfGTDIGOstp0KPjL
dCnfuYY8paPywJ/nSQ1Wz2Uz/nDXJH6TKHSmk6ZVFZKATTxQVPdqMMsuYSbgt7nk
xsGZkvxTbLD0qHD50w1MYVRAGRnkhwuCjHAO7tqNwAA4XM6MIvho9SKC3Qakuuiz
tqi3jSAOLeV2EljrJ5LCM7tkTQW1y7VB8SS5Gwo3ZXc7C/67+qpxjr1a+Tsw2d9I
09PdxfD17OFXVVrokGCpGu9hbt/qDApm5ku4eAD+NSts1ZYu7Vo6np4oFklqHlJJ
XBIXxBmrv/OO93+SUSW/SuuPmkRLa7fYiHUfNiOwPDoHED2CLJUbxePs7XqNf/Tz
gc5vzKYAD1MN33BVe9HebCwVoAPO0Edsf3tsCJK3INOjxmHvEP//oNKEnxfTx+ps
WsoBHfjS1NgJPhqvNCUXcmAoopyo/Vzo1c1nXnQ+Eud3TFrnEpdqXjHfFO+jZQSA
Jp5OUVXyAbIAUaQmIWmpN4QC+tvu0fHJ52QZh0FgShliymVCAGLneAUPadnuHzzH
b6T3HDrjSbE/zYLLFhZ8aXUkUOvMnlO5s0LUDdcrFCZZjoQtbTHdppAptD4P1thu
lj0WDZun90EOjABcyTH5mEjze00fq9IgWjrYlAUvNJiIp2e/MwyY5T44aCmt+9sa
/fceKV19oxnIKgtyKnHzStnge1lLCS28LEgmtPxiN/emRu2XQcIvdkpHu4i1XeeS
czYglOmMz4CCQYmdlK6nSVXAiaTFLKxxnwwhzTDXpRTUvsntHiwPCZjNW5s7TD9w
7YC8t6r8ovAxctn+lh9xU8inLU/+jwBKQUQ1yaWeKhmwRRI8qcANL3kkw8XFY77L
2zizB0IYkhsIegKLAAFOsHsBScZNUCRPx5FeyiJeVCIlwXgrksdW32iRBxRsdToY
izrgKvyVSe/Ffr3LVfAZmfhsQ5aZNlBEh5tFgF0RdlZzlIVmvyGUYl2sWjKhm5A2
RsMkUojUhcfpWSWJC2HB9eluGidlGxl2+UPS3f91ZvpQst4jOwpwM7cLp2rICUgi
iYbPbpE60VqHulTdGRQtw4BP6eAZYfkVtIVlcmxCHd9nZZY5fexLLO+BzH+QXVME
lfEAv/ZX1GzgHCdYxVc0VYhI4WqpKAUMbTS7ZBZASOEfnStLTz3J7LF/5FtXj6k9
tN3wKKbuOhufTizzlYKYJQdkTXz2DayErJ8wdc7h+DVIAF2dmq9icSxTSGtzd8eZ
RJtQkCdg2RlWhcGQsx+C9IZ2UlKFraiuTVEEtb3v6PINQy5GVCMYQCuguGLFS4Z3
JTV8dUypWqX7E8BTsnOXz7E+EywEyWYL5Sk/sBDk4JnC5dWAsfIoXuCf4ceOwV7h
ohmwvKU0/IC/OAw41KKzpYw4+wVtaqxOVzdc3XCL2PZQu9KV7l0VWI7mEiwjx8Y7
rc4yGWGRrfmHE8yZidO1H98j/Zf+U9IMyla12OcqIWOwwP+B43tyJKDONL/MRpBV
DZQt79gcX4HWONIq3xt/TFUxT5PdAUQwenKVymktIw83XOhAgjZLLeJWCO7g1gPo
9RMMXJy2qjnlGd9u4mnD4h1hMm7hmLWE5E9wHg3+muwIxhUJYJLckABfatrELD2T
m0V5LrygphhIlHzuyNrXJcmIfmbOsme6eILbiF0GImnj0k7Bzeq23f/PyxZDBOPY
QebhjlUSIroZ7qln4gvSxtdReF28mK2N/ZMnolWM8IPFSqP++wPxDMda8l/ZUuQI
Q8KuZS1aUMikohZvIWoN0FmP3btZvUJQf2hPPt3OShzmGTSGoCjrJXbIfkWc71d1
lNkLBYHPZWW+1w6y2Aeu8vtQoTFhdVdWW7r4m30IUohOPfGczeZrvjwPLnUrsuL+
RrpX0NJ5wo5+LjphNbZZ0slp5xucx7RHl8oKyRJ0ivXo8XmHJFaoCIkglfKaWBIj
0iEpU02UI2CBpyhO4Yydn2CFW74Pke0tZCy6Y35dZrohxPuQeMLcbtSh9sl+Zaii
WcK4hf+V5qbZE8hQ/5E7PEmYah8UEKf0kG3X8QzsFWY+pr6RNAjcwQa4osazPv1V
zLI+WWtlKVYgIjBZu6dHLIb1RIqw77NNj2esK+O/eRW6kgEYOKDpdkaMk6D9/btK
OLQ6lkVHD5IJtHpn2LNAW9k8oIzH6uZcDuXgpWUOG/wpaRZtzxOVVQs+v2452djE
3V6pHg6KSzLWZ0dtD4ugi9AqgJT+GFDqeYkpojdB34mipv6QyujIhxglHDbwzVmI
5FPe1n/faTfXqy7SNLG4YJjUp23AfNhLi6EkOzaPr7fn45+yGe7WC24CJK97Gmhj
W6/wOTD/LjG2bVRchI4FvtHri6jZ7agHSePRduOKAGzsmPQqBCCAR9hxm6Bo3r17
WdeDcP7PjSqE1x/kmwdAzSO4vWzJn3WZBU/sMxWr3GnczhgLnnhRKcpZYtoOd0Xq
b+6kvSS91A2kYWD6/eJ/T0CxLJcjTFrLTo9w0VndxtmTbB6R7H+dpEKgg4rrCwQq
VngHU43GXNHntOB+pFr35BRoAExXJu/Ira08eQzFlE4xL+v5QUKBHqNo/3esajGb
J4E1VVe1F/gUFaW6BtVtk5BSA3pHj5L9iwJ/b+xpdBAvI8HI+h6Cv3l6vSuZavt7
9aBE+PhwJud821afjdNjuH9ybtF+klH8dr+JyJo2f+bLG995K1CH99t9cWT4STnb
tJCmlB1rBe51Dp4aBV5/YWdg3lhde4oS3WOT/wAwnCw+tS6l6Og5m2gqOi6zfDqo
Yc1HvQqhf0TbiH6k/ld+BPSFNB6bz59S+zQMYvQFhdQQCw4pH15zH/bJKACES8+q
7yXT/ZjKcTwlgvswNbz9i6yYMs6+X9ZT0IWNdx99/Xhfj6wx3dG4OoZ9KvsusjhG
wZc9oknwshUp2Qmd9X6bY1T6HxXk/wIEpRYCxvgudCJr+Ok/KrdiAJHjoB/igDc8
zJ+CxibZmWlE6eSYUoVFJyjhWKt2VEjxGCiG9m0xKnYCuNabJ/jwz07xbS7zdXEU
ogQWTJZeQYoI30LzfzHaV/9LIdn6AD63a/khxGWcaHZOoE4EjmmcUoorKh5L8ZCQ
qMVmiI9FUhT9RfTkDvKkIrFCRjS2JMpB0T3zsjd61JBtcw5G48V5qxPAHGWX5BlZ
UIV8FnagkYIQaaoRdNlpV+YWQTEqPM6ombjfaXxJ8y/Fi6d3fGNMF9sdDT6Dca5p
bokTbPw473K5Rxso8izzvm7NQuKvx9sOzpLnLVdwswfxuQDa7o/rgMLQZAkvpGPO
Lo00iWMYPA1KRsWLEDuat+JWskdGX92Vl5z6w/tOdYox5AZuFrj0NHoQqg+UFZl7
yWu9dO+Kttmg6kUM2RhtEJuXA7prUD4wkSyPcB6nUMvZGtSUmH2HwnD/XeoR0v4a
7dtvyPglx14UKfLDyXCR0BbyqnqX1X5ydea456614ZZJUN8iqOGw8C3zhHOOBkan
jHYDUEGkjt3fRP5bPNWHW5iZ15+meUyQIKmlwaZFQcF3M2auA4DM2ufFSeDcgvYe
qd7WD34dLa1fUEuAFXblH/W2YXqI4N/NWqewOOcfNF8rpYq0V2gb3H86HwxGCTvV
RuptC8s1A8+uTaMVMPnjHkVt6V1XpApTsnozdnhTDbd8zYku2e3ZksNNt9qwzeeB
elqZxgTqFH+NeL5FKkHsRVoNqqDkaWiLnjYgsamYJBImbdelkrpJlSzIMOh9ZNQr
eqDsGA9CKpaD0sGQazr9xttFIMd1gRxBb/vX+FTatSzFQN3vkS3VS40KrJ/urHrE
uDNR89hXvhmN7TcpoYetIRpCigNr0r6j22Pb3ZbcvOMX2++hPF0i8c0CcO3+R5vD
Qiss7IZm2AfMNJBIW3Tiz8R0Hf7xCVusH44M+ZUcCF8JsSYnnuAV2E6B7D5NVx1x
HaUkHvhsJzE2FtkwNZBCb5lrclS74soU+n/7L2nSWI3MLnegioHf2gGbjHj2kLep
vfiQSFeIK25mr75S8u8gBHoUtQ0UE92zLYRG7+3jee+RRZqYR5O6FjYf0lt2vEUG
zwjZACiA2jxLXtal4lETQx48FKCCsyV6i2PI2ppSEUXKrBTWvRCMYjQWZZLOzpuh
hYsu6T3LLH+SPdANpvFp7ZmuK602jOOPF+cAuM1t628qltkP9QMDeHHJvvif9pdW
Nkd3auhY2BqFIRE7rpwCoWBkrhmno2Msh98qpfmQTsmKfowS7CFe8yQw+KBXy1QM
gnXbEIEKJBfDMSuizj1B2pMzD7VC97YRdQU7xviZfmJb5Yful1eAwzC1rNKP2oeH
n0g5jowA09d/7pzVkK5WXu5WOXYPiMqcmTuxlREokA2fRDlz0YetIBxr9rM0LrP9
ey9GnFQojmITOxBKa5h6drl8qP7vCCtLOS2uxHP1hb6XAF+mOmymXRKg3lPudZO6
8HMPK6oTKUaNvvWzoi0Z0NzeaK94scej4aNdg+8rJehAEEbB13RADD0/vyE+bkaQ
/qqPykus2xRdv7HOCbAXFpAQrEaU0FNz+MTCGYYjaFsmOiu/3ZkcfdmSSIY4cxxA
Cu+jchZmYlgvbfiKlDEQeuBK1prLW/NuCpxY+EiIfDxKBqZdSZFhJfto31Yg/Qs2
1//+/v6googK5H3LV08z0j0xUdpXDxUQ3/ceP8oYnouiET0Qz0OU+kZz3rNMhca0
3HShaI9kXdHMaVYo7UILHRWTEG8yfTSNfHHdQ75vSLrPw3aBT7t9b6kMcGAosDwO
hAWL39k2dNSaEkSn3nWoOCzr8aWlJLu5GLyRiVmnOU+mJsg/k8z6o2lwOC6Md69c
hDH1IFESf9ZlF8Wtp/V59KJAbzU4Hk+dLAxH8wdsXuK0kDHSI7FYA1FI2AujmyMU
/Tkb0GhfR00NvRAFVBiBcRcp+d9oVs4N8EawGnnludH4ZwBKth3mXp6Vz3G3IxhM
OvCbBGdQsxL900+LjpbGq+LWjEiswtXHeFQK1fwPNcH1ko/HxdYLozFMwIdYcKBy
Y1IeLxrBo+bjtxWw1JZD30tzZjZTUiBAzlsYVwE2AICSiwJJCpJWxKPdmLURgKre
aTD0dH1xTVaT7v2/UjYQaIQlVYJ/5EjgnU+b+j7i7Fpf6c2s18rUJYgn/EN9HDjI
L+ni2sUuC8VVN2emT5w2P8790kYTgENeDGN0auo/NyXT7x9PyXxG1UaA3GCN7sTx
NwL5nVr+Z/o95yJMM5obQ2Qi73bL3gn6QvlOQAU8Uhka2bvuF5INqEg/4sNTKBon
8EMSUbVMXxIaEB4JwKCCLYVDk+/LGtRS3zKyywLtC2K4UwvYjUzIN1ZeWNSoW3jQ
HUUoRyep4sLztFRiZAGq055iX5QmgBuI4slPHIlszC3/kVDxY6/eY/iltaO1RkDN
9E5jw2sCxXqpcAE5P0kAXZAcOSJR/IWVg51mqNNvRzc3MJ0drUYAP+lQm3UPSKNj
+rnpoCl+n5K86wqzoDj0gmWNowrgzoz5cIDe5IHg0hbfrf4CNM2XO+Ii+k7RhuLM
tKfWu6pBgij3F+x1yZCF9naPB3uCVM6730kCEGbeS0oW8jMMeVc8ap//8r23klmi
i/Yxvs1QcocoAtrjoXf1kHZVHi6P1zTQ4a1A7ovYB9i5vq0+xZB/bYQdK93dK8Mp
LaSDkQGC/K4h9kNn13w4xK8D5nzXOPEuiTj1T8eeh0/o5aeIiMNI4GNbmyXO+SS/
9FpGaVeCBcZJxAYSnhyI4WqLcKW7T3iFqoydAIGp7ku6lwAGsff8cnl1GzGLJZg9
Imzc20bS0DBXPw96JRGjheIaXc8omzKuc31TWLlsA+g3ONvN0zv2Wl8Gz7Dlyqtd
jp8L6TnMVXpp0bl3ctms3aukeHnwIIYk8u5BrN2GeO/GTV4siai+SjAO8L8ONcKf
IR5JFwaLnQa/vDpAY/2bdx18+7ZFKF+L62yryvdPqwPwwAZvXDWCqE54WjTN9LdF
BiDz+Uo3cvaOFtzrwgZTA/ET0q//NZ7eaXpylBWDzc1jYNG/I5p39B/cOsdhlWAU
kqU5DEVOWM2LNWzPxEtjudP44YzjzcOg1nxGvWex0td2pT1D+cLgwceqW6VdsAbB
W7YvT1xkUtYyW2uRu01N19FVfHmfb/SO6Dk1GkM/mujnzwzR/+66SUXYmPcYO4tK
5nvAwvbtpJOOmrMRqtTLyirzKN0HltYJHUZpO55LZ+3/jubr2/AdsD31rtyaYozg
ch0LbQHEM/jFg8xtDfiN17tGNR8WzQJh3E5jhZnhrLv8AwQrANz1FiNeoocrvzzC
O+JiaUZ4ChPVhovI8LQ3YBEWyVhyk/+F6rM+NYLyJFWyV+vu+UWmhaMqV1y8VsH4
969oiOyiVYCMKLuJ+pTTLWodUq3VXY+QB3FKF8Pl29f4JBg0XbfWl1YgiOPibiTy
GqnbCqqlf04MskYm1/mCaVELCx+esZXl6fE8p3WTI3zI0ev2nnhnuRmqQInhPhkK
Q08yWQiDgrFpkRCGQaD5VfHa/6kn32fkJYkr519YC+NgEDTxhitWWGwN/yiuEzQt
v4aKzFHu6YJLDs14WBhfQ29HByv4+qU0RafvTAWYsLbkoX8a9+Np4fCnNGjNYtyb
xcPcniR3TVBwiTDZxqr/j2i+UslH+I9hbJMHMCiSczmw0Y9O1fRhChEbxZvOzhuq
FbmXnX306OLVjYQYKelphASKr69kTeb3ZkC7d/hkbJtDMfHRBHnmVR/YX6xdsWqN
40xzuAjd6d7ksWRr1Sjkg6R/NYf4QMfHYYmvgFRynA1UT4AG3bQdksx8DWDd8kGD
43HmYiAWycJRt8wQy5exhd4hdJoxhz/Mr/m9BrtpDN/uJj6HLORT7pjOPCr4xurY
4x5DRSk+4/s0hs6VGp9ciMgXhyU/7Xmkr6KQFmxSeKK+xDyHqvxFD4nnNyLoQCct
EERjGt+KIZKu+DWMvzz4YGmFLzIWnD/g1UNm8kI1yHxKozhNe7CymG1coGY4NwAP
ptGnaoJVxEGv6VfBwDRAN6zuAX+P2WnCExMKuy17Nl5UPOAttMW/atUbJUUXiN4G
UEabHDNfeOr/ZgS/ufBocgEgRA2XcgpyuONqLix5cNB4AnGmQhgLZADiNj7OI4R2
k4FeiVfFCGbKXN6lq5Fu+2/LGAFXpdjOVXLDlvGn16na1PAoeSgBw7mwBg7LG306
i3asVu0jQDjvZDya1oKu4tdo2cvuhrcsi6EgTp3/BGonpH6wlYcz5zs1SOVOfSNL
VGVh+kaDjlL2hoZw5SRarpgh7DU7xJ9ldUtbNo/zx5sMz0uBv1u6B6k70ENE5/yL
SdtkRfKmFZ8LhzJRxt95lakSFeK9e39RYSAEgG0lnEj05sFffto/i8mBzS/W9g7k
p0xwSKVa3sEr4ogo2NPZKGVOMgliNWAR9C/08jH56DpJinN8v0+XV/0RIxzWKS0S
kLQ+AvMwC03sxM+8WZ2JsPwP0ArK+d/RMDPP9Ma/h53AMf3CJ30xuPjG1BiG+LlA
Y4mWEes6oWwnYptKVBjg5hcUVpUEbvVlHqjZjxiXYJzOUOSkFWPhHlPprXY8xlC4
A+4djJKsWxQbA3tXTX9UhHH9bgKFhTkiKxBZQJB7G1IbwNbSiegl7TQbdcC/Ha9J
NyuXOIc2WJBHuVdtISdoD1FukHv4+4XpaxD0hcMoX8DLzhe2wwe7rOhLv4GnEXTF
dnRxEhnV5dS6MLu6blDnPEeN4JcZhsY6KNT1hMrlTvnzKoTaDqTW2hPbANbVSDxZ
lfbYUoCruW9nG/9cBja2oes5d4AXNxDxEacDM0XPZGXRmnQvmAI6uZEOvMHi+zyB
Q2IqaXOUd5dH6/W7XHuzDRU985yQYjcqyqXW9cL6jUBKkvzxUUVo3x/OUmOxdraa
SBkGirMuopH1PFEZIY6T2lG16w+9TDCU8kReis0CdIVw7+JOuhLIRSWRmGluKtcG
Xf2Ff0i6YZY9aJg1U4PbthUFES55HE8Oma6O1lGQYyzi+TEgXGBW5xYPBLER4WVz
ofrgIlkfvvrRM5DMVmuS+LGCYDaQAL6+D4AbSY9cdk8x80tMck/nwd6fO8pDE0aT
qFnZr/UMqlGqM425ueqonMEZtEaXQPeCgcacXE3qilYYEjvb7kLDtT+HyuP3GQ5n
8KYxddhotWayxJG4xVfyARGTFftnceqEMTflWdd3HddtPY9Wc/BN3jQH6rF23kAY
E08rE2XTxouPf6RmN04ocoiETVgdnEjcO73LNsCOtgQild6WKkPzofvxrLZzyfIO
3v9V++dlrJx4FWiR9wPDNVeYvP5skHBHepCxqkvUB0UlR6sXmoryLOppSpmjdhtj
BpPCC97QaGyrP1UHA+elLowZmeLW6hhACmBf+bRdYrRbre8/kIXD/t6CmsL61ykW
/iYBWK6lGl5uGywaxBeCIgYWAvpR7UhlMjboN4jFNvxUFNtLn7Vcs7Bj4e3FwDdt
SPX+4xLrpGcnSlJwfFaU3nOgIvacCduFD53iMjmXdMauFfBW+1nFQL5cl5B6GwIc
MomgPu9G9efJlfTjS2lLonTOKbSudQDouZcjMeEjg2O2rPqS9xbpQkbYgQQT97Rg
7s9yzybyBIpPw1DbUw/TaDpxKXb1KO2DO2HNjf3B47lcraEycXdWdgWx9Fv++kfc
cMTQMmMcNoVrQ4b+Ub3F/xjLQqySts7ICCWZavf77tax3vOSmC8O4reFWoN4lSck
DX4z7JLzWjwFLepOXM8mqCWe3lKMEYnmMxSv9/CUAse6/J3PmsiNDrSROLWPauZz
Ctd0/rA89/w+Ax8TXSpjsT8dOEF9XPBmpj+NPjANbdmVUzRV9/aN6bMIDTnRfHOA
GpnnrCcwlFBjwGdhOGrz+faeTVqG1mR9zfdZLeczY20u+g15qSOV7yt4p3y/B4EI
MoG4DbuixdV7uQpDyW+pjK7RtzyU+IlUNu27I2CqGtkpK1V83jk6QPpebcQYCJT6
N7UVfYL5J8yUphaiDkBDsOPquS8sCNnFC9onD0oj2B3RL3uJMY37YFs/Afrt1BiS
mxKJebJvobIy+jUrBVXOXsCChHeuo2pM45tmnQnlKKCTgLrw1BMT6iFcQGSKgxeJ
kGXst9I22wAaLyTc1l/BnDEL5uSpmVwylrl7AYQvIPhvvy/8VZSZYuoleWghsTlR
ZhxSeWBxStLOjkxhjU8qGIe1z7bKO9nibPZ9gzK7qky+Bc9flB9C+EOn2JNH9orj
JB8PiqRIWLvsGR5ufdDc0BmnXa/L2izHaMLpmVS0DUmfXdW4ak3qNks+RMgd0Cma
+AQ97pQg2XByd1g8KjpfJxsEsvzXbbtmjFQiqx71Omiw7XIMhwNCXGK/Ry1t0gVR
9F918vQ/S2yd9IpJZq8eMSc2OOBOVLeGU4N9Xk/ErWihUBV5Weu9xwZcAnRUl+wT
to89MpZPsMO08nHjXZT93Vhb+bsOX34fTb3P/rz83r96GMaT+HOaIZlV2+QnFwoV
3bEAXUTY+seCIlNkTqD4LVsOgqSmW8JqflUV6il8bAlqo7W+rWW1jVJtPWrtlr0n
r6GBE6CKGE/63iniCyOwibkRg4V8cI2UjrV9hN7KJqw9xz41LDHPgfGznrB1/mLG
iohQpNaGjwdhskFfrkveaMuytZ0UJzl9dUb6dfCaeFXdq1sdnJaZp2eGAemXgoso
Hi8ockwR49GmBFADa0FFa4T6eFgB9VfAKzqDw0MzHXZxA3gSoHtyB3yLHVC9/K2j
2sZ3QH9jbL0GtE8KyZBfMYWn3CkQSFitcv3CLSGDShSHN0Y8Po1ww62yp512grXs
3HhGRER3w74i3WXy8IkrZgl5l7WyFOk3yWgK0+itHd+OTj1b3ATlBJZR8+JXZzlC
FQ5+U/zFAM8kzn+YGY8kJ4yBmN0UcIOySqlkHCydvW8zsxKe7cz6dXqYzWDulKyu
yKprMswK7mlgWJNkPsO4C75Ji4jUwMEtO9IiXfb7PLRkgHeZJoVmpZEDX7sb2NmL
L1JSov4ZatD08t1TdutU/ZINLRTUvE+dgRC29FznX89uoet7KAVwKeDtDdHaPgqJ
Hev8p8LT/9DsBWuB2tmjIDL37jCodAk3u8BiIGh3Msqszf4B8oLryRfgH8saGZ39
L+jQJyVw7QD6L9CP/FTsyGlQtnsfJFR1dc+zpshZvqISD7T/fhLVOMX74YVRnz9Z
zmJunPt4KRWXNmC45r7KM2MGWnXbGNDK0ib9Q4lUPkAV12zd8SXqufo7GDF/DkR9
z7hsNK4a8ux3U3CA32UquclgORvG+frZa34dGCw+BKPGI5Ilu3rsxDvA3vCoEkuW
OIMaj5DA0DFaPO+DoDmp6pKAVAkT1pdeNVe1L/Q/PURKic6dSn2+EpGAHUzY3ifj
c1AG/ToUDM0Bffrmk8tIVUmwA/MavGGi7KQxjDMiNj0WjO7m7mz2py8v363Ywetw
BN2QS5f6Lo/32POrwIMp2IBnvT90vE9MW9G5OYtyDpBtjpySug+oHPl6m/L4UFV+
+/F+EE6Ka/D0pbOuorKjV8CocUsKlkGeCntoFk0GrPfoHnxlKcrie88Tcx3PIu9U
XY21aOBg5S4486RaMZsY9NbzXSxIVv0cqA5IFaeILYZG0C4++DIW5KcXeFs3AKVW
VrbKMYVNy2O4IdAfLKatPFashxSaqUf6O1tb+HnoHbuzFxvKyyqutEZnwPJC37LA
MLmWmA+RAz/YvwTXULKku+W8L3U5UnlHUm185FFL/t3OEatD00f/hmDADK8SpEcE
AB/hSO1gdnRjl1fF/4lstZstlmJHROjvjm8pPoohPNuGurTMB+0zOPtZRJtKzOO1
4uzDVBPOKtkaD4sICC53KNiJaUwZ9HHEDNPLZ0vWsJoFFz4x8W2T21fHvf1h+enl
Tq6lUR4EoNzaIWZeJfJuZ1XesLyaxwm7IP9me62zzBv8u49EasUMz5fiVWSiFho/
oKJ2RwfVHQjb6sWWzHgLVez3bjkBxnA/z8SI1/AAtDFphR6t4VGIyhqLsdwJwrHr
7Q4lXfbvlhNArJqX6RMwsA1xC+QEfdkPIM5YSFgfQgglfUW+GFfy/yY/u7kO2JSz
u2ewEuUxB+2HikL7rhvFy0u0QPfXe9/CuaVOr62hSt2XD9oj7UouXzJpnfdWDb1y
NEhfF5Yfed58wF3QKWNCBUEq1P/kHNYaJMU3npYyU1cQGj7s01lxTI2IYLHBH0x1
EwWwQW0rQ7TOVJ+Y+59jOJ2gCUeHKkWZqQUrGELMbqpSjbnxAQOGO6JHK0bac+Ph
Spn+HLtyhJv4PGY2vmv+wuIt05reFxFVpHZQajgZqA4b2W8Uf65qYyzrgDRJcY4L
1NU40DzQxOR0ZkpWiVyqly8ztugbvhzsDdKn/r0TD70iQhp01EPzbGLIl21hDovm
6KYtLuJbNltsY7WZLmtAQ+g+1VHbsnOlgJ2NseW6nSABttZbUOB3ahRMg1pIPrzc
USOVsBLHXiUoIPsjX3hfvjQ0lEW2vv9OqGl1ryQCoBBx3IEfpQ4OKZbrrttYZK8I
hZnktr85dqhlIEKQTWTZMGFTsakuNFlybri/JStIguos5qe1oSJvUmoGr4XfeWNw
U4RWLDJir/fd2aEqDqKo+2OUDrmCdKEqDu0eP/nlVWtOIbEN6nukLB19dceBce6s
C9RlxFbk5Wz52i1GPfxtHdA4tN/D2HmOiSki5eRPH2NzuSdAazWg/pH3NChhq2rM
RGpSc7Y2AlLGomr1aHZPidctCIaRpVtflCy8IzWH0p37UTqN2tMlJKIrkSwnIoz9
tWN2N0TRtKvesQW9eoSOB98F8TomfaAMNd/SdqDNC3R2ZlT9TnvrYNw7hztuqVg+
mZ0iahhfB/djbeABl+xwm7XpWspT/wZx1Ltq53SYQ58gVGW5RvDjMdbD8YEst57A
H4ZZ5WngwgpYMqM63IWUz3Yv0cr2M+aSveuAWXrTP2r8lRAwF3NsAErpoREaU4zi
/7UluOiz29EsYh1hFDpZ+cujtL4K8iM0CUAMm7psrdhHTR6RWiRScm3KGuT4fTNv
mPQg5AoIXcJ7cq67xAiQorrzH2wxEGVsC+GgKhIpuJSXFaVN9igrcCCiZ6BgDRGz
Q4zH33OdBtlkALdrlp3ybO6B4lpDV0BdmeYrQjICMf57D49i0MWecmYKmvwlOVSa
qoj+lBDQklHi9F5gMLozJ+8BDT3y+arD19j+3akJ/WGPbZJrKFY4JG2AfOC0LktE
2sVN5do52Obm85D32l6R4v9m9ouTq1fcpBbw6egca4yg+QiPnOGVCU3jdPJZ8FUq
FQBRSgAVJ0vSXpRygrTniQ8D9E9mw4NLmfPggIPvby33IXwfEma4OyXGtDvnns6e
QfpEBYzEo6Iij3RVW/v9ieW2vKxF0x62v86riFkxGHNSUeWaIdqDHpdv+NRjLr73
7q8UO35oi7iR75DuEco8K6NgvocLpMynvZhh/6hJu6MarL311QkdJrQX42vIjIqu
zwwRaC/BT7VEEn6Ai+WmgMA8+H9taeO5O1PyOCFKh0/tQ454gB1z3VCfUGfXmK6Y
BfhjUDn4Sq0M0IOXz7i9B/8JW6vELarH/EkhiFhC/15edb9a0cFGy8DQjuZU+nN7
43F6Xt0yiszIQF96oNU+dV1lvJmbqFWaMxdmLmfFfGshnOtNiP+0csBQ3NEpeZZj
TSCSvOMCjwgpm9xTO7zIb3phbZ63B9vNO8k636Jcou2wdLePT4qxo8fasNJUPB4A
bD3vI9SIwzTq7MucPRIZ0euLhYs41OsEAByKXnOw4kxNKhZWKU8kfk22OzgGnsWv
YNTB1s4/zdQOn9aahlzvqLvroHZs8dmybyrSQ9bvlBpFlA/cZ469dswFVLshvPd7
09//S20Be7dQ4BfoNwDFOycQ8A38sfLoY1xKt1Hc/VcJ6Z5QlrH4imbQLepoIzpI
DmyfsA5z2SNtFDkt3ff4ivEaavr9NElIfG1s3uyE8fn8aQIK71da1ehVLcL7n+8f
dZFySNCommq29Skh3cV2aTKQsewNY6jlvS0H5/pXySrA8kUDSeMa8Q1S4/oUKuoQ
CjF4IJdBK/t6DrbLjFJxf2cFgIK/inTo02GypjrL1l7IQKU44xtOEYKEV9cQ2paG
CXFygXof0mzL/rvxJErRXALARxYcLFhEpQmOtde9S9NmDUiB7e5yGlcVAjzMUvMC
SU18GtYKfnMLdd9EQlJPNglCOSlt2ndicYJPhCQS+jWyiUiBaroiuAnOfY00hJWp
wyxPvTnwP/Kpj0JHaSh/sIs6ETkpy1Hg3nVPt4/HxTaELAkBjIx/vSxBnLkBt377
6REiq05VrNc+l80iZWuvaFiCxC6bdNBDudyxtvj6YLqh2EDNTjBOblTLU1TOHYdH
SeaqC4gyhlgt9w3QltSWfa59I4tPaVQFd2oESt51x6xCPhHDAcP5lfWIVB/yoL9h
EKUZVha5z4it/sk20n+rSoeEQr+ngfAC0bGLpWyEumoHf3PrjkMh64OcSXhBTGOI
8Z96eiBKB/p5Ik4eQdosIk50t+DSDLD3usbHOWf/3hUYU0EcBZg8LW0vRuPcgoYu
tu8vCcjWgKM14YfPZh0xCixJFYFPi/WMRWhL2iAf3IjItkId0A0eA5TwTOFVbX8J
CO5ersomgP1/rE0TiK276CCbBtEhE3dCqTkwtv7VgMYX6WvQiiYG7BKT6O3yWDTp
k/GM6oFtfxYDBCXdltaG/Cgs8s7zW6kBQl8eTGenf2y5j+A5iSrjfHCj1hgutxrF
GsA5610djRwARSTWAozWWlJ88N3o6dhS9eB3crgRCGouL1gMyM6H0ZcGF4d7sX5e
fZrcpPL/Y8wch6RcoTHExHMCna+fc/5Vy0sIQZFGAGTfeOW1m4qe2nM5jJqsLkQ6
09fRloKbsP+IP4QjM1fJ70YBhjmOkhlKHOCGjy8XdkVTYO1dkZ03Kg7GZKcWpsg1
B7Rzd3sW8Ds1BzMEYNFOzYfuhdx7VGLDT0voh5lOqmzxn2DBFgy4JJjt+JSphufE
lWvEp3gzp6E99TMbGqZhMR7+PsWhqZUAAbNxlGX6lo/tHaJ3yG2q3TTOBl1pGVqD
DMU4XYlDnw2cHC/E/W1D3bjVfR6pe30kVfdggq5/PNz4J20deHrEiC05VDd6ns5D
pFu4blfEtNXpnEZr9DQWFx4jmf0pTyfEHicM9NMAYnN69oVidsgjl4HfnKmkw0dJ
9kzTLvLWGgUbE8xZ7/PwuRQ9ggtEUJunrUKLZJ+y5ZL5yKxks4ckdj6c9aN615Cb
GnNUuCLU37+kXl2ZmWLfm3u4QTT0W4NFpLSjixfW9OshMFa+G2y1G1XjptUaXqXT
sr4V2fOOFTEn3Te2Ok45H23mwh0ys/LVvsSPoK04HrErvyoqKR5dIO5CNxWtZmTV
+Npz0zyJ1l0jjyJ/wIHhpiH7wH6tlmie2SDP6bDOGgELBmJmf9lbUVmBi3rVrfim
WLaeqcUkoDueKCr5/rijyrsgLPhWWRnndDaf9WtjxS0B89fnbOJBiLy/AEHzaZBv
VljeQDlHYJgxO3ZQN43hOEieicpaCX0DhfhVtlmiL4cZkxrPfEBiKFb7wv9zjpHC
NcsEeHlNHSwrBoBCgNC8PVhZp28nHwUNmzSXoB0tK+opUaWx5vXu87oRCfaH4Xqf
PsdWDWqY/nQrP49Rh84GEOzi3b2F62t504s6cEIzoIeJzHvBPX83coK3pb4vd7dW
1D8dlqOJH4gFLP77/1sN9S9E2j/y5yZ0qUzlujn3nnY6UcEvnsqFTtFOGzeFsDcA
EbygWtKotEpeMjMaD34eyJH7AVJ3eBlVe++fxiFQZnBUjED8XIIatEisMYhYWV3Z
7I00K54kt19DezSU44Ow0599y4xv9kysN+45P7nDXVQbTqtO4ogipocCaw/b69Z2
h7Z6/gh/hjF/Zbxs1JlNw5J+AWhKaPpA6SlQUMrGRE0YBlJcryAsQca/nHOMvqmg
dPbdgN2ORWYfRrmM60rZ4w8zaEftg51SJ0ckVbB8j9iL5nzhlaplXUIlnnH9I0us
HClvxFB4ENyU45Xi9VmvN7zubPnBSoIeGdUGL/+7C2D9zKpwjjLVVYXmdPYeUnC6
wbN9z8NkgRWipC2UlaiFt7z/FKnDcuz7uHvo00lKpU/MyvQTW6KEhYB/VLkkd4lv
01XpfoVJHmezjXPQ1FXeCESpekxNDP3FbuWYbHZJfTp61iSF1ddAJR3HIxLEcLae
Qn12LTLEb1p/4gJ/F2iqYNLIFJGp14sgu45wg3J4rlZXYNz8VcIMXD4vuula0Mjv
UceHvMNerXYbshZ8ScdDF5WxqJsW8K7KjPR3CygKshR9CTrxd32E6o0ntE2Q9und
gT6+9Iav9JGU96/llC1Foz3Ezse4uKqE6PKCACLGd3QyMnyItH8JA5YxiZfcp8zA
aD1/EbvSvdC8IGML9KkjqSLvm7zTpNFrjGnaFH567EO2CXEdPRXCNt3/iO5P6jEJ
wK/KkjmXLI2FQWQs1XbUvrVj0YH7kwudW3O2xsyXvXjllDXv0BBDtC4Fg4XvGBof
SyibHz6rx2uOlOcA8MYnSqKdUZLQDoPj5LbtUjwy6PIz4AJSTTxqX40QlVyv4yeg
2NPOcYphqnFuYlcbcGfu20elYv4hFb2x8AteKqK7FabWE87i7VMxmI3AJZzHKLfF
hS79K+L/FsjauG2qCHJKf0pkEzv0KZdoVWKQpWr6krodDksSDBAnpEgY05ozySCQ
n2daAj0ceO9rLpJObCM8wd+gbolOEelEKvtmM3HAsRRJrhgyi98U6uZMVoPlJDs5
YF9HEmNgdCCF9zXIDgVmSTUA6l24cm4h1ZWa0l4eo1sWSYLpLxh1szk81MpJ6SFe
9i2W+iad8bzFfMjkHxK4PaAVATQH5hy+lq0RGGU1bMpLCAXoPXQdk7C4amq0iCWO
1OeKNeQ2IF2S3QRkxWXr+c9wXpDldHczofzVGt6IE2VOA0YYeFRTim8URd99WeFw
eAakbye2I+yhH3s09Kc/8vRYTqOsClHmGin7zoTGA8rZ5BSf1wbkKrMEdtefxqVf
Jy96Uqz6IrCzkvlQbHnHwwDyBO1c3MmN269vElEWLzelqK8+LQ5YrAd66+Kc0lHm
ANqqnEf4bA8k1cM3Sdb837dOw+GE5dCBq+CSfvuAvBt6fXEMXboxOPWam9+gr8pw
K8dpnga+OtdApSakuB54bfUNpa3Hu3w7PIRcLFF6TUKMasVrPPDk5MiBRYsFcgxD
GKZ7K/gtcaz/7H/8TjUI4T88FX08UXHhx6ayMSvvsh9+tRi6bZp1ZewZ+zDJ718c
lXpRNK4ZQDsheKElnS4VyPeMEIlw27/KoTn5Ed0giKb0R9s1Zcc/ChGAENFlZyaf
wBGEjX1eyf28D44uApa92lez67wFTRpfVMm2oRO7e4Ls2FTyB9Ke0/UbnZzKgAC1
E+J0Yro1eVK3TMxCKyq+b5nWBIHNhKxFWKes0pNSX7u1Op9MzlKV1L4Lxh6ux59Z
K3MlvNC2MZikSJaKMdiBoABxViy/S7z8f+FTSOSt32p9aM1YHbMoymfVSUZ+vcW7
SFieS+4w95K5kKEy216XW/4hMwNsF8gSosGG5faHxR1e2pXVJG9uaFXgC7ZkSamU
RLD2kSBXAMde73miXz7hieAgT5hKeeqYNfyZGXHMkg4H8/YcUbqNFdKUKK4uZFV6
Bi4JZRdGWUiams9IBCHBYKHkesgkTa4J95mfvLVCPHz3pFcsAC4eqKKbAndoLf1t
FbrMZmHiZbT6xHcTHApAKCvHpc+XADNxiKchDFtZz7ghXLfcpEzfl1CeHzKaF3ls
BCgNWR7MEN4WzcDt+I1YbdHj7KT/p8jrfKbewAvKvBUvyF2X+HciOKv1HY0Lveu7
owGsmddStl24I6QJOrl5rjTy3tMIdxToSpzYFwusECbDoC3vTWoaKMTQXu73uxWc
xqx2fYM0YAoNS6iQCeXWvFafA195pmOekVv+bPnsjuie+JYia8JH3c+pFxt1URrs
QV+mnEzx0yRJ/0lQFkX7zOERMV4GwRxRpEo5hjS4E8ctUeOyzXooBoEL+oMgbiMG
81d9Wy3GIUdR++hMqT3fZHc7l3Vn6WKmugrIF2HINgik8BHoBs/1JT9f9sBueHdc
AG/r4fqAALMdhUnN1bz6K48kdbCGal/b8PPNjrOXb5wEoRYB4QeRGW3OocRaqftG
KqTF5QE2nVqhUI9rHoEGnU2MYqvJ2ZsWFLWLOiUtPeLFnmiu8N0SaobPOWGTFwLE
gIruDc2JhUjnHrDyVqVmXRe8reJ6kXkN64meb+TvF6Eg6Fxtuh4mBK0Tom8S//wz
53y57N0h8cInS94r+g/r6hZqiiwA9TZZP/QgADZbldtCHkdwaZ0ucbfPAOKw1/mQ
jB+4ca2B1KzK+xxrbyDn3vpHCF9kL2gFRUWO5kcdkW3kdSi0LDMvPUScdF6RtVcK
RGyeuknwc6yrdAwx0+5R5FYcWOpUiNH1vHNaq9xdEdUHupR+KF5DPGbPIHtivQQP
/lPc8TOy62d8AX+laNf5/nljdcltdigwF5yVugqzg0ZP1hYaWOhRbABL3i5PZU8m
6cTd70/v/OgeiWE4HKb22+sVXf799eYdgE6H1Zt67QBWFGwCm4LfeokcmiE+juSb
NHRKxAiIqUVdkr+AFRaPOK9P8LrOdgq5yaL1jNE0uoKte+61C2x1f9cQ73AQ8n8T
h5PvoWObCsrq2MKzI1sfRFnYzCYS9+nNEnyMlmujE0c6cXlZ7DiSv/wuROcle4RB
+1O61Gyc3kVqrtW16f7Cx0/0WZ3Wep2CfDcnQZbER5Zv3kVp7LrMnyFAwmLzjtx8
gWIX3irehIBcTeDCvdirj3JSwpco6DT47VjSqEd8OFE0EomnfJAd6ZjMYepeDjyD
rxqm4tSmME3P6/cDPEOgiN92F0Yx991hT+W9yp4z0NGky0ZG4U/JaqMhn9NmkwYk
AV9C7M5gM1JxK4eoLDGK8lC52B088pPMJGaTYJwODozU8przkO9jf3CchPk+IwOo
vaaK6FMznkjpcjL3j5eiW10H4Eu6BSbBmKy5xBNf8clJ+RxugIy4OONp6wRat+c7
m62xob3LmW+LvnX69tl0DfsLCotDeWml+4QxY0Q0Dx+AIFoxw+ljaWDyRd0TceZ1
Qv7hYAWYCfNwYyuOpdf6aOGq/n/Ov7G6InbL0vzIuZtyzkoAqYeUxriHCFv44r2F
o43MxtAWFeDRSj49ddvCIkXzvS3sR5CckTipyfc8++zEpr2/F2X6cOpYx6ChvKIS
FfOXQPVLAxyaMDlpgJ6z+aiUV/Zpx5daRg6MpvFCkVT1MgSWN4Y764Osz2KXVU/O
yoBl05tFBmBTHfPEHNZtTRfA1/7fsJrSjkJQd7CKKGDEEuCh/Jq7wQ28mDNZyzj+
MBcEaQVGf6RmfeCkUs7O1S/QO57G3NSwE3A0gaw1WkrWCx8n92hqrWn3g4fheUI5
XRAgOTLTLs7BSJN230Gv+YzBjk36HC4xFbtjtnvUAIayGLB0X8cW+g8bP/WwHFMA
VG+jy1sQXDMkVjDYb5iUgg4r8o45FsKFm8zC6SCX5Gtq6BRt0yqt7sg0hkGKCtvs
jjHcE6fWFn/MsWqkEKpfisdIdM1EE3XXwUJdfEhaR7OFPLJ19FMKxtRPFRzvNskS
v5PwFZRsE/jyeHtasF8A699FYVab5SKuZy1b/ZcIrTl9jjmP7DtRWk3Tlge7m0b3
Frk3yD5FzDSejEtPPW9/vyzk4Xjq2tMDjGd6mgLsyIPPnQgSLiYr+2OhsOK6qGbM
fv2nmD1Ypzy550+qFwLvhhAu0eQg5yhz5hItxWDQE4rqHrnlnAfONhzIuDGl4gy8
LmZ4E+cuTJvcEZ4NL1W+T2mOdNjoUVdXq0ai9M4xk5HfJ+N/lXhxfZm6L/aumELE
ICqHVQ3ZrNlKl6ExQDSH2zEyihP+QftyVxHt57pOfpf/hZUXE/4R4YBVrxkdaotN
LsT2r47zT35OWlbyt5riS2aTmeXBodB5EpQH57gFTBQMkfYmSpnlHFqBVOtVtEnx
x6naV2ieUg83gVv2jJCEngByX6PFXlF8kUFyVz5QYZAg8emiw9uQrsPg/3VvSH87
ztToHfBr7YqYapjmeWbntagA/ZLfWEmVUeu89u4zSMlHCA/9R+wn4zd8Xbwu7dZP
eEEm8rHZg6e80dJUGr+dwGW8D9WxQJ4ha6xDMaA9aGFYNJqZNMfBgAGXM+zH5EGQ
yUJHaX7HVW10L1Gckwi07PMcEv1DhcIjCLey4LJx/PCx9t4EMVz9A0KA4qdDa4kF
Rkm9ntYhMOuHdueX2jk+3prsMxrBXVjVUjpgNFw+tTlytSXveXqP2TLafZppEFMM
X4pZIh5kSVdcaz++ebtQhxQBic6bi6AOigM6//o0ST8kiQNh+IrGkmmjg9kOeEpf
R38y5S+bHl/ljWYjsE0LBt8ZPB58vG2MRVOqXgZdCePj43/9CUyQEhOjFmQy1c2I
DX3dgrJzU/dt+o7U6pBvCOy4kRWJILMdlCsAsnpvipFK2qnTm3PxD43Lw2UnqTxh
FgIZUsMQtnxCgJuKrHWlbeYnx7lxD+H60CBkdvOW8HecRkOCojM7LQDk8IByWscb
hlVuROISEqsZX+hWwGIyVe56PzibRc0F+LPY5W/SVLdTPCVsKPMSp7FIqGjEW8u4
sY1T9dOyUTu9s5Xkhlcm9x7Gk5Wo9Yhu1pIbG7wLAI7WQozwhw+CQwEUUmlkbN7g
KQ+awTOqYkzoe0AUlEXCO9ZLPOrR0e1RD9LeAuFFoGjVeUd30dfrzJHxIIxi4qgt
QX6cCAlSjc6ygClJoKyRKXM1jnT5s4/J2F2A9W4vApzNqcpQoIpG3+QXf2w5U9fF
RlYUTeeotKt8eUhgfS+MR0LLTElQPwJ5P6vC50uIeTmQnK8AzYzljeJ9/uvH2RxD
czaZlkb09nqjcx2jC9vnWzz1MOAWI0IURzOCOBnShlWj3cF94kFw4OJlRwJ2zjGz
xvmAN61bp10NxafsjyrAm7rmUZwno5IYf/SkFlBe3by2IknXAq3zgpESlEBGqtgn
JwPicjORtbnF1BxbxpW9QL68S1gjYAEM4TCgqIX87Ib6DbznzfQwWg5H7tzsXWqO
dqrxGToA49uqoxsdrz/CGxJ24khsaCHgLnoYcDIjnmVW7lS4lS/O7eZ1z5U/mEh4
AsBz6uYEb8cdDsY0Sst5wYcrxVri6An9B1u+FkXnyp4ybEYuHDbk5KrmGfoOeLcW
HO077zBDiY5VZlG4XGGizk6pteo5PkI2DXh2oa1GHcCYcnPECAVgKLPki1B3ruQu
8nUHXRm+EznkL5cP8K8SV2XW1sks5xIekwWfERKyApzHAOlLzPevt79XWme6acw/
QKz+GNmeqV1T3CAzWt4lpFQ3vL6A7wGyhDWAzHdu8RMAN9hIlMiCy4HLFG+MbxdQ
L4dpcbmO1WS3VE2iW4kx+/Xvam1Ns0LX3WUfqoGvN8OWPj31sW/M1tMkuE0OWBZr
40QiLmS3MdFKJjPGDmLXeQK/v4RT+jNfUbReIWC6i8TZxmYsiVEjVJcGmxinTgLT
fasIGTVq2zYOhbOfhoMcA7MluKTzj3E3lL/x3J3NqrTuQ0Jz8n4vaqtVlP8uqofU
2D6LfspE+cpq3PYdFG8VYNKY4H+e+Set0K8DZXEdB9otn6h55gsdYNZPcs705jIk
B19XLTJP7zUG78lMTjkYTt+++JOPIyUWKBOZn0xaFNk5YINY0ad0AQBnBoQhZ39C
rNDnnq2OKT7pAUF50Qiihdo1LOaMcsyG0T01vDdWJEg/KjR+HJ2khLMK2XESLsKo
8nkrXrN37qGmUr+v/6KcBIHkkJpTYIAn4d7RF71tkQl2tOueuZ61e4dC/Lv/KuZc
Y3moxIupfKrt1gAg8digXVmsHmLHS3RNKCl5YPSpbMC+Se/oX+8oS+l4TAck9jIP
qCK2jWxJCSL71J9qxZkjt7+lNiL0CicVD2EYqfPV8H2OCzqvDf5FzXklf+e6dtSv
3JOa2phOUAzINU47jor5k+tqkdzgcAWY1Po/XFtFb412rcr837CA4zfthh2VW3Ar
YhL2os8blUtCtLa4utVfPlyhUINg7NsTeqQ+/1tU5l+mcyOqb6FRRzMdPtojAWfG
rok8taaABAdMwStggrsKXWFmKZE/l6mL4p62Dbg3jY3hh93s6PMkNGE976xz0sbG
MCWHPBgIQWzSHiaSsMGLjG6wwqP6I99vRICIAND0hbIrF/RpNLbVa5MFntMRPQ9Y
IfQxdeb17bUOtc74UKLVXjIPTXwd3jkzfSMCEM9ZJ+3onygM+3EM9qG+OqDbmveH
NnFPbRr1DiVCNprOnJzv3kMBRNLpFpOMAUrkprSG3sF7JtkIhwJ9npxTGV+dYhiQ
3OCZ1HXGaU/GpHBXLkHcMdfrQbUEvKJdip/jRoHGSB9a6N17Ht8bVYx48j6mUTJP
xOItT8oeoFcXrnYthvY1gf1P8REatjXHBphgeLSU7drJABHpA44+PunhdGSbsc3h
12YlOM3lFwLTzPtDkreemMHnXZ0CllKrI8fr3NRBPqSm5ph7biH3sPq2y0i4RLSw
tOpklD8rPQ+mrNcYxePDE/Z4d2YXtqMjT8TgAvpXhAGff5fSAQCKNnGZ27m7irLF
94i4wIgT8fGtYREhzp4jojcTAhMzozwl4JcT/yw76SZRsJYUMogb6Yi/UJbkLpoR
EkQOLiAi8Su/6wzXz1t77KGIC3uyZyjW60d2R1ctkMPnJBhiZX9kRl1PrkY0cnZ6
5uzq8BX5s8J/p8nnQDR/8+4Gc7UHX/MRcn8nvXTVGm8NAPn2R25lIc7QlyBwvLU9
1ctq/ICwHqcui/4nig5Si4wTlX2UlKl6ZIQO7SnmCetDl7XJc5FzN0Y+7IkDPRyu
rGv67ZPE1t+lSa285e5q3DCkmokFr7ur0IrqyzQ+stIZwwOEUsXz0AJSBsnJ0vxd
`pragma protect end_protected
