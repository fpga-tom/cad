// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
L5ptR8rOmrntfooLCuX5xRIB27i3TiYXlbCgKIHfe354eZOIKtOtX9c4L9JhAzbS
UdL22GLA4kbVQl+jYSNaB1mlgI0KeZD1ib8gUF2I5qzcAFkDILLhVlGzRvwIkAGp
F0V2aWe5lJOkEq1rC4mmfvG9kEkzhC8ZFoW/ZrEKcKs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11648)
l3gfIQOfwEoR4yVKpEoXCXKyxCweSkEoKweFr7lUbgGWY3p8rSf5a262lVHOs7st
uoTa68TEHtFOSm9/IKg6SzhzUedG9knvryj6UQiCPR7cTHr/koGw0fTtxhbkiBEL
5S90x6OtYrrOTJTAowlKvDew1l2U2Uq0nzA0B4/Np4j99iYZOsd+i3YZ89cGOFtK
Lg4EnhES3Nz8QkWrh+/lLm5DV/M3OlapghXcg68GeOdV0ubsCRIfYV5RXdDzDK3x
oPPoDyRobMinAq/rCTZM28/dRWaXzPlCe/prin67SV6H8rWVj7NowMbjXi2uiaeJ
d8+l1KQKkb6m2cCkB1AlfQ6WcKMVyoCx3uG+qQ70YkYRQAiXsVOP8ztWPnn7AvpA
Kzaz6pH71vpQKvk0MHCjyITuJpCyhgcce5oQsig2p/iExJhC+XQ/Y+iWJxI4rVxi
iUmSK81ynCfREdHFDyJ6XqGlEzV7vOTHiS5SWt9B6tDy7xxe7cKTlf9Mqr+xP6vM
m1besQe9Bwsa/QPfQk8PVDwEL0uNdRpwrdzIsGyUFe6L22X5jutcTXHPsqc/P75d
Wzn6kRKpk0tYkvgA9hChxxP8ztJSeIklqXVKqq3tF/7eGKJ7iJFEf41TYxd8pJqm
UvEZlb4Bf8hY+XKUZT5Gw1ynbBFT1yBVtXvFMnseH21Wh6byuYgY7wg4D4SmkLe3
xHjjSAyPfUu37tgja5cXtF8D9awLTCHUBRUeysYIOQ/0GGiWurIaQXXy5nW02wiZ
Ofy+QZ/ix4Zb46JHUNwDPcZ9+R/AJOOg2SBb/eyckAw8Ha41R57QFUmtL7C9yAwf
F0osT25K74LBefk3rc3leuiDXQzhE07P9SQcw/3P4iuf60ut3cC4lHEWN2HcdKGw
h3ivd2jzEWunvWepSeNrFAaKHoYcMqhrdes97Jak3CYsrDUJsTLiBrmIvtXWuz2w
LRAlAsUF0XGOnkT9R/5CHhwccRCAVdsY1wDe1fi270q7UrXNUcJPUErsQuLNSJah
4i2LLHigu+o4GWBAY1W+z4IJ0tCwvDI6w7Rg3G+IzNKbt+3cy+L/qlwqYLKL32Zo
irxt/KeJD+1rzOksuT/FqLqCfzoOvNJq2GkyXZdrPOZI/i76Yjm3JfvCSNZk5YJd
k51dzWBDb70XrubniZM5TyFXD+ZNSHuXJxkakfQSpwepFlZxP+cuewzDVw94PBJ4
gVNi98HIhmcwuMzwYrg0758nyR1IQw/ldbqHuxOZOoUc6mP2EN2gtzzM6wzzXc3I
ji2jmAChtDrqCHamR0AXWQ+EWRcQ3WFVOs5JWSqG9gqRhlGPp04Xz7sXMwusWLNg
dDnnyNGoFH6w6j3+Z/oOKrudJG85IunN86iuA90XkYEJU5ZJfzI8iC4CW/kn8D4y
b9vh7AlrStCvwPuA3sVb/ktWCPsIrKQBZC6bqxvLu4lSlkcrtBBVPGqbCtM7Q+yS
z0mEE5IZECEvgtHjfh1zzUtJXOZXnsgd1T3RO1PNlw1MlaRXZJO1aT2AyYJlaBm1
27Mv4x/vP9lBEWAgN1qJWGLvacnCTNloa0Z+r2+3BS8+ka7T1ceR3j3bkTeWQPTL
fTiF/kyvKruQZPfGfVrH595u6A6zlBzwCmd7dkEft/HSXwFP2W8A8TFrulOUEHpA
+3bhVLuDGH6xrKwjRGtylCMtp+AIteFjBoxKpoOtNFjPhPaWxHnztCizw1lhk7pX
tS+yZd+qq0gP9VHpLN0aewi5YLfk+Ir6QthkvlxtJqAV5R/3l2lM5uI7KDJGdss4
8RyFRRHB13jNfZH3TqL6fc3xK05AjX9yTln2Bt/HLBx8XLvMJ96OF0mLAUeWexZ4
LXGnrFEVKFDmC6Fn2A7iTx+WQMiMVwimpo3m4L8g4iDVzG3+6ldcpgaC9Qxkcl7g
U9awAFnmpjaf9kG8rUQhO6npP1EHiSN4FvUOYs8hTtTIGqFDscMaNU110bXAUtp+
lxewozZp+gkxqtNN/S84PdHEScCpHTAbussiQ0YAKKhZXzcllZ1K6jLvDMR4TX6E
Ilvy3O1ABgHbL3M5QSnxDVZ1JYhs6r1P7XHxRfV+/4fpaW0vmWB8/lin0sa24uY1
EDDbqAmknkYJ1N6BewIpyxnBGPSd/Bdy5lxKbvt/mcZ/Yfkj88gCthYW6tOBrOEz
7kZKLpvqMykL/8r3J1VHCkoxe++EeoFEftp6k/vpkHIjIOSHZSj7wO/fbYgxq1ap
lMGJ46wECVTX4Za/4mn3sgbSkj9r6SKIKeYDV6lvUPEE3wID8COB1N4Unnxn5QT3
jBvBm15ObwH+HQgtt77PViaCPBbRCVq/xwO+2ndTF2SVYXKwkTrCl4hhUi57BGAz
sfNWzMM2AXqVFXOmujtiR09u7RAfZugIXQFm/VZJVYExrkKOlhI+I8XIAXoVta/E
ZSQyVwErvgH6FEkK+p3tyIlEaf6ePL80OJ6gI8ygfAJ2n8pK9NETY6CvfaGYqL8v
4lmmD/C8wVgxV+uM4PXGCCRPq5U55rmH+VgJO0AjuimVNAhkoon0GreGRDbyCVfF
W8FdLa2tTPNubprht28nnFi1FRiEEqAv6Cs5JTqNwFzQNG7b4O1o5e+n52YSbOmy
EzCNBdFoj6RnIJo12oeWULXo8chQCv1c6CXT4QKCL8uoPUUmhOoUgQqV0732BCJc
oWb7O1yimUZ0lbuscVZ7UiIQkOLqA31U2pgR558msyPWNmNXiXNQQrJFRyyUInux
S6GrRAWSkwV65b10/sQ73J6G9YVcHVMEZZJOGrxnMEY7Q/3BN9MoSigXVrJQ8IoQ
2hI7fDgTXk17UivcPX01GPTdmyw9HZ+N+B+lBg2PG4LPFxt1eZMGjW5fjC3zur4A
uS9k6TuZxjwLplzyjo/MawV+4MdhgdmXERkQ3g3GKqCXF/BjY4mR+QEMpVyZYjVb
BHPp6YUKec9VMhbh6VdFUhJI3FfnD+85SKxnmFjZb1707TDuW1N7GvpKOdXGs+lj
EBwuFP25+WSuQyT3p47EYXHlGlvAr02rulmBUgetwie+jQkNI5/JuA2C0XFhCSo9
HGn64uhj6foA9DFu8POu6y+LLr1RdXWOt+yImv76YpyJUc2CozVpKDx6IkUhKdie
PewRGKpYVfd7wJvev5clTWUDiZ/j/eMgCvzed+lzYOKnkM1qYAZBfLURV6NSI3/Y
/Z2M8tDsiru45Ka2Jub8aAhqMVi4q1fGjvHMZm7GeKoZbqdgD2MXcSaau24IzQIu
uh8bCP7JqlDlUlb5Hb+bGtcV2cpqOXu+psBvsdOtvQpXollCn/viFgSNIdD0uFRH
vOzwFiQ5Uzg4oso827o4VwytAlWhCC1b1FkJY5dW/FbCfZpa+57+S+h5czD67PaR
YLgH//+SkrzT6F6+mz+oKRF1zS8qjDXj7cVVJHSo9kwOsQ3i6gaqZCosrcpkrW6b
XqnzcIv7lOifs0EARB9aboqU3QvkKpFHw4glNXg0cYudIEb4sA5Z9qZB4KTZUtKX
y+zqH0tRlZs96ZcIN5oNiTFWW8OnC7T9lGkEtf1FtrcIPwLMMACBdLKSMLEcZf25
6bjQVWxBnN5rxspPVB5jYNxfek32GZ0tqnTbNV3794YrAk0Xe4pEkL0FTaK7KNpG
gGahN22sQUqn0gTkZfq48eIUWRyD591b+NetHZIiVW4HRiV7amc5meOjQ6ys7V9O
wCZI603TMSA24kyeOVR8VK3mEFYzPhqLwvOYCXZ9Hk+itGWgek94rjtvldudw+dk
qTwY9Ub8PJiiI+31w5jalh974Vc23b2EhBmt81vlN+9vDueU1MpkigHkVmU5pHFo
bkr4xTNHWtqfMC5NSLZMBFTeWKdgq0vwFFS+gS28Uzwz89ip5qiL5puakq2odnXe
Y78vPS9Uf8IcfltnPzJrmZbvlZWJhICXq7oAvikcmh9/DftwYEE7WZYT5lgii7Zq
+Z0cAYtUVHOMnn8/Nqz6k2BjRpKxC4wREC1v0jfoBv8bfCNNI5tkAb8+V3It34j9
2HC7JUM8zESo9XnaXPuPAe9s1T+hltgX1uXSl8z3bmvaKRvbkhMHAhCbFffz+Q59
+gdOrzDlcNN97AhswEWGfY1Rtl9cEXaXpaUo+gnaGO+K7zIijfy0yYd/7P0YGumM
FoNARBkDvgA37AQTRoGYL6/cYbyb4pb8xA2Kgp9OnN1EaTZpz5JN2wSDdn4Skltc
8EYCDGoZk0EMScJGwzz30KQ95eph2HAeEZmbyq12y8p42CAmorrNpgwmgKGraBQH
DitJNlFY6NluMe2hliaVYw0fgi1cpSkSLBPtXQLmRqi2YexBvSf9sFkin45q5iEK
ndId4xpm1vHQ/t53Ce9jgy8WxofJzloqhB/F8557PWX99ns4eXMtwdBHPymfS1V5
3VnIlb28GlxDOhrymrqyxWjLgp4GhD3DJr/4T7yuukg0x98eut8zNuj2ztADVTfi
xzA1YoXCF3qqdUq4RFFKHDLr9TRSYlDbZ5ml6Ua/eAI70KkOSjNt7ZhESffsRJT1
1x4tMDJ/utD3M8nTEALsOFjKrbN7e3FSm0qpqr14IDPEQ+YfDmzxR+GlNZrRTl8T
tb6vdXLMcSZiHFxhhBEjhGzDTDjhVQFjgh51NvWqCrl+MF/bSNVpQi7cyPLP+53w
rfiLd6gpGlE+LnuvwIBAYgU0Dbsqbx2VQKoWdvIrOkCmHH9OiAVBdafPFAuYS6zV
bn0lr349MGr7hn3m4jSwfOGoDl7IomuI7sQxE8qdINC0jRH+mWdN93dQ66CIL5WM
SNnNzby5VnOfeWE8wGHV8VNZQeVBkZ7OyRpD/1TQ6W4C5HrE1eN+ZzdFMIZeKmMl
5yb5jYfGFGN7fC3lszvRVO2SQWp9QGoP5UBWM1OxFRRweZc43YoamQG1POfeIZ8x
7vrMuchdigS+PMwoJ+9B0Xk6sO69gKSfvuoCoeWfy/etqU1cpx0RrTTZ1bO8stBl
Zp+LkM66O+6f/wenc5oEgM/7PsfOEdweiZQmC3CeltNI3fGgT8XhWc3hyskDOimI
9A9raTh4fy9ADCZ7S4MSDSCCR+rHtLeG/iXpvSaiNhoc4csOYIzLkNUeVdKlzInB
/KZV2GNBmetPT6/iVqsRDXQTToqCaDrQIy8Ci0mhFanuTtwADGqKgDaquWYzgA8X
fDMZlEIZFMYS8+iO9MysijimXHCwBMQytye+K7LVpKvfERLjaHctEfFRFdEGg2+I
CvSBqJUa6Z1xrAI3/4NiSB/LD0dFUQoSvC0NcFXP/cndc4+4EL++brAwX2+96Tmu
4Pvvx10RnD4qIqQZOFFqoKMhuIBZRA4KjeQgMshrHU/SrxvUQzdCRSzqivgtXS6e
niApeacNE4zzDZYcSEbZfZ8leFAUHca1wyZCNXPwXnIizcPEuw5zavbO78KXIfV0
qnU0PEpQuDGdJ3lqjogvPqzbeSnpp9G+V1J9iHcCyfjFZy/brA7NUrBCblrcFDqb
PkgW35UTiShORMONCUSxsiefJTsxBVMxiREiq+E+RDufDP1eR56iTnpOZGsFEhpW
VdMDgCV5ZpWmZJA8m2r1mGSjYBK9nBGZqfpkK6J9RQ9XDaKBvtPbic3YP+p01ivn
TdFg8bY07CetMwIN1lGQJO/7PvzpxXfrqT0DhGiXn5ds/QAfHe77TK8YAqrG4SKX
hfC1aREoViHtrkiR8fW9AywzJGG0HbJOar0KHB3U3n8foYXjnsl5Tzu+YJ4BLGZx
Bcze8Cbd5OHTy0WGoIV0iz+xSfPm6GQ17LIzNPh+FofqWVR02n2oB81TsnU2HhGf
y+/aQlAVFDMYAd56lHBlivOYF+szQk7lGJqr2DpaXx9ahD0wS3dFxvQp1NP26hOu
TY9Xk6yInwVWQBEiNy95MEd81G4uVsU78lIyEsuUnfvKuVUMxsyihIGnoKOsGbrP
W9AWO7Ztsep80YQ6US4YO8TKvEs/du6/MdPurQY17dS4DxzPmKHlw4j3PfqRAmGy
PwCbFH3Xn4egi9oJEQ5OxITkkSi2+j2PCRHZNXVNr6F8Bo/RxvHSU41XzEWfjAcY
EgLY/rsNLvGXjDeFyiFzgDmTZsd+MNMb3bqL7osB0rkgqCketONa/B1I8pA+T8lh
J/9/NGtKMS+8w05kCqKr85bxhuW2gtPRf3RR0dPbjr5AAYLDfBdkh7aDiijYU87u
zNurr9238+pmgDwv8ETpHOhCq94zbs8t37VQnJs8gFieowm2TZPogXS6TQ2IfVRX
ZhL3IK1nQH6dQFxMaUSaJC1+gbtiSh21c6KFFXZ96l11A91E8dnlGDjXUeG2gDZf
odEu27GFQwjEkrwZIxz7aZVpQMjrQGAeJ9WW2iy57lEKIm6T9pS7hdgzCT7pds2B
Lr3THXWr9qCvjIPJkq/KoDpIiQWPY+4qSOAWUS94yASVCKl6G92Gxw4q3zuTxVZX
Ox+mOMISPKMty5YN63eb602aF+2UWeMcMwxxxojgjsyomXPzg818+Cm+Ud15wshP
BYi+Q+yPT+g/AFO8iKGrRFdAGdiQm7X1p0ZIFVSKGLg/WD7aWrcULATh4WQ1QWSH
I2WjDgvOCG/S1cHP1Zm+8mVyVFYlMZYHsx+1hQrqXcfshfKRjjBEJI4YpY843kPz
42JX24tvRepgtNPtN/NTFvAM1AxQrUhVgoNdomuqzN1swsh++lKRsW+SGxDYy31X
9pBBZBsD+lR/URiNUkufizL9+QqJXGIP8zCw5R3dZVxYGn7OKVC7j8b91wSUWX5O
ZZlFhIEMntZOjnuRmtxcsJV359mpWs/+uvqRm90FgZmQcKqvKp8EKf1z95mziv+1
7hWjoo41yZ8BCay3B0yqTnvFsxiHB6rMoaymXULBpoL2ZvH8Ynpk6gWYnxFVEy6Y
pRJJrzFho67mg08rfq0qMCxT/vG/tZuNdBVEtD189mFRF6cC9rkUR1V82lgqt8aJ
J217PJg/XckHGYJ7kWP9Ij4RgINODNKynIHvz7X8X6YFUcO1VJZfF6Y2KAbin/B9
zYLDs6oim74EbJj29s8f9hZj2Yx2/ayxIFAhFjh2ya/kDHQgWzNA9FJ7xVBbwo9z
JICXwI+QP4yhKLuPtsADN73MvJAYgfUY3UA5k/uVqgH7U/krGtJRa6nVl0dO3RTM
aPHCbN3sdz3OTJ6nYPFOxCZ1pxKBnNJbyezCWfpjN/wZpPZNUNc5ZgCt0Ir9QcyU
KFLPiovgCyCXTm+eMYyNYKWNoBUHubdcO+8eaiBtJ6XRToM0FPL05Y3G6QF+eHb2
LnM6yk3Yc/b3F60dbIb8J3prkCIB1nALVGwUf3NIl2DnqZpskOWxjdcaO8MzDgC1
J0Ct8Uj3vitd38ZPCLZoKbRLEPjaugLct85dw53plg168BtblYVFNIj2vhStMNNS
UN5sn/xjiePojW/jkn1sXR60SQQOkKZY0ae5w8aD3x1zZWMQ+1fTZLU3tFi07okP
2CQLUsfJ4j+/+HD52pSIPQRAa1KQlRff22G4cbNDKihZyNDAaO8s68voA879MeKl
lXdkr/d8VGius9x8adpGwqQjaY4vEGcEwYB2209sGaGZWGqHHHuigaCuce0SYQLx
z5zYfb3oEWpdgLf8g0LPLprCcmYrNLDL+jpEBBEmOmuVXgzsAYBY1ot/H0X7Etjg
NWwexrXTKd2grsEl/EqwsFdTSiV2jECDfQdP3b65aAQp0DFuJuCIteK0FE/oesHJ
0KZJDUUSFqXAt4/WP1SzuWDm6ySjvQbn2DD4quZqp7NjRsflwjfJe2K1BTn92DAh
rwwdprE+tX2iLrQKhJVq9lADNV5wczcK/kvzOMST+MUvSt8RGVbAg2vU6ZBV6tA8
jsN1LqLEK0JPKuzBe8/xEwmqs3axebT4urKxcA2bNIKBip5Mke+aGJc03DUPkHNp
y0qKMIEM1Tt3pXNlTxA5CZY/2YCcJF3wSaCZSgtLkhPR3MTI9DDGxHHBEhsS2Sd5
zolmEVrhX2j0+4wD1Xo4fWuKJlOnEc/1smy6Ke+QcGlmLrnj9Oq9z1p4yGtnILX7
vXvDOnlh0Wlp3+IJrDdgcmeZMnt1FEtBK8RT+jXepGRp6GI78iQoeG1/UOnPgrii
hSIRamh09ghsKldupxoKt8w4ocPKf4xlquSxS1uyTNaizigP0qTmsZsHFDCHdxoB
UQylSHAIrVzL5srz7j0UyD4t1ihtfiv1i90OgvoSwGXohKOIXmuOs9Txr/pnxXWl
2yvAN7pyKbRwVIrZ5OHnegFZThTh1RLBBMfXiuPbH9tFNr6bjmE3n7zBIbaJaZKB
EkrWrKoMdyEdC+Nm+NyntzJ5lZaV/c54OssGa7qLEtoQTfD6Xu1+zfgHjnWGF22K
G2PfTEHDMBr247EFKb8L+6wlRrHA9d2NvYxiBJsHEmy0XQ8hHmtfDz3sIDcwNtkI
S6D2BYgUX1O4BG6bJNtj/52hhoqxEfVzfIyol4S8Y9HrZ0EiB+m5SZgHnMEctM0P
JfQikBef3fzPluExxO6qvLdTDjmJJI7p1xMDsE8qlSznJ8PDEoGO+8xfnsigueEo
TsukiV0ph0AhjFnSVb8uAmwBHMs1Xv7BaqhyQwUP7VbnWeY0sZ5ghFvuv2kX0YXx
UYuHb4AACkOrA57rwgj77bzvjg4tn/4E0eJvrvWyC0E2b8NBMXqcsPbuqG+3rWqe
MCqXFXpIqyS8MFdwfAparsGAJFxDzgxg+3YsuEFsYBi1f72MUHLyWIa6nFSe8qI3
Sj8legco7MEA3MJ4STSyl8QICxN4UXGDDvh1JggjWJSeiMrvnkTsEbhW2rO/MscL
dCeJT8D3b1LjeVJG55hcsMDOkgHKDN5hQBTLYLmO4tHHu4cO18W5/RiI+EWRp9gr
CcfN7uXz8p5EhZS9eXB/VAZy97GNXGZdC7Lr571wm5i/sB/wxfGG2TcNvC9JzJds
iIxThIeecF18+2WASd3+NMr2DslJ9oOeIN38QcDyp0mnnL/ozqmeY5ZdAPW1Plgd
n0ylNiutI6j59Y6tkGu9SBrNAsCpdZPFSnUiOLYZ81WFuvyJzE7imD/7+0WZ908M
0pRKDE5dU/KtLfKFXcflih9sz6BmH67P89Le2BYc4fZWywxqD8ZVt1I7Q7/DldZS
WoYGmWCPDO5sTGYOlIq6DghSzogzJoOL0zHIR6QqZsB48ZPfYUxdvFesQ1a4ukET
cy1LsIpaOaLQE99GyOgEJnTJpz3phPKXRziZS0+zGMLGLnApuYVFWPvwJNLDpmhR
EWaFsTX9VKAwjIDscKGG2WIM8vlc/YU23f/JKqrUclMUZOFF2XoWvDuOIGbpLgCB
z4rGFX3wl0ASurma7GjgUmZqwC67USAKOidEi/YpECRnmaERgTqgvirnqMg9o0fU
EXStfw0QX9qTbcqCL3AVngjMGvxdF+uDPaQjE3InE/R2s/s23t419MYMmWg4V5bi
KlVNnvJTzCCzd2TOeE1j8uxZnTEptPAkeAyh1/310XHs5cghSneFMGCYb1ZToi6O
y494i9JqvAn0N4vACYDwEcU89Wq7yiRGsrvt4Ciqg3T6+iET6ZtLCHk/Rt9XCI7G
QoCg7DvRJ1DsE1KY6aAgVOh/EHg6pnNwUb7TXt+yE+Nz+ObdMj42zX4iqivzF9fJ
rKGfL9qLTKGBZ6eROLz8K846olTtBCkpmB5QQTw/4JwzF9HFQaroF65XQCI4hyoj
pcHIQzwIr6J9Hz8Ukq75Q4m6TCHESlSb0m91jawLSgfGYmWRiNWwrvBJoDKLp84L
E/saLnP1wi9hfjOnc6UxJvsz27szr8Iy+q1KevXxnRVEy0YHWphjsRRTJyZv+11S
vmLpj1agcZr31R+10zRfIIVlyoO7NWMa9tSDq+YThBUeSrMfxaac72KrhJyDZnwo
GcwU256Mm7v8K61KTiSEsMoXJLezM6CYUux8sotohmmKNZtWN++c74lINxo2Fgu7
iHvfVm0WGVGr/m/g2EvmhM8HtbzFM9uOp4aumrFycw/TeX0WihvgxI7Cwyi+1mkS
LFK+GZ8wn4kwYGI+JUSiJZg+C+xYOUNAtsFbUKDxna6hSfOF/8nboUkTMbAulKuS
DWuxbMDTD4wNv7Spv8Drgta8iw9bLBzfAjHkkveFf1JH5KZ13YEMnFCXbStAI7fe
A95mbtCnYM3UXAJCRpYkZ73tEeg87QEeJtcgbDCZMzVm5TGMcsd5aPC4H+PP/Fvx
A+cZAUGScSDft6biXaKE68kItCFClfXq0MpHqy3QYp2wYeENazWxY/U7+ue19YLx
TCXXZjPcUpu4mKVsRcqoDMqRNJa0/0EMHvA1r/sDzrDcO1b0QZC6I16c22QnWmPG
0UK6goYWA06H5tmAkW/ojhN/o2ItDFCj5PeDwnSdQb2j2cOsu4ibQXk0t67E/4YY
V4JTIqJnzQRr5hMwcMqqKzqRUVoo7WqHhZQM6sVxyn7m7fPrZWyoy6FEqTlQQg6s
DqQWM/ixIJQvMOAZASffB/CAm3z/NTe/oD7Q3BC9DjKXqXyiIkro/SUEgV0hCoPN
JIO03uJNxDWzO1OmHWiGiEAQzdmBwFD2ArF9drAwP+D3lw4HRqXrobJtmIeRrdbw
VFviUKBYivFdanxsetfA1hft2VGd1aLdNCgMQUYMpkMK/K/NxQTaTIC7t1Wxi7y4
vbV733CIp//S4MzMrmQImEczMdMUnSQYyrLFEMpQE0EDaFUp1bvSsam8OouTk9/j
mo/wGuhJS0c7jhZEvkXnU+DojpoB908WKAigztIqXEdStCTS3Ty4p6vdXtQMWvRg
ykw8hgPOK0FuFdk1j29DsvyqAViZj2IfEa+CLEsPayeGA8m7H5nKAd6/Z7QvGyv+
UdenpVBCdtxqeLWNdt/UXU/T7U9pktTNoLjJDaiIx6sp/yzodqyXWJP79xvWydIk
UsDFKhaM+2pjnZ5O0ajZZ/bK3cdoOJJGboGRWVhymoJF9S9wNYjFoCCYwhJk9HWO
M2DRe/cpBdCAo0V9TKfb4jj4TjethWboBY5RPBjY97IWpHMmnz+dCQIy+g/xhPFC
3qEyeX39G0YOC4qi+PAXzyRx06eIXf+sdCgjDu9IgV39x/Cm22Z7un5T9XKoPl/d
iZOi5ZbeagFtdeBZ0hOfOd0MgEao5WTcGIov0poofRb9HtP2jpny80HLzE1/OFBv
UHSPl6dFwAxscwmyI2TRP4peWs2rVHzZUp44Wmblq4+tNZEhIDs8vpgPw9gP2RaA
pCu8PvFJiEGeSkPaZ8Ey+gcZqsLv2FGpvaMXJE+Dyz1PoUVEuHUzuRxAnKXjtF8f
qMhN+reQMWLXBNqdLJiT/PAGISfAW8GQQClbppBRLNHIc7MPZsjwuVBe3pmF8y3+
izAoSzz9lsmCWc6bhEkt8XcABesRcc7TmPUx0bWCcoO11G5k4JbDmJHFC0qKSw8B
TkHEkITQJYHDslG5WGz3uyVYHeclzjVAY7KCJ1++C2lrCe3loApDk7DdplVrsFZV
UhBN/YiBN9FGS6EWyh9TIf2thQntoON30ji/7cSpiCOhAlx3qDw5ZrXtwvvPGMXq
IlVtaGaAnLR/1TBJuHAy8R2u44tbi8JqCIOPAom+onpyDAMPNLM3Tg/72XEvrbLC
mcLDRTDfSPEj1uNkMvF8XqvTl+Nc3EDwsW27FL6WQPMLpeOlnuAQ0oUOrybBQRYi
p8vb1/Qp/gVLdTZo29unF2+U5uJX1ckcaO+wvm+DQ5EaNkx4Tn/7nickHAUZwGL1
99pmfDqVEIrMSg1W/ECgFRgdwtmVoI6cf81u7ktMOwCu5GT7Cs1Kiiy7UB4w+69h
fzWUpJ+VYeFqCWQ8NgJ7Z56I8QyvbYvKBYvMbZtDvk/zwAs0JLdVo4NDxwywaIMT
5ivV3QUH7NgUu45E0xvMEUwtANikUmAZCR2v4Xm9m6D100z75csE1ykd6IUbptrl
3UVdXHHpkqQJ47eEWD0QTxo0Apd+XHZlXsaj7QrFYUktn/UDWJg2cueJaltFv5Tw
bz1fg8y4GfUSO0jLCxODh5OSizsoxZ1axZ+Uu9rZhfeDry7PDiHn7bbROY8heWUF
CZFI1H4V/6XYzA9jSD+A31JzYL6Jt5yo19/Dm6hA5WxC5srgdpwjA4els84jbKfm
UnouEstFLf5ddyes4QZVRQk1Es/JF/PNo9QpvrD9h1R46fUvCT6MYzBD6ZKvcv+k
hU8UyArG1SvE1j7vg2vqJsWB62rJb/NN8SkWgN9GL0xFmfIwFTJJwz/0prbmG6FG
6vAhAFMGP5n+XkDgFCPebunZmb7fTFy78l9XhBR5xGzTap8hr4Anx0s9R4t/XYAY
1pioeaJLr4bLnrWsgxO+Cr+ZupHH/e/FRpDd62MybcIUIfVrBJVVGRyCGguZcXDr
D9DyJRBY8b4H1QP7ZX8s5ZT0EaLebak7uESFz5s84KTqttDKzcawpOm4gs2MlGqT
MMPYA52z5hriwT1VhV/5AMtT8DIpwU1FhYf3W0W0eGrsdJqSbzrwy8IOId/D3fgA
GMZiU2z8PNOywJ4roSRyZBnnu1va3tOK0x2Dr4EZpX6k+20IPjqrSIl0FG6/dD25
wkTkU6GiRzw1dxvh+RXQz/nRot5QRqBwwgp7+SLb5R8tROTi9e3d79WfJaMTbF7P
jA/1zwjokJC+DPJ4Das//o5io4amfGxR2wDiFMR5EEDxdNDJEBMBnzlfaTiZmpJp
SqHPHmyj6eYggOioNHnBOoyBwKgqXDvqOubT9VAURi78DCywBoZimQARLHFrMaQW
P8rpdsYOgZj2PjKt2mlu0IhGri9o042WIztX0hXXuWO8UIGaGZGwH5w8euEML9FB
JYjNbbhfaGtEesbm86zsMJQUJN6PCT16BdZ+jyTItkB+kvdBRr7mlmNhOnjMs3/Y
BcUPopOHu948++n9EoOv0WGFYuF2fLwV/FJTExrkqhrV5OOA2muf9JbiYDK3c9A4
Bk0vdCOyb6YKNPYYu+IHTFDb9uBfn65Q5bGC1XPKoSVFXdHibS7RGvS9FkG+2min
Unkym+TMLyKyMvgifAhJ3gfQIvv1DCXo3AdzC8ySNdBer0gHk5RwHmXOQxNmKpF/
cM32u+HgAx4j9tDru+GYJ2VjVgyfvbf753fhaow0zrmO9cn9174ZofPRd5Vy/vzJ
HOK5O2Itwnzcr0BghfeRxigAqIFyuwRmOs6NrIvPgfSknkDC8kRyZiNQ3a4Oog9k
O0qP/V1nv2QomPZX/jKN5q/DA5oTXrFNNhpB7nRYOCGv6VJE+8o69xN/uMgXMQjz
nkr0qI+Wb50mr4oBCatMaaHU0WDO8vqgtm3BFMEvG6B66f/XkbZIGWJptXAFufr+
adZ0D2c74vpWHYXGJG64oQ2G0izWaoJRheYH81OOVPGdOKLGUHgadxXAoaklC4Rb
KiJ6dLFYr1wK2tFoCxL0Vn3pyg98oGBmhH8EFMDfEhmFMc3wCXKu++ILp3fbcDWn
6q73JYGbyVQ1UKp260hIZRhtY265aXcBeu0bxsShBKw/XUebvaWTmhKWqwODh2Ls
HPgpkT4R01Oks6k+3slTThErR62u4ySg+ivQdFwfxBIJTr3gBJZQB8hPbbgosN39
p2gvefuW/7inrXmQHa6qZ9fpvNgZK/qdOhOJbJVXl37Ew175PfbxlofdFcHjLx1E
4hQTO6vF+GTXSDGXoXIpBLY5o/hKa+/AsOn7OzhD73wRwIhCNabp7xjmb7r+csTb
lRFEMdaC+ncj3JxnAR/rtPoGqSMz18VMDhIpLd1f1vqVXBdH008pNC+ja1PbGOde
KSmv3RvvRewnMsgQs+87vggqtXFrRg1zHX4Kk3y3Q4gF4KavF8YkPB3HezKCe+Ok
cOs4aL3hbfnCN7QuDrTZ3u6xNyz7tQYgS77rLJ6QvtLBUawZclefOAIoXv1sMMIJ
0m7X+1cKb/ey4rdWgzfOkeH9m3vdrFMO0gyo1hPF1yCHp2m7KgXtvwJVnPfGRGEs
ABrNMG+lz+Du0VaRzKGr2mrKdNm572ySP9+VZyLNWUs9HItB+TTT8Ab8dY/kdL9/
dif7g2BzMWWhRCiy+Mfys1u6gLPg1N0JscewHK9pxe1nIqa89FGROzqQ35280EQm
U43vqM1IbFaT4IUoNi5r61pe/KF5byE5wcmtBBUvWz750y+Vqx1nEi8qgdqLFZFK
yKlTB+2aBQThciJZ5ahIUXs5oudZZXDojc1TVK9UfUq2ZhvUA/O6Ca7x2D8RIW6H
iA8BTYIYWqQGN56QIV9A7YloMRUVQ7drQYUC+1kpWQYCrWTgLBLUotyR114e1lUL
w8lzUyrVNdwh+b9bdBhGa8WWbwWG1p1zTqbo+XHvv1zXAbGGxce9MY2a7wsG8Dyp
McisDFh2fh3lkQfFEaW1P7dhDQB6J9dl6i9+3HUwXgEsdZwZDZdGUyvOccl3dEpu
lFM0Im86eBYqdGKVKkh9ZuYPfgYDjzSGZQhp2zrhc3wn28za8HBlMJtJyx7pq8nY
Txic+ZK1MsMccNXR5gA4mB/G0uYt0V9KGCyaOi9Kmvbnh2cc0GL/LHi45ffNKr/C
S8HqE0LCIZFZ1KwqreJvNoB1Q8Q4lxxpaQ59aF0mm3BrW1LPpqjt3OVqwlQdgu3t
Z1fP4AHVUT5KKL382peCL77jOJ9UuIqXjmQStVQW7/gO8diRUpiLjwGGLzSMVMh3
aRn3l5/j+hXaRWknlwX+IZbd2hU9Jg3AbekUnvgDQRmT4S4Z3veAqq1c+Jyf6va7
vU6vAByDxFksvly/DLD91DfaR22JqvX3XwNrn7TqmvhTPnV0qb7OHfGRPkl64jQu
D7SEtCmKp1PJydS/BZ0E7d72qCEmEjJj8EUealJ1RnAX+73WRA4z8husam89e5/X
fMauuuQwEpdxArFulEZ0D7qyjthYqMcUzDnXSZg7eHrdhhQz63ZZ2HwYVLhO+mlu
WdH+C5VWnlAN7b2j0psatpOnCBUu8yzSDphuSd0fjopWU2kuA+z9Ih+/VFVytonD
7afG/V0QsoWAXuhSx/gBn4lxRgK8P2VAkBTtATB+IDXvwWKaquYjOC9M8tgQPhtj
88EhTWhZKPcRwfomwWmOWdEENHEJMszcE4xeEQXEOsWp5jWtDuP07hQRdhvfHi2V
+rB1yKDk4iKkAPJX+BAkuFIna1fRaOdV+UJwrg1eRJ7h39rZSyQ7iuAJ5cGnybIw
FkUpb6/hBmvgzEDAIBcd4CXCFX7Vix4/pHvuKs2hoJiTi+JB6DafQP1LSNPYvTd0
afPK8xamgZmOhYptPV9xS8pQ4O8CVOe8j0mVqc/mrL9q7Tq5gv0cIm4I3P/nApGO
ad7IBg3mLYZPxQ7IwdKJk3lxMNJvKmXLZwQ4JojWEfN9urHTjAhIqjb68+9h1jln
QxoSF7RT05RJ4vQuvzbDdWglse+UcNU+6ZHiqwAJRMpdTYqkY9Ahs66cOLbrR5Rh
ltGmTMHe8HhksWEGKPJYvxX7MmhghELrzLtzgfba51Y=
`pragma protect end_protected
