// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:38 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
B4ou1g25cJYKp/7pFG/Xm8eZY1TEA3M0WILUmE/gIvWP6S+oBosA+OPueYgnZw90
9wrF1EE4TzBh66L6SeltLSRFLHkn6pS1uMuLBuwWdvM1XJKn8ihA1WFkpgxufHia
dI131COdFZg96yIiXw9r4OHcWiPpqDci0U9mB4ZtZRw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8272)
IhhCuuf+j6+E3nmCJQLjWUX1XUnDyzHC34pU+2dfIy+uD15rFd6jchk+HVaPDBE6
j9MYiIh85WL/WIEbH5eAikzEE41ZnwhmcyHME/F0aewrbW2xPseWcmqa29ZDGiSR
bNAuWgULTdATC/SQPaUWQQRUUBVMSagWzReLnKex2qQZTjy0xbMrJ+PghHcrUZo8
sdKmPo6TbnwJPmcSA73Q0py+arOBu6bTEfpYv7dwHyRpnWCsClpBxYYsSyn+pUCY
rV9bYsG1xqR1fh8YqRqGouJXKSFpMnKd3bsZKLqqtt9bi+hrcs+B0i5BOQaKgk3Y
NLftyVFRoyOAv85HlpzZY2KNWF8VhaMEmm52mo5DFo45bqpXpw/O9YIexqulwoGl
ZEaH0x/mMtot5DoQjdDbf/B9mCtVJ9WGMshdBpVYOmMM6n0jMl4J6P1iBulEDBX1
DcN0YFov3wo1VZ5hPUcNisNiMlv6hRzbM/NSvjJsTU4+HP5WjA6aF1V6RZYtFo/N
GC+eEQpPoyKxMlyVin3KhKHOaTuNrTLPg9uPicwT/00T77OrE2Hhtiil1XTi8crh
EoLB8qf2NxPi5Z9JgfisgMD+m/izNxqWfRQ3OmZqQ1ct1DnapVON9X0/StCtJsnj
4jZ1pc8ARrNfSPlH9MQhiZVC7DLR78G7WhiHx/mKWlAPOkXj3ocr/Av2mxp9Qkwv
Aw/vB7L2PzVMjpNER7PFB08X9xckS9anVyEmmuYQ62V/2oZJyqG1p2v+ENOrK486
id/xcNw8DgdZs9WOm7nEoYNR9A9zqha3hGKUEIFFyjKPnjuHMUMWjq18AO2xx3Sw
Uo0rw9iNXk9AU48OTLtb9vAfOTsbrfMlP7A59iliOioQifXj+29hp2/OdsRbkG41
wVMOnFgV6TNpiURNCajjygCez34ez0fhYAUZ/mFpSla7gbZTetkW0WQ+ibOb7xBi
myG3z0VvlW31BNomDhdpSD9JzW4uuNuaZ5on+AzVDUgkKIgpQABfQXecbphtwD4c
UUHi6vAJ+eqry8Nf5VavEsVaISRqe1E5g5rEYeFHCBhMKEbfhYZipR2gc51wf5xH
9ic3S1lkseRzYkAgB9rZrA2bfAl+gAQB4bGcN2sLDhnoWATosodG6wI6D0cTxZoX
wVUoA4Ub0tljn0lFI3SAP8cnTFCcq6dlVcPFuLnU09GUZanTlmDLovCv9JtoVLCT
N7ESOfQFdVsRLOi1oNrMHS9Nxb5fBCd7CYYmApzs4wFmji5ukdIuApkYWOdxU3aB
U9cKZAuw2M8G5k1/qSlm+fvs5MgQllbT6nyPYdH9WTaA7zMNYMHkDvDsaoL5Bpr1
3tXUt952P3eQf4EPUlI+5A3zKz+I5I3hWGz0fuWZXKG7zfe63h7uH4l0OWq2cY4m
0rka6ao9FuzDpB1JH4i8LNwVwlah/NgZImEubqfxgmR5aUh0Vnbhf8L8zmh6xsDS
cTnVJ329uTRinL9PiY6wAk+Uq0P5OpyRT5xcyvHjh5cU08CWbPG+2aHG4rnP60Su
0QxG+UkREW+xM5FcOJqFlTRKSVc3e1wCLM0jaibC0E2kh5js6FBj4DF80BCT5td/
xrYWUEDexM+pG8KUCe1HNzrLfPhQYz0kdMjJEvQjB/2tl8faUsRERFx/4j6ii+gC
WVD1aN+BNx9zKpooRbADN2/XI6AeLQYLoOcpEvi0JFU8iNg7NOj26sY0ho74U6ay
WPSlkpYXAnVZ0vKVwOm07faOMBHfP8CyUUW16iJ/dvKa7SARACN0nDxShN3PJKPR
s2YPMnUu29D/lYVKueiJxAKMCvegLrt47gG05bz82VX636mf5VzB5lHX8FdEiWCD
rKVOxzM5PG05RsPnaLBP5rel0z0tqvBYcdU3//SdR3EYUCxLiWIdjH5SN75JWHmL
tb9eWjnf5iYUEaUPvMPPEfA2Hb/HYVbNYQl0Geb9n0R+fO6YoPJg0q7VVx+zUgPn
g0g4iTsCM0Ld1KqH+kroIgbJEEzvAlJRjWJ0zRmKvQoIA3nqaoHvEOo1EYYs5wJz
mxZjRNvGapFNv2BWmtw7HkRkQXItVVmyLAuA1D8LG2FuNm4Oo8ty6QlPlI7U9a2m
gqs8sXFwvcLctq8VhHJHwXSccvd2xQGo4CvqcPxWLQL0TIJnfh7F8D5uzep93ed0
K/IgORYNGT/STvZdrhcckAlCAKhmk/I0K6BHC0jxLBInP3Ye7IM0CT2Se/dtyLjY
Tsxc3QxhXZSlK10nhujdWTFso0RGIv1GPSjpb+vs7JDUfOuUGM/JWVF6vNgcg20T
OFrkBDfZkPw2ecqjH7yJxWL4v80H4JQXH+5SifymmA1h/Ty6xGrDvRc+3Tbhxo6o
iErkZ5R89DvVFOM7mvw1/8ZD9WkdeD5H+Q8osdv37M3bbcZG1SB7pD5Qto00Qbhh
8lXhENM+vT/ZtQnqUOXkKgs2gZ12snz+AMUNVcjRtewLEYrmDTwwpFLyu6aRosoh
SBsD1vZ3ieB6HMsARVPSLYcIVOgGZSAYuoQty3YSGFTbPm9O0++cct0qh0KMQ4TR
KeZh76CVaKP0bvqsR0xiS9iCzq1x2FpQ3/RKAfqqz/JXGtCYwv/wy/VJLv6ONC4A
9RZm3u8FjVY56hsPkQljJmZgMZkb8/fhBWS8SOTKtTrbAryEc4A200lezuUQ1SmS
uYPpNf0qWF4EmDO4jBTNSVAnu7IjB9/8YfHBwqq0+i/LTOQIfeX08wJUz/7BGETY
vejEbD9qK9ESls2pSVnLhUxFOMvixJyKJ0vS5GYo3JdePoZLPq2h6sVavhZW7nO9
hf8W2a8NTBemHZ3TX1STLrlZd/dF++KxDf9W5FhRWPvJ9DuyEMO723N3yaCP99SV
aU/VJyZG9ET51M2mZeOUlH3HCDNjW5m7/MaY3txw1QsfevFBUb6QeAelC/Skfo9D
GO2X/VU9EhvQb3AvGYJEaIMi7g+15lv/nBgvu+gNyv1rogLbavCx5hL2t9gGqB8C
ce1NsXAG3RIiQ+8Dhk0O4F1IWQO/jmAq41Dyag/1Op8nh3lopqO7EwtsN5CjNIPS
2P4WNb0t6z8V+lZeUZIwd9Mv9NaQRrOLKNPyVddwl9LyK4VjhUXXr/Q+ZbDBgpdW
2RiqUsOAbP8w1+yu5y+7DjGZGyL329E3Gzo1dA7fdtwm7TIiIg052/wtgZBVgNzu
6Slk4bpHwItUYSZPx3Gygg85woXsMgb4636FqmCxjSgSYCxb66JlF7GQ0TYdFT4+
HGBI2WmFTRiLboLBfpEaWR/UdRQZW2dgogWPaCSnbYnpYNiTOVZThzzorozkP1YU
M4si3td7S/4ARVjX6DBZGO/xVTVvzKPpBGsZDq6ZDQPgQFJjiigt4GOOm9xA8Nbs
gkM0hO0WAoF7sgPdsGpew15A0YzIQm1RONM4Wi2N0XKZxVbL1cUl9AdFsTBRhniV
+G0PnO/zJSvv1Qars8xyphxdN4UitelcUZnKNHON9hK9QWbUckbuAq+JsnF8rWLC
I0UGkd4pOv1CiFhmlLs2WxJnH9Ao/1lql8aJOVjd6PKGzxvLtMun07Ns4COeoLV3
zxLcGuOa+5qUtJVtC758jm/N8pqi3YIOGWizBTWa4Xg72ok2LItLSaNBsEJh8H6p
DluTsOxHe+SUQDDLc9U1fWITn49DETbJf0zxK3PqliDh6iN/+LmZCMtFLFdWtIxA
qO90boULD2SD4hkPKqMCvJSvtUOmDR5iKjoEkkYxkHt0EnYw1mj3whBFlyFSlVYe
zoH9PYX4i3SHXQ0GMMLKVwfFg/MU/cbwbuqipvGEr5Ixn2fT3FyetqFQx4OHtZNH
8lHYWtMfk9mpAuCnsh3+Ea3qnj5HF1NywTE8SUii815SOG2dl507ruItlhpW33sA
pX0NuQdGiE+Sp+n/7f99s8istvoT4V/q6uiyW0d+wgt5/arprZnZwYUpv2fiTDrm
Qvae/63s+a/Mt1Iiz+FE7FqPpGPf4JQRZao0nsAVeDUnsmS1puGCL4mSgHb/De3/
WqcsLKLqs7xEheP25B/gJwfXqsOQKIJchxVqRV+fHgSZcFcHvqROaB9VTemgVdw0
c7adR++X8afJCnxspmMd2C4LUhXPxzPTGIzbnRMJulsvGahgh/xBKEcvADf3Ury2
WC4AbZhfG+fx4Lw8K9mgJS50Giw/773ew80XsSYf2X0RhSv8hVB28en6vN8Qwl++
fpG6TcglFqRh5W2eipoYG6OcpiO+3P1JLS/h3hnzWljDr1TzhId+BHbhL55RsWSe
Au+Q6Il53bzEu3/g6ELo199ydnovVcMw7cIkYPfst8XMAe0lQK3nFs8D5bGEKk8l
7gNSa5FmmIo/3p4VYNw2x+XNRxmmtJMXxEJU2b1Q3cl0nuWhRhH5+DoUHvV1uBSb
1gLm6obvARB+5WVeNBch+dzY0C5xioccCSpFBnyER1PPFECsXA7jvXrByR/l7yKG
fAf12MgZWINSSY5l/9OF+V6eRFHZX0USGaZAko4SdgPdK9airPtpne3mTRCPQ5mg
BMvVOAYvtxCYbOZ16QknXTuTA63Ztzv3baeWutncADR2RAmHO45OyFQQfKDCsj5M
rp570sF4SRMu2h8ULL9iXvAcw2hi25VdNaDu9Ne7siuAE6zf+6nV0FPkyAubu5+K
gf5B+iOy29vn7ugMOF2S2Dzo3ar9hoySM8FYMksg/ZYNGP1r0Q1SO52QjH0dAOLT
UDJ89I+2EDgoorRMlpZvgullyrmUfwq3YoHlf/52/cQ9XBEDyL/ucPiclzuD4vaU
zeXEMmRrRBF4PA26tG/umawI8l6OG22I6M7wkIOemHzpd/zPXpV123bTiHD5L/5y
2e+ihA2ZEs/jDVPP4gAmAXICbLTanooLRLCdbpiGBNrNiwrYJhQWS/uYqRgDsCVA
17SPOc/qeJwWzB43Aj325TIt1bDIKfAQuRwM+999XjtDb2Us11paewrwvXZQ50HG
kYI1U6QK/qGpBgZthKp+0fFZaa8haFywxx+wwqARTweTVSM0xC9BVtbqnOh0zrpg
QbAY0HRa+doopNxHlv4LOMyJbQDNeOvV58LEV+n9/83kQOVhlder8FZNugth6KmR
UGOo+Bbsaqqr/qlsgP22w7uKgjXhmuWvjfYyp5gXHHUXndiZ48FIK20r5ARhIwQC
UiFZ+xY/edetfUD177tKar5JdZzDiBkjsTlEtaUrE3qSNPaT3nQmf68CuFbJHZRy
MYNZABXC//cW2FkaReVGUuhx0AWHBPENrnRS9S0ITxwMpILd2mXLvDI+k46VlsUo
SY/BtDJDkHV3tHm2uRsFT0bXX8huZX3K2fnDA+qg6wU5zRkxbUawZfqIqguFGSEn
nedG5yyhHdWrEoPOtbnayE63NOfxLADSj+Wk9lVtsvcK9Wrgib9rVWMJO7kSxwVt
PR4pM1JZ+9vEbbq+KNLqdICGHGQVhzHuh2NqVK/mQ2fpVyxi5n15zIab5TiGIW6D
aaRFVxH27hOd7JqwyLPO1lUY05liKeefuI+NuJvg6/PUrxVdu8eGtAaw8xQCuvYR
kcZ1Q/jAB7v83RkML2uWFCVLpw3DLQVJK96CKUCPTOCCFmCdZf3Q6elJ4LX+SXru
xLrCyrNWQxjP29CGmfIuAj3ZUwSHcKV63SCDxWlZPTTr/u08G5M8A2w9VuF7R0vA
tTbAKEbLWnIukeOe6KcnDsRNi1T6dGJHGUoV7aQhP6UtVEBrLBGfDwxgc3BR/ow3
XTqCBPA/3i4/D6uqrlwvLUrgdH7/qkqOcUCWGsG+7rGpd8kA1gkksbExYDPRZWgz
3dmMQBNUMILva96hoxrHJ6YKIA6XSuqOJ4QtcrlxXzdpj6OBlCrR9HIr93a6baQE
W2DeSOwXBZwaGwxJchmQnemtJN53lu2HY7YObWEMs4yTmwAEkaMbbgHDC23L7B1u
EhheMqC6sBQ9d65v4m5Dj4BiY/skAQMKO2WA7XlKzlJjg0QuTifz50aY60tsNXYP
TJHEJteOhikpAxwr21CLR/bml+WhwORNJ154rQx1nLMFTNDTXADBBzsbuq4vdH3m
D7hcyjw4173Fg3KK/R4JGtLjUaFoJomITGJc+4ZFa872u6Lp/NN3lOM2ri616NE3
55W8KEYr4nZ6VHCDavwORO2/ss/6n/BI+1911fHaebaV+JWk/Gl7T7UVdTNRIVe6
lc97yDCmC2Jg9NePEmEMqZlwHFuMzNisAAkD9jLAHxWbMGHU+MmfhXisivfMI4lW
Ihd3eT55FVU3/DVfqk+DyBfzKmGm2dyF5N4wga1ys0GMU/5miMCS+a5/wenfd/DY
ySvnphWAiquQsHT5zwcTQxlAFgVhZj1g9qZRJrIJqmY34IjesEr1DmGIs3r+azYV
GRNkXOmDP7n32YSc7bVIgQ7qVUc+EJDAf4YmMyPlmNa7E/7lbXgUqa7KO70lNTrH
yZoyLfEzGZ6562090j1cS5zGS++FiiPCzc//NJTg4j6aB9z64rPlWj3Afr3SvMYj
8N1hpD48kcnSpuOqNxWaygyWypi86UXj2owKG69o3G3ncWd5Gkag+idnV4cwqkYv
AGPPS0vS0IWh9rvQHo1pHN6JKranbBLGVpL55tTCm53NeBnL3Qo9JN8OJrnknhtM
7F5hyIPXftQU4/rtN7+87rfeLzjezYYM/vcJdJz+UQOmpTv/ls4h4wqn05rQhu3H
icv1WbCLqYd/Q9f6zgT5cfebbxtuFj8/s90v/e8h+JFadJaYYC3ajJgAQ4XKVCI+
oPeOn3S0XIphyDkg0RIQXGTtqa/An4hUmL2zAtMaDqz8j5GDkxsUoQxux69uW+qG
RJ9zXkQE8fSg3TGhe8BKTTNVPa9FQH2HNfw1ldjGrcT6dRgWEBb6P/h8e1QM7yCQ
bfhnZAcAcvhkGt2qjj7YE6+pXhxe6wnSoKa5xt0PvbiMCb3WC24w0wcCql6caOHj
ZVZA+eg+7eDb5muv5IO6JnzMW/8PECaG615yggyYKaTKTZuWaJNuNr4T0/z7q5+6
0Q4zHTCNNNbEDPpDp71AIkXr0in/o17Z31zBYukpRsINYvRza6/5tWv+HITAd30r
Le9FNj6QahSptbIzII3QTQy7sJewGxwQ+uiHegIItu6jci7cqx0/ILX3RTbIdshP
ncoXXgM0Btr2VFedpAvhYa20a3fDjCnhDxivTieBwX5AbsuLS1XZnUVSdsfqlovF
N5EcAeAkZ1lo9uoV1pbSEfFRmYoqm61PLTDGCEapT6Mup4cXUVu3OKD1NgTWij2B
mmoF4g3CELWxoUOtclp3AfbNnXO+DZefhrehjg0Zu5q9oDBYfJd5ybYBTwMRAbyY
h2eTuTIoYR3mB5afiRfvG94xAPZw5DlCZfV/qyisbj2v+fh2pxInWR+byeEVn7AU
MG7+c8V2PiFFZ5TcvcX4xhdtyjpdTenwcqZ2os9jj+5N1WJCX09c2EvClw5IE8BO
FmUYpMsXRvoBjSTUiPKRF27aN7gknL5cbPojWLvXaZ6q5scaLjPcRzJgbiE+ZC06
ofZmlEJ7ImF3iiO/nXUV4AdcgE67ixO/6NrnXZkOZZCK7MTGsCJcRzAfD2mf8wla
sWdNNBVS1ijqelJSpAg7prUwoXDAX4nFscARXe0hjQZVS2AcwdRA81SeeJ41rN0Y
I/bHJg/gkg6sjY5Clpf8a4bJR+YCFLW/l9aK3/xHa6WlH7pk2kUFQuk/M4pgZ9eR
QlaGirKOd9OFW52c8WlKAtO+kjdRbmHvPdcauDZWsRf3fe6ozkKfwO7x35ePPNIF
Xg2w5dYtru8GcKHyx6vGPKebe7O7Smpz2OMYvtJOrm7CJ76IJCKpYfq9NIBNkOXS
UksY2lF6HAFIy56ac0aOaD+VxnVNI/wTOe3Z++d2+j45sHSvmwVKPZAdBm/AD6AR
+vnQ+yoTpw5fr9IrjtEUh63cZoDf7NNI2xaDkmG04pQLK/VAA2dvlCOQXI1rMDlK
qx6QaqcyWAPZu9yirr5oXFJEeA2GjX7Hi+7iTeQBJST2NkDdJ63A+UuAUm2Nl9aK
dg98kH8hcaVuqPitn/JzkkVADcxU8+dR5v59nEEJZHI+K4eC1eMgQj8zYqeTXxa6
/CNQqS8hSjbVv/mcsyRbQScZgdYhgenoCmkwThtOQUUa8pFgtdulcsN77bMxywKE
za2U8FQSyz0pRTOAcKYSQejGT8BQBP9p+W9VBK2o6t6TGLpkyUzpxLhLR8IFZ9Gj
0iVqKmNogDsd5CUm/oWvvocknmCFBCg8Ex/DaClu/sNKeehVHqExoJVug12lHTs6
Kz9avBY654bLacd0MHHpoXfn9gZIutqr5aHUWdx0hs2fq8FqWRZ+zVSARLWDBG2Z
dFXqgH80fz7uoGIOVAXvMDP9QrQnGQHPJWn+rPOOoXZ43J1SaxlCVGYuQz3+7h4I
1S6gGiOvLsCaHJqwZdTCa8qHhzXaEGie63xjKgzKgxlpUpFlFWIYYvdF9f6duh6l
Vwzv/lB77NcIVsx8MO7xCSwAH9+z7yXpTOQauUfjqrCu1qft5ENkjOXNj8Gk4vG+
cLb47AjOdrtatj3D9iqojzRjQ9C5vxrtPeMSvfmbv9fm7U814xW7kYPXPPrLvyui
m1hr7oLisVmGwrrqadCALEr22hlPmxXq2bGcLnQ+yuMfBtm5VGhLG32SWe5EHNeJ
7uStokIAjHO1tL321jKgHvUNfkZ3cvBIEYGv+mW2iLm9+Ox41UiJAgFJFz7DWDlg
xi0h4THE/C7i2UWdrIhrbNqn3bfnxedUEUrKyWvTH0yc2gf72vag3UbPaxjtuwl/
T2US32hQn3PWzG7TPErcMfOKGUpGRlIfpFbrNEXnA5LGlSYD3SlJuoNNhWAOGmwT
E2dbaPdCsMHf+fgMp3MT+zv6COrpZuKa2ds8s3hIBWcW5+JwR7DNMzYQZ+YcwYAq
ECD/Pa29UR5OfqlVGfELrKq5pVAZSJQ7CLF6+KDe9ejIMVmLl0EBQ8YSIrLDlRcn
c4ltVTrOUHVB2oZ+rSmXRuEt3uoHBoUUGsJl3u1UXWfEnoqNob5XAZuc5uCSTOYX
gbY9ijPh3ZLYjLJoCN3bbIONmGPCkKyBJKwqgRarsEyjmb5QflOAd3VNFGqtWBi3
mzIeAFJlezZmFzwOgqiR5trfWHdApaD2d9HsBU75SPDLiXUFL3Z2pFy/lfzCrall
LvxF6qzn+O+IDkHJg4ihZpcKYNw7+b1QAfZYGlT3A2Hok6uM5Wgl4W9PFIyaVS3Z
l+PBj0uWSCtISBTXkG8GwYzCGEUgkZ6R/u1QH4dGzmA0ZpgxTUafAId3UtxjYDPq
WHwdz+ZZCU39Pot01QxKW/upipLwMDHcsKOd/SHV4ICL2xzK26E1E+N9wL41nsdu
KBEGgurJo4ASO/QQqxHAw9t6EK8gD9BAqV78nv1EKAhnLWX8TTiSOe0ZBKSSNWQf
cWdQaMAfOGsGNH6JaEJCZvCS6Sk2dP2W6FljgPnmHf6YRR9O8B45EgF1VY31AP7t
mDDPmgkE/RG9nB9eEfMV9YYPxnS4tnk96PgCcqqJ9qtwzoh8gyh0i0xiDzxG7NB3
WoPepR40KC50CyMZ4CQw2tGnY71JF0tx7UNPVd/apgDUEMObt1bK8mlWcsv8aFV3
i0twJf6SDv+YD9WVywqFHV9yh9X03RlWDlOlkxN7Qp3MlFEyUH/dKtyoeaASLq4X
hjo3tCyIE1Yl2LQSya7RAuZo46k2nd/DFOJ5Q6OKgLaQr1fMHMu4VqPuVTdpUHtc
S1clGwBd8jwpKHSE8qziIYG65NnvxS43BVjUFoi1Iqa//eBfot6ppIP4GTGw9vvh
pmKrMnHtFU3yvA0jDnIG10XNkwJtFldq+3yzMBFkgVBI3zK+TsXgjYfum9YR5uaZ
a8b6qACMmqe4q0tMOG4pDkAPVIQZdTuK5F7pwcx8ArsEFCHGcmqaj9YWBRnLPS+Z
kZT6TDKqydE3WGTgXN+gREOJRNTLhL9la/8uUUFEv5VjqW5wVNRhf0TfYfXRfQb5
w3Bkg/SUiZ0cXCqKHr8rVgtsuxgf3Fs30QQrmZj409ntYUUr51eaBaGtm5rY8U9w
2Z9iXw9Z18Trgljobeh97oVfybyrUYasF2d0c/m3GswlQeqjdAgB+XlktPZXqdYL
SO+nUcF7r1yum95Kf5aUWB5duP45Padkbmno4vCsgGh8eGJQav6XV6NAswL9tncq
0Ayii3MPO1V378EuzwJ4HeORC4S4NB0IBkt4wUAdAxseN7bmPbwCnVT71zIZW0zk
0Dct0RwKb8EdJhoAKEkY59uGkopPbrAFCplteEVOAnIJMNEN5PKiI0uLi3oVJoHF
w0emhXyuE7I1IuKj+H1SqnkbO4Y53tJwwxgyOpoM4JVWtCjuA2EpbbMnodLFbRvI
W780FCmGshkbaenQrEPR3GZz3NmKK2GU/EZjAJAWbn8UAzfqf1U9GrkYvQ95ETRW
3GXUWbwNB2WnrM39Dtp4zAfiwQ8Kotl5Z36BtV9OAHbxl93yGvckAAvQeaEHrv9a
5V5/BJCKPcxF0/9E758QRSd4L/ZVNOrf764fTMUYIiRTAsX55PPWa29dQ/F06eHo
4+DgNCAX5KiCd1SkDnrWWFApld6LMjylDYcq6Wsy3GsNsI5tOVboSqMdflJF/uoD
IPwtVegzERJ8oJT4D8Q9QwpK3o6c3pORMs89er0dA3jA0HYGr53RmVM6/x19n5ck
2ESHMmFSMiM1DhvvIjr2USbcrb+DCxVhgRO0C5epf0PBWWzyrzsxEKQfgsDsBqxj
deD61bBil4Oy0ewwCXZj+vpxRohPIaPL4OQ4wG+preO41kqKe8Iqxot29jmfPGQS
XTlYQzLHbPEiJSGzvl8vLhNindtQMNeA++/sktkbOH++2MCsTPPjyBbHZRt0NazP
fuqxP49oJMXMgg2bbkkz9pBTlFGFQ06j8BnSIpAAJiNM6hkovXR0awilvhts7X0x
MP5OyPCS6ZQoGhpNfrFodg==
`pragma protect end_protected
