// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:46 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oLorV2az7yzwRXA2hEWBGDJQmHSmZwAbb3bAqe/Me+N8oUETexVjDr3IsAn+QRnb
EkFB24Vqvq8G/H2i9C6bWjxgxsrHLLTUtlA4NHTujiDO3afkEaic8q1Yp/Rz9KnR
9Dx7IrX8hEKmj0ppIXW4yQY2nDY2GeoalWHb2EOTPCM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22384)
PjkKChObUZXEZWaiTkGI4qtHh6m+vAAW6nwmqh2dSjX89k41hRJpMe/jdqmN9pYc
K28joX3/MeivMjFNG4ymoWyNMkkTtfVpAeHeRWL1//JuswGbj/lvJwn4gkVgfJC6
CW2J7Daj7SM76xQiiTFZm6BTQ89imA3xLgCJMKGH6pc0McYrIJe9ukot4R+jpNVi
hrYOAEpeYcGAAS0jWxoTZ7V5ik5cf4BLj9cf9V6xDUxnEYzfS+rl+6XF5F5X4Rz3
m8t0g6OrmjcoAUyDE7bWJO9hb8dctZ2CBwg9A2VGi1xxI1J2XumZUOucvTsTuFZZ
p/Dcqaf+XnvWtTr22gG4LmSvQk8nYUCZyLyPjkxt1htPQSqjuFkzO6HiF7FOe5gS
taqH1tqKpQpy6RI8oEGsql+mKVPmsnXeDaNf91KsEO7u03Vh/3HigD+zx/7NI6If
8e6i1wIHssrB/i9knmADaMT5eZR250KoZe+qamQSivHJDnOgem9IpilPsAZhVKqy
ZXA5ta5IdxBCc6qvKHp9170SjWQN1bKYt6TVO/4DpJFJAOiBgAd73Qi9q7VUE/4X
uCGYEG2R8q62jK+Ikt5HS0V48NhfO7N+vfff5GjIrJ5VolKCPq7EZ3YLKakrVbh9
S4IyG7viUxlI1gEaSgnIFkrL1Uaguuu45ePygvYsRkqJgDKQuNdesiiDPe1dJxuQ
yuZQEl65toFf6Xq6yUMmL+FwTfxgbIdydnIbz3LrJsXyhiKkFHf8NFGvDzSWMTd9
i9cZjJpWyhJOL3lLWRInvqRUvNRkpqaarv6qv8Ar/4OxpswbQxe0+65Fj9i4be7W
Ncr1at1h/kRVaSVVUD4HcKi2Yla9SfSMTCgW0aX1FNuefQN7NfOysnqSiUWwGuPY
d2pKwJAN6nXSpajq5/qyjDfSQ40k6Kb4HjJo1BWEDLz039ENGyXghhWaAZt8L/R4
0n63sjkor18X/Ph5pugAUcQ+pfJXIlh4FPvo5b/T6/BexXcBXVaLhXuKNWD6kmmz
bSaAMVMGdZbD+7HaU87Y2xIrRgo5mKUUrrFxPxlsNQjoV5pdgczAWOGZghG+E6mg
KviggBaLtgs2jsJyoLBV300UuTwoHKkqzcINLXZGiB9abZYVDZ+Ki4d2G3IOlY2e
hZcjtawPYb5nBf+kEhfvdhM/dSFeb8ACJMi0B3uqq/IxYTBtkLlQkKIxITtf96Hs
MASyrSk0wNWUVSNEJ6+R5aDt1UGk3vtqfuCPOd3+VE7TixCMv5XcR+IDNmFdTqLP
jnws7Rvz20tVnveHTId1CKRW7ESzH01yuninuSRE9fzOTVQfS0Cr+on3/hwYDvsA
J87HIaMfW89eOTP4yv/LEC2doCy1ETuBG8lER7ME1ro9bfbtdUyhWWXHTLymqvPm
NOg/s/N3ALLdsyfZXuUBzkJLcjhd2bFl5UTAlPW8E+PqZxu2Np3h1MaPo1DPayGf
WWYogzUrtSAzDxLCVXch0oxEo/R4/4xLyNUWJZpmUngfYNpKv0wWs2w6s8d9ywM7
1HHJGHvPozPd7nGpz9zjakNJmm4oX4y6xmqqwEfFxcZTO0SsuGQ3ZXFkU9dXlBMR
PmRmoamqferRfLa6BW7ODfxhrpLqKBt2LzMMPTVCVy9Q2tTdRFRcJK+at6qfHv+a
kibQcGGFTHWF2RiYO0GqI2h6fMf6U1XlQU0io/xWf58V0jh0dOuR2oTZQbKJyyvS
En3MS6x1Sj5Qj6HWSGkbCRqqdEg8P+LOXhtRi0Im462Mq1yjphZ9rWlrD5xq39P+
b/I0ws6y/DfPHcfzqoDiEkZDfJEo5rgGDq/FSkUKzpA8NHCUngV2KNpb3CTd75Te
qCV0T/9wggYWNk0JniE7dtVDTwBc5inc3wlJg61qP2HaFErhmU4eg0zWa8JagAuT
hLelPRtbZG92V62cXnmahqe+cetW5RjbgjyIKGG3xCvRP9G+CevcoYOyl3BZ56Ke
s28L2Cj+B6y9NcIvtwrm7onUssWwQUmkR+a9mL2vAK+phwY9C2LOgrfM8p0ogETg
nFVTlRs3CG2vUtgZxFCiDLHR39nwwERkz4q1CGjH+iokqUWndAwf+1D9ul4DS+y6
/LjdyJyD3G+3weAdHQL/HNUkl1pLRLMjfdtmyJoXYHY6hqplWnvlvKb4uz3DCYgh
5bYeyC3UAxP/lF32pW4TmhV1+naGinKSIZCjN8+v0/kTRzQJQ6NbgQxQ23oC/qV4
/Ov/1s9vmC0GhIfLvVW4ttazAJoSYMnWZxEZbmb3BXE6QpK/SiqRNoMe65Om+yXO
MoHwAhBeaMJvrxgUc9UVSEhxuCCsC6osS9rI+7W2ALOPRMClzthzc61wuagblD70
+KjrmLcXTFQ4/isCLwPdL+dvt7ZlRVDjdC5aRW5aGPspacYMo9m1GWl03vFDJXla
LjrW/UEI+OOfq2D6U1W487CItje6M6z1jVcadv/v/NoogJyQL/79e1+nw6NPBwDd
84TAUjJvkTzpUWNcqVD7Ci8wb9Eq/FMpnBaeDqGFdDz2mJkiAUv/hss/08nQgF2C
k+I0NJ+LIU8JlmhHaR8kEd27yVE4c2oO4RmMmCB9slrikvAxf318MmQgDN/eRiT2
RjaZLbm4w88VO03hjqsAenB/Gc57V6kz6TIIoHk9Lz+nrGDPG4s6+JgsGDxcVBjI
IV88cMsMoK4PY/qTnr0nAwoUksrGsYtv0L4RLu70hWEmFWb55NTF2hfeVejGnc9v
g9FzRBbr4RDiO8hcEsJJGVFfPEEMxgDgGyeSQF9/JC7Up23FCCBRGghVo4eI5yp5
sG1Ozse6M8rFQEpn1mXFADEtiL60wAEtWIh2A3HOz5+jPpbsxbrj/Gy72DKbEAC3
fVLJr0dVKjvEqYwOzMAJf85XMACmUJ0Iwp+xMrhaemOqtGDQlEjWOVWHQ3I3iF2K
HAJFTj3zC6kEMiVGaUFqZLg2+ygPa6jOHZpvPcshmd8uH8qGz7O2pbQ5jA4nw134
XJAsCW/G0UQAoJscL/HAX4ZrZbntwXWrtrnZd8Zj4GAjGL8eC2Ry12LpkrAbOWGy
A8Vyz8eredCvqCPLB0kwwoYwrxF1Dhsdo0/QfXJKyc8pOZWgM0b0/f/rs+pKMDmE
Xrv3AN2Zq8T15JFqkQabUlqS10mfNI0/rHy8L7iRL2jk/xycpEGZLcLG/S6DI/4N
EFtPAnEPIJvW6EHu53tzcbX3Qd+5OZDtgeCFtg/4n70ELJjefqcJz+/R83Droap5
2czb0yoKmmhQtKBbjuBuSKevmKuZ/3cYALSme4CpE3qBsI+7kwZL6enexG/do7K3
9gnHlSazkqaR4lDD4rmDTDbH++uKxVM3q2aSXL8nt8la0Qw573uQuag7jSf002Zt
vgA1EHvhvOSlE+qX7AKPzxHNhtWZIq2FH72HYDfeJmsE6qmBeoJDLFeOUcZpNjWw
lCFLllvvHER4CDJfn0eKWkZSQSL3xdD+rTpmOOB54cc3RTZPsO+U+deeaQoAOCnM
zWf2vvg9AuZjYFYn1iRFx08eZQ/P0Oxh8FbOXQ/fg61D0pa1+zh69rMGc0/4B91S
qU0Ro3OctUXsu5qdsg2nIqdd9L/TVpbiJQgExVIz4T7btmGJvuydwNOWK/BVuAsZ
CbE2gNQ8Bt/moHk9onnW0RTsE4vH3jzV/SJnDjYw3tNOQzxr1qX8y4W0pPmUlLrt
0r0mjCLlw8J8I7G/FYD/edusaIfYGTMA2s6VKCMuViP2FUJ7Iyt9RgFa/uoUICEy
Qjv4Gfduw4D5mBbnklbPieyXPtRC8v+hd10HTo/J30IeOxsI/Wn7Hwn6wnf0hF5C
2cogqzz2/IqIzY2JYrN3WsiQWjEMEG9qlFx4Pd9u7GuPs/ImBvHsygVv0lfygKRW
yDMIbjoxFcTaQngGF31/Woi9B6mr075Fvmb7TEk4Wk2BQFF3SFrFyHEUdfB2ENi0
5IWqoOZYtgb82McXOWfWuH6gXUflwrzOEASRIptxEuxrOxGiTDcdCkssE2BTF8O3
Zcz7m/Tpz9pA5FrEDVQlYQI+WFnjQdSLcnzEe9EY3nMvYlo25p45+QO31ob1uW+f
iNkoLsTfkf3dQPs1Y9IbxQKuyjDCh4po5F1+cwoz04m04X7PjD4GWcUfaH4buV1M
BSwAG++1yKQyYbuQnAkB188Hyz82wwoN7AAm0wKDuF/90gN16ROFpQQbFoK6ZOM+
w9/fpGsErD4m6Ni1uM8YI7BUH2Wg7HtMgUBzKZsS3kSXeNiJX7WmaAsQACASJKid
1czPNISQVMXZldB06hZ449Yi04Sk/U7feDHsJk1TrhBXBsQ8LT5oXWtzTQ5vGBnY
Tow6Bg/SsaA38Anl/4O2gIJ5ZH0cW4SYx85nI85ulFPvfzrZhyjLiUKMnVZaNzj6
vLJaXX51U+qUHZpJiPyXwYQ7ni2wz6FEm6pTmSFTjr0H3iJKQrboACUxiK6wVuSp
3CTwCX5wsIs88bISuDaSWoZFBxNb42VCbUbH7GWTLENRcS8LqjWcWe3PVNgC28nB
M0gIfEki1L4z5EGcuqRCN5HJnapwRuSCQ/YGT36WwtBOydi82NlQMQysml3eZpIL
BLotibByDTsqNWLc2sJlc4GdQEJEx1/h3LqhichDFh+qOKvmuqHdGnVDz5JVtHHu
dz0iTtvgFEapUaj3cCT6z3Z61GGlr7BV2kez3GFIYrBoz+vfIm5TBYVx3HdIvBAf
6Fudn/rq72e+bymHnsbRNwnu+2EclR78RlOgpQZE5e0dCkCRJLLSVgyHYiXE2U75
Kq5vYUyfNS0O7wE23sG9JJpyAyhDlykn4rl4qBDd2FXR8tSDB8QQ7SLgoHG1Ifk8
bo1S6Gq7/ru//cOBQPtWmBpzvKfEqyaMtDPgozc6UDhwG7klRvjRIZRA8KX9PQuI
TL9OQT0Wqp0Z7g53uWzOgXhaicL3Nxo+sX95U+STfiJR34GPIzwuKmQ/6Sy6jNfH
+24t9TAtjW0abHMRjfoixQyHDVevfVPlmwVgsdjbBV9RKry4FYCMJl0pwgNBAa6A
rSbT8mBFJadfNRJ4Z/et08CmYD2xGzdFaH1DmUuB4mQZIKRQ5c6tTEb7ExdG2wXx
tY6/wjNrO/IjxQzRue/d4H73lPiyL5acg0b3QUEhrjfM4B2wHjxv+eSyLY+IZPBs
kHojbOTBvtYviwvSRa3ghJGm9NuboD7bvSxokDrAlhMLzn8ceju4lmCee4KRQUO0
/6C1XDVeoFPCW/RSHRi+2qo3HmwqAdjIMVG7oYeLzMmTTRD4BoIFpJWyBclzjeI1
ti2anhOZwmF6VTpyfBQpk+p5kINuZRYERZ3b8f1ROQjSUNXCD/TmPrkFtgxxQHmd
iMst8H1ett8Z0f05ln307K9cmP89V2wMMcHlTlUbwhOshJk9vXUcpnWdAhWwujeg
AquX7vRLVe9Up9qTrPF9qmiQwpDAfoBbmXZcIMXOR7TUbMlV6k8SkOgXuEqktZ1l
WC5LKmXQ1telLf5T6Ds2Usyelcf0NQNrB8MCqG4zq17IFyHGVrC14DqWPlY5NyVw
nE7aPWntqC0lJq9dUYXTmyixew3mP0PbKV1MTlfDRBsAATqjt+fwdNN9WxVcGt2N
mi5T9Y+JktlMc+yw5UBSKTQRTdOrtU/QHQ6eF1rHiIl7sserG0AWfZokuF9FjKrB
JASuB/R42JOIA1XNn+BPwHd4hKZX9stOmaoF4LmuMcD64yi8eZ5oRNGjEzX3wywz
aDVS1TUh8Hlh1jUiPdbppxnTC/v5kGRcVn+owgztZ12u8FBkRRVOZqMedMPv98B7
DQeelAe7kvN66NaP9RPJNofyT5G33PXHGY7sEwBGGIXu5xnRQt9hOEIqVrsQmOMx
x0Ze7j6l5UsYzdo/S9jKmkmm/G+QSN911Q+ntCltJmLFq0pn4d8JugVBlF6RnfNa
UsHLV+DSEphkCwIuUobel47UuX/jaB5AWtm8BRHyS5Eybb9bx4UUigabPA+LCmqO
8mCOhD3yR/HZ6VpHzOLEgJ5sbgTixWgjtqAvBTJUccERFnRVjSnFAxcgtz7zxFpT
RiqRbjF27gN3xVXwbx3+7c83DMmKkOZn1aWDdpUcYMAwPoslWZAYCucb39hAyC2m
CejncfTWrckHk9B1F8ewAui0lTmv5hsoo1x7en4f+nT2MCTX4O8EIrQ+Zlre/8QW
JcQ/4p8AuBTv2rWFFd+KLXyRe8LlB/3Q12JmYgiCx+UPJtu8rTAdq72UQx02va9U
hq1yA9SOSw8C0osFfbTla07HsGkbSP+MHO6034/ZW9OwuXO60bf1rIC3W6xLpLUm
EiLs9S1OpCfj7FdETj1iE+9yDXO1jZ4F8XiIUezHDWpMOus90Z/wlQT6OiRJNyD2
ByFD6vplYMe9QJPe+6MkDjMqqJcO+uMLvca2+1KqFRt2z9MxHZnlcs64cEbXOkiY
C57SN5WtPI9LRKarVUo+NttMWWDV5e7AClnI+qjdeGavhCEE2/thtuRA7nA+9xSI
rnwAtWcRtQjFqC4ZWDkDip21CyXf7Y5LjDu5ZjGSWA4LZTGpkYePCKsJskq3kAjz
UwKyGZONiKOvWvU7Kg4AT+4X20C04uZEeFH+vpMbBzytQx7hl1osQN41mMho/4/U
Oe+D7CuoUUL3j42Hcl8unRE2trCy8m1nVTh1+YEt8AkGwFLnA3e+efeAaCOxeAKk
H/W9UiubTwfNx858XDlK1OsSn7nmZoeqkap0MujFoHXMUcBk8IpWlAg29DMWuFqh
9mE9HTdD3f7d3C64GYjRUnWSnkVO5OO5BkqThppOVdYO69a3Fd3B+W1phn8QsXb/
WfIJEKD3mqf+oIyr+dFp0uIvrpLoacygXFfoCcrsyw6PImNy+/QnDXPIjstgrI7h
P0Po659Qe5ctrps+VhJZiJ3M8PciORS2cHwI2IySgzk7Z+iJVWOJyaeVib4aGyee
lMSL+tJQnlXcU3wn0rtJi8z+lPa/I9aUtjkmxURXVk+kJlUhB9ma+u6YyVVELoLs
4nxhm/Y1a2DaWRbMPH6RADh43OcEbF5/yhBQcf7MW/jFaFQ93ZKArMTB8xKvwUwv
dwVucp3uOwZwK29nfNHvTjnk8wDLQvqjzjnqBsq8ezGJDHycVm0yeWPhgGhDQEfK
O/KaIeZ66Icd8TEgZVjmJU5ukPzpzUIh5ezoXyNvTBQxpU9AB9Dm/QAve81QkX7W
dO6GCaNB8NZj8166wm3OkJpj/ra3vS7PJBVi6Q4oWnTMzqK+ingpfW+GG/pl+FQW
cG8qB04ZbzC9NaiaSE+xWX2jaltzNIthey9+FyXC6k9OqEvU/NEXcHjurAgL3ncJ
kR3SIJQI5gx5AzcvHdra62W/XiiZMDokRUGyinOksFD6F2hFvL/7JUdzbwiGKKIW
ws1AhGhSXoR4ZB1nydgAZELGCz/NwF0ngw/Kk2OYkyDUHYqXkc+/sZCPHTKX51Wk
Bn6IfRNhbwuyPC128mv2FRyCm5RI+nXxB7MtC4WMxFosOcI8pjK4nsr1mAtSjMyg
mS66DYzhj11Pw89p5V9jI7mbIexpWq3Y5harBEBjmNjW4HSwLo8kpJH7dAWXpPWZ
YRCEbdhBsMYiUyWq6QVXa1p7lNcNGsJDIgovk2WKc9mwIfSbcwvZ8s/nrYt8LJXd
AjQMwHV2Zu5k26ozi6E0+6PBYkuMIbwd61hzJvsraPeV7QWi3mKyQxUAZg0cZQ58
/w0DCr+eb3PlcC5ynMaM/FIW323SvPEhNr1H1EtpmJIUrhP//oBRwGPMiyj6nmNO
YqjiZekfCsIt3G60+/RKCD2QVYnBA1YPmmOPysJfIzKriQDy/1BMyOLJvIsfaFL/
QRstYi37IaHYWBKI+ME62XAfCtp9+lURyMZzAuK/XhmnASURgy1/eZ5mpGucfLpq
ZPg3AVDEtoZ93aVjyViMUI+AWtYGTZKSEsHGn2t5g49E5WBz4nFXhpfWjSNjTm+Y
9iELxyrTyb3IVNrcKPEfY/TzJqYUZEFkKWU9w1fd6/BSaDRzv0TcMkQLAHFT1QJ/
yyi0x/N7dGpJ3xtmqHnLGpQ0l8+dj3x45AvmDUs+6N0/l/3lryVIRJaOmyTpz4kB
6rE3/WAU2uuTa6WrbuPzh2FkNz4A58MRwHyGyMQkbwfeSp5BauFvZK8TAPipUcev
m1CeybFawsJ8tzxCe33KP7shgeS5OFgdUIsoPzCLJXx+w5AamSSveGL1Z3F+ww3Y
zYQnwyE+Aht3u4gTki1bSHtDq+mbXO3acqTmcJROVtU0SN/mQkw0pZe7X6e8GVeN
eG+68tqSZsOtJ0Kcl0G0ME0iL+8Pu8sQzoY43KoRsgNFUVYnGDmgC8Zyxkwk68gV
iDupJYwuNFP/+soCiwNEBLssrbphomyxwISwrdDHCcUFQIa7aB8xxWMxcVRSLiLt
EF1kD5AdxESl7V2OB+f+r0Ebejr86Rgsu5PFrrSdQIDbbg7VwBhT8tRQum/W+akJ
UMHx+emBT0UDCjlweCFSGaUmcOZIVQvQYIkz7uhUg0m0WN0AOJ7REyWiuJx8owb7
p5YoAwQF2YBF7Vn+/EiVlV+92VTadKck5Rdvq0BCsK56yueG3aYrFXWB4TdfRTPx
aQA+XZko488wahATBufK2XJHlO9dOKLr63Cqwt3SFcCwXt0ZbhLKVMYIkcY/vvI1
0xJp3Xbrd2Adh6hQotVtjnOyLSpcJPPL/GihAmypHMFJGG0aMA5l6VhGMO/bQU7+
AUeEF3xG5bllYfEPA610o9j7OMnCE1o8IwWZTsEiI43a4Ydz505fH0KbBrnhdA1G
WpUQu4FFHnfCPha12A/8qTLRVTlWpJjCOS5WCI7Q215aiO3W+XHWct+XApKOEIsR
fioyLHWRwonWZXZPRDQ3hUcYnkCuTyH+2bOCwRUadqdLWauxI0ywa+jinsxZokDw
lpFfd4J2Z38nvKZJ5caIgfZKQVmniIjTRvXS7kaGE7MymBLzvy0NMYaC6xRskGiO
N2ebiQJNCXNCLoHAD6IYOtVWjWEnUd2pgLRK/pfCpGIIj4NoUvrAxncj6ZDqQttD
PjeSoEkfvzJ2j8FtF8r9WBpALOyGnaaoe9X7xvYaybgu5Zh7wstjhfZW5VK/WIx7
I0k2ZVbH1r0ahRQDaDEp1AVm6WjF1xMsYa7WrsBMv2Ym6f7rCtVwD1898mBx9SMV
idfWAdUSpj/4qI29F/ZltWcdBjEPYEt40/ayejUB4l/kdn45R4DyL/NdE7VUwCn1
vSwLDMnvNnnyq5F31Ri9xFrnRRW8dWKM5gsWFb0quIWA23YaRVFuTUGurz1YZBok
AdSvzv1hXpj0ObqP4+OtsbzeHqhUaBEhE6IX26P3vZyOiD+GiiquvireHwFAhG1m
lSwnQ/MYA4cYZdrJ2gPjHg2oAfK1wBlUlHcjgAoGe7nhudtWlzWy1FCYLMWOuGgh
Pg2wvYAZB7XFplg2sNzNGf6hlHqxC5ngeg24qTBXqQ1dBtYDVnKVZAboKPJQiDak
vrcLTipBNVs3ybHD9HSE633YwbFT5QBd0vYPtT88S7RJ5Q++bcSjP0308KAkFGEL
vTpGOAXieUmHNwqmLMhg5jaisyIoXPPyQf5lSUofkerEO5FLu/qiokyykDCKSn+r
SoVkLTAXNEtYkXGa+sZLplWTOAq28FATfJuRulZXk29zzMmGrfvLyzZaT6hB6zv5
4AQGvfvF7Bb36mhQoYYovkJGFzl75wfTh0sKDMd9erzRw8D77RVdxTP5arwvj2Kj
y0w38E0aePjlospn9Z1pwoqhnLaXQ2cYhzMgSoMFTY2IsKKYUqCMXLkDb6UF3Nxl
s9AJBfm2NxALzSlIWdYZoRDBgjz7hB3pqCFdn20Ipbd2O6rUMj3zBlJWVz2Wl58V
Gb0NZ35kCW2Xj+ZFLHt6CObrGiRK2vjKctegP7E4c3A2c+KDs6vMFJXXYRS3dJk4
c3y9ADJa/V91pJH1EtQveURYOUTZSfaFL8dc0d3Y3DTZdPsus8/E9xhgAlpTdUT8
hoCxBYlmUpF+Uoh/HkXSrOdMEM2XQefFOTyl7TUT4JnuUOJkWXnuWTyRcM+Ed75A
Name7DC32FMr4UrDJrbFmdold+rpEBNPWMssf+VN7i++8TwdKwRRv52AMm8OCBxe
MCxDvxt3m76QJiQPB75UMBzTMsDhhC3fo2PseK3fBTtsxW+Ldpa5DJw+I+kQt8/Y
3B//6fJXsReMZY8vKMGGK8Ixjwtku7mmVuTtNDsXz9X7jLSDEfdLp7/XMqji9HWe
Z3GShVLM9Nz0vuBzu+WtQb72NlU5JFmy0oBbkO4cwF1yI4HFhcFMU6ENgWuyt86z
NYqpQ/m2LL5rPpCgliIda6lu7gxTOYCBkgN+pn1WAFHJuWFuDhui5kTUIOYslLdf
SZ/rC7OF2FOYrpHc53kmM1p/OapKcaMrAzhmYWvIK9fnkMA2m8UaerLVzV49fWeA
5ycBhNRzwmsETBiqtXX3dut12zrAbWwe89GSx3XP+Jcfn2jLVu0Nes/rqjcr3ZNN
5KEaWvmm7cNQQ5XZqiM98mMcfqooX6hrIjoDNY1WteRO68gLtggF61nP4zxFWD0Z
FdnI71L3YWsdCEaBVt1lUQBm5X3ouuyRPbpcHFq1XCiiJYnpR7RxiaCvrTAD8n01
oYncOT6fsNUIMpYqNVEaeHdaYgBUOCa/fkc4tc1vgpgXyLe2GQuO2J8nciHmurFF
0FKe2hsPLwQzZAeRwlZ14SgBQdXBqYL248VW75XZ+06HW6S0mbqKF5D1/2ViPY9p
nggzj7kgcdmgw4LViqyNV9+7EvP8QCeb+VLEmBRrgn4feIQtzGQcu2WiytTFVRlM
a21Jws+xORBqsZYUQS3h6uSAoJ1cfCzPHGI/8f3fxUlJCyKfqCelz7eRTHZWElav
q7NG3HcuTI48rSNkGI3eEcgIT4NV3lgnETYXP85fEPyPrU2I8bZ9VITY3Mo7TXpM
hYnam3MZ/hqSnln8vou6iGxhmKi+y5RA8jb/WsInDmIphbm4OqmTI/vGIfXn8imi
yBpZ4I/L26bfMH6Gr60d1nsh7i8a5J4vAN45NPm718mlfFATaUXBfnC0fkGE35V4
Pel3aFCoUQMuBKmniSrSrSnAyYqdkU016abdj6L0s/aMqR8V814kJN38ycy/MzFR
TcPAF3d3/w3SjcUulFGwlcnZldi8/nEajhrHMsKnRcTyIt3Qiaobu3u1j8Au7WUk
vrLkNy7luJqz4HbJMQdLZE+uzZoeuWbAqPrR7YEY01qmJJKRh2ctK3SBWQkIUTuD
/JXgBM2px++ZMzuaeM5br0dUtNos/MfwXvbaI0vwDFsLwJ8KKJyl3qJjMMO4Q1yt
zNZ3U0dYUto6M0urpnAcP3igzD2c4V0PGs87urYSlMfqpQs/kBUdnh0Zc0ZJXAmu
fFVSERkqixCIvkTr5pz0RtPgKp6Tu84OGXqzqbdW6LSJMkdF+CJYBmWS50XXQq0M
CWAvC7HZIICA7fCFR8YLg7cM8f29S8zM610F/tGW/Ibwex3Q5o1sTRf3AEjXsbPw
+iVHSICX+dOTBvaH7qrNH2No+v8AMwmuflpCQ5HKVl/XiCeJz0m7zhRhuLmXmw4f
ubRq0H3JuGTILAzcMQAbvQ7e7HbWYYKbr08rEs3FJHstGMIrc1vGzbzlee9/cgod
blmITeF6wnnxyAy3bR1817zdDyWmJ54+jx6CMEsk3sbzaBgfKs9UQ8dkNsCSVkTH
TvOsWHW7VRqloB8ptf+oZ837F5VPuPVtBeN4u7/k+O/yO2Va5XzlJE7tI8Wgo1cM
G2Bg0rcdX8PtocjfihtuK/9KxkCNNpa26qXlJJN9cT7bV4N3ffQuYUatpjI/FFXx
C7ycV+PCAOv9T7IVtMRX7p6SIdFiDGQqecIR6G9Xl4mmAlUATcYhTX5NcwRSnCLj
X7msqXYXKcjlT3g6OvNZTroy2TANI+F0/KQdILwgkGO7TGdM+UZtoihu+99hjR4X
kZMMBFdOcrbAqHu2qX91z+3tQPqzD/QHioDF9KOvvAnehcEx3o+QVtfON1gAbHPb
axy5cs22C540eRU+vO78QEGsnDYfZvmj6GfZyYJX6w6ADvN2cKfMUy+mMNzv6LRv
IWUUUbW4KPGT7qCWPfqK9q1NLNRElMnPh5W++1aJsdjVRZFQpvSSc35TCBPeEUf7
buYJAohGrVl0Svi8KJr2aVlaJXU2NcIH99WqLrBTao48WPlXxS6JOlwO3S/xunEp
9IdzVZmxZR61pAJNDWFzm2BQB9ggxog/S4DFPiaobhysaEmOl5ALpSMtpL3GnPsL
ZrF8MB4CDvBcHsPi7UzA3w5YDyApvV2rmj9P+EOPX3Zl/N7qYeUltx3e8jBeQKI7
6TW3RAjDMlYGEuXLpM1sv8Nyfywmc+M6+x9/MNUENvtUVm6VePlKl4U15iDDgnr2
7+KkvEldhC0W45WWGLuAFvWl+8E+sppNAlerNJEZcvRwnXy03fuQAoEZTLQRSy82
gjgIX2jVPSgKIsfKwBx7DMgpiM0dLvdcsIrdy6WxRc89zw3kfqoQtE0BDUEberJF
JdJmOvDCmgAkj3NXAHWe6iLfpHB+SlyB5RcMmz7h18AN8JnFlhsOYZlr5gHhF9r5
ryDLK824S8cljfglDyuIsg9QqCFJcM+iuhBOgwXujlxZoV6JywICMYISmampW2yZ
EVYYCCNmuRXmT+7QtDLqhKOdw7fa0W4R225jdw67WWtyJn1IMPqqXkSW3ba7bsmH
dIyQoXcEaP8uDJE4qre++jBlET7wQ2FJfU2G10rbgpNT2J5eu9yTTdyZeny7MRHh
xBz3SGq/xaBCbF0yPG8VNF9pujCkLLtE8c7H3yZvmCX8isV19fIkQAcGkiZXOLac
D6ijeTOOva9m+bBEUYu7uaNSg7sOBYIVoMn7vL/3HqQYyLZjdz5XlfYneOovU9YM
77Kz+j+cWjpRTWKiz1HyQG8W2hWiJdTgMsZrDEDUhDFdQtJvLD0oSEPkzsXLyQqK
Qznnlz/e4BPBIBl0UjozTiOzlLWVSg6qr7FODe+HuCvSYLL8Z7Jtvx/4L2pC4Nvu
kz5xZMrWSFAjiiksF1GQMhdCMwIVkTPAts439t58zk2ukiMK0qeK0Jy0/ZU1pP7o
GBZCsocMSWYExw5wDlknIIB6WWQvXb0DoFWu3pCq1BarsZjIHh2d6j9vzriG9GUO
WzbNjhch7nKt4eGx8T4G6DhkZg43vUd5WQL8KIZNs1xAtBkriitycS+2Le9kOZTN
CFwnzkKed8tGSONhmRc/jxFeX2Ebg08yRkKF04M91AZ+83ehmLFyo/Lwhx8rwLWH
+3juq1LhI+HlDvIJR17P2xaEVNOBMA5SRkUMUOT0XLD8wY/CQBdn8XnjtWaxCieX
0lRmhNkwDuqQkK122lvP02WZbVvgXHW0HLpMaevfRFusb5QPZKGqn9+BPEXnBuF1
tfKDxxQRXl8EG+EL7rtCwKIx+ASqbBIwC7fj9r4cwbvI+7j32k7KPukPBVOmV53m
WPj3qLZxS/g4QBP6ijVV9D3PMBso/Vfgo1Gz6Ytu8d+bDGjtmzGouBOensJ+PEw5
UG7Mls6OniF0/Z/C4otP0Sjfu+m1O5jbV6aS0HchaaO1CKMgbujjvXr8Wk5xXxNO
Te1UGbAgLAhNh6YISaksRelkb6F0Jr0blir6Cr8abnYm+8oZ+vNtvT1PTY6wJTZG
XlJwyrPGV/nNwkW4LPu93Aot5xVodQTkXIKcCdwdMZIsRfvR7H6dAECS++KC67FO
oxqXV/IQ9tiFHAoqHAhYiH/3yu6iuBneY6l1Y3saJg3Q4wgIzUbCr1FNGn3+jMGe
L6Y3okK/bnJYU/ZluwANbhvbPfzpWQar4vZagGR+2xrZjIpamJFHepP2jYGcdQ12
IYTIGYczkRw5zPeZCLUaPdgcZSFCfcoHhwB3W5DsXnfoAeWMJBxKujZn+KqGPIZF
S24V0qKWTulhx5Ad1kNlTTzveqctOK/yQHyqlfy7TgK0mCW2RzG4nK0vc8YXtQkH
6y0WGuNSoI3SGul9maZJ7dld2rsSW912422h7plupges3ig2UfqoWPXxNjTWk8wG
+lDXSLjEdcyzhFsJYUVxDFOvC+Yz/DZ38FuLzmGJureRV05noI9aQr2YjnbluPg5
N2HlNG71i3p3k2axxUMXsdgXyZk3jrmEU1N6g+8m5sg5j6/rrMONzBL7jEss59Hw
VASamU3vOm5U6ilW0Uddhk+EvVhWA/rYJjasqohoryvh9A5mDOFHlagL8i6oczd8
TBsvWslMP7eWqf+/P15YB9uqXiu0zAyirKg2x9KbDpTGOZmDeB7r7t3Ff9swJr1K
t1Iq9nBqc1GsrIQfXxVqdpVKBpP4maFOROHc7WEkmtsw/mJyMvsjI+b1j15JfItk
kC6clxGo3NRxjsbdiBYRpY7/P2IE1G9bK+7PQIrXNsZf59rvhvtN8UiT/r2KSy7P
cRZNUmR6LumGw6mKKU6CnhpXXvEgdfTsAKrg9GR1xWR8ZnMMZEscF41yHIeuiTkh
nk4+A+bpTZ/FNJu7cJDgofnZ4qsINYmekXNarJojB+YGNI9lspBcHNzdFiXldGAo
Ma8zNCAUpY7eUL0o90gAxopz1maIiwq5nX/eKH5qzZllmjEJEAeWUodAYAmsdV0a
AFlsIYvI8m5iODAnXhGEpzC60PpOWfCrWQpkvsjalgNtt+6viOs6dXB/RdwFPPH+
lyEWqpAHQSoMQnqIH5DwqbU0+asqw+ltl3z4vP1ziLH0tyZyDJ0ezVMYEKyCVSck
MU+VBznHViUlKx/3Qh/RwkbknA7UYOwJnmC+AJPxEBdsDsD1rER+wR8sOm++czk7
W7b0FrJ3crGqW4FHjtnUmvyKh8VWAjL1HZb3w6aRNCZh3PVHlBP4dS3w+mmSrCuo
ADqrrv8GGt9BgS0URe8Adw0pDCY9ZITDLEiSt6/QM3RfhFLN/Nu/5U0gFp6lgNZ3
eJrMff48p3TJMzRHIGNr1Ghbo0M2dZ9RAzvHAjpDSJY5B2itqFaNUynY+SXRdal4
nsDR4wE8oHXcsruIjlsugg+vyFWxY3MXQ/7xTxXY6Tiw97U8UCAOrnv1V85JGgpB
JT7MWZjYho/UAxRUlZNnhpMW+e46rU0E1sy8Khhp3KU/s4Y0xB9ffOi1NYqA6le0
B9XDmq2vrPceoejS9WRexW6aEtMLFXlxBBQb4AmXGuTJjOVQWGy6nvr2GETlPXnN
BLs9V90BTsZlWgsnl+HFP86didd4Aqp1jj7eCMQ6Ms/Kg4YW9MQAPd4qBA1weOGG
dv4fIawctdC0eZMENdhfa4oyCGvc3KmPZzl/8dNzM0VqyKboZPCVldJnjF2iHGlZ
2RBTSFqLMUqw7DzvmWWSr2OdIIBULyhbFieoF8XPfFZ6S5bAGpWRkK0MijveKTAx
To7Wt0SA1As3rEU8qUMfMUwTNX2Sti1KXPiX+CeyU4hKOVF1IAgbjoqnzUXe19Q9
am7ymWCBf4ye6v93S/xSEduOssnhURaHLDKYW1WcP4LPE4h11kaE4GwIYu3a9g+p
YPgD9Jh82V36gEj8tnNUYfBkec2CsOTzhnZARMKRwM50mc5yfhmbIHg6gwOrrqpD
QcCrV28Yao2syeY8Q/ODB5fE7XfUTzRUqXGeiK+KSGo5MJoRupuiF7u3908eH0Wz
jGKgjCDmb08Na+yj4YFg4XnSqnOBOoryUmYoNfDL7OuZCnsXBl/KZUR6bqBzsnCJ
/xJ+iVg/igr9V7k1rxD6wm/f6djN0jJ2qeyiuZWh9CbD0LFpivVoMm/1yBQTAI93
J5YwEPtB2+3PloL/jrhqHhJ9V4KTl+fj+oVgBr7LqZeDAcxyh/NPHmB6GQ4aojXC
duqv2aA1LLX+REMJFlH1wsd49m6YnGPs49d9311jSzUlZS9dwguYj7d5DA3ABW3B
dulKg3mcaaH99aiQcvrFIUebi98uEZ1b4HVfSga/0mEzl8soVkIdxj8ClUzQTf0h
Q180NokuuABryTxwPJBCs2dwRQ7kDYe8faBo5CXUPvDaPMyexRdmqeNjQxXaCGu9
lfzYNyfIkhbvN2xliRaiJv2EmrXnwogBwR/lnCZmLS1os4HPPShY4qWQLLRf33mR
yLSlZVJLM701lZlPkQDmJ4A2i+WLYf8aW4iXG6HQO2imJkbfzlx11PNqxwU+fuaa
9Jyli0lan+sRey1UouIfHJzq2DLPYysEfYX7EKN92wQOvCPeX68pramTSpYOLnCA
Jm4xDMSPlJV1hdPLtlBn5s/cZbr3UJ0exPYJaN26Y7kj7yB4/zYn6MkwuP9BimiG
eWC2v/K3Vjwzv3UcREnuejIKbRQICM78JtXCEZ9VsOKikjJicFn0voRJfGalxjya
H8Qlhzn7p4CWkAS8UomdnzOtA+Q/dtmQSP08Ad8OlZQrn7I87yyIEMQXuq6374wg
Q///3J4OtW97/sTJhUpErqHGZoS1hkO0RK/9WKNbiYGH27aG7Q0vCoTIVPRSXUGU
Yy7uoETIfnl2l62zCjRLiHZpXoVCVncPWTnKrP+rpJSYci96Pt8eTQv8vPccb/9o
ZtaMBDPgt12wMnuI7sl+hxbvb4979EVKFYgeBvENtuC4iSxMP/DqFouvei3jVIbm
WxK1v4amRZmHlqRhJyIEu7JKD7CtKtpfmSE2cE6daGhYarKD9X5krUeGoYHrS5ZA
hGfN0qR6JLeGqvrbmjjo0xSy5Ydb1P4ICIsdaufV0zLqEo69kZUObuU1YgOurHg6
Ps2GkjNiGDCnrxA4LbQMEpvAQlAaLo7ZPNvbCRFbLE+eu6274FEg0VJ+WcExT1Vr
fN9/FE+6BCsxrnuJub1K+a3PIAJ6v1GlbG60dmDLxbhNC7y5asHpr2TXCUX4CVMi
XdAGUqk/X4O62ZGzLuzUfndNeMS4ULd1IBbJmd7BgEfL1I78Cn/GDsSo/1nQUO+R
StA2+mRS96ugBbmEg6G7LkIqym1XMnDJrtqOEm4+Zg9/05cSmVjyftGvXY9rMyio
LrJAFtlvGn4ekLSF+cr+KUDNTgMdBQJdYi/jqEtNbDsEUBrI+CPQgtcNumicfaCK
mY8DJkdIAzonwmLU52+CKFHTPu23J8MJ0f31xADl0kGW7iRg/6pZUj728/nkvpXj
8gZb+WrHcvABmNg3csXUv1fma7vJlqk8Esujsa0UvIeknvWcJXh/8+FtsUNs4+Xi
xSk0r446+jy6K358+kGzKK9EByAc/U3teZpW4MsW4AGRbWRhNubiX448UW3yckS0
tSAjhTNsO7hiEmtmXvL3PsGRJuXVtJWy0Iw9Ws00OlT4kPTMxXBWYnIqIbGdh5E2
lJ15Fq3sKPSvnj5LZIxdVJkoZ9YedNid/kUQ3S+3Jc7saQDSd2KYgMS4JjQ1YRhq
gQ7P4v3LeQcua5PY4/opdQYV6LlHOYp6kSnK4TmDDwEm6nSgy2mza9K+F/3NuqiI
fIrs0tzX9dRPZom7eT0gRajXpwUZ3fNzg7IXir3AeR3CMsiWeKTToiIVJjbS8VM1
IhB2Fl/jPKljnGzMB48CP8JqxXxDkOxGNjmnYNSqZnaaj6OOD2kNNI0Ls1BK3jBE
/GkHPhpSORcR3fU5WYqMI37Y3a4MC5Da+fAsg8f83vbgOqvej/EyIoglOyXIa3tY
eLngUCwKr5RKltI7UB4DcKZ4GPXbq2i9dGZS1xOMPwp6CTge02PwmLDxIioPICBH
L3H+kMm7jW72leKvcxW8LCe0z1fsHU3RRAuCMN1m82Cbf6wT3T0VBRJ+2jiBecNh
vY0X9YVO+55wL77ssi5C9VaBeuEDhx5DenDUt+5vG/bC0ZIik5Hxib9XhL3EsReC
NZnHoi/XbtLFpksFJqhTqqk+U9lx5sE7PbwkHeXbkaW4k+2THGRSaW91X9khMpC1
rbS823/6XZXwHv82h5llhT8BOfC22oMORokM7xK4XWVdu71B/ssY6b4oUqM6q7el
84Uc+t8jQHJ67CFFcfVgNDd9mJPuZ7jStLME6x+4gT7aoFRyO7iy/lsy9FbEjLZ0
X1YckZiErF10Oz8hNocEALI4jnOO4c/1NJauFBnWDzP0WTzYSl5zfzfjzgamBTBC
rhbNfcpTu7mciJQjimw5j+65Urq4eo7184052KQ1XNXzQ9coaoqa3ywmmISZFnk/
BODh23ogwTWAAMDHwopQA09pAZAAOrZCAjxlVyB0tolF3zeXTD64uzLM4PeBeXlz
Vl/tUP43ln2vAx/Jo+wRSxUGLPvKPlT3F0g8WdNL7LGG7PnLQgpPssiqPy6FO1xZ
CRWKqPHqbuJfr8UTO+0+xidKQrKl6Zg0zX38LzXIALl0EBz8v8kgQc0x5jkLL0Fz
w08/hBKGCrTmPf59TWaqs2nr/B7plMNZ0PMTdJZQ5+TM3jmhwgBjc3ee970qInUD
yriVy85Xg5sYJIUQ/Opr3BqxKDH2cqX6Am6MR+J3bMRlKvIas2/XRh2eQJqlZeDq
GuNMYcaVFLoVNnncOuUwTPyKIlgtA2cH9NVc17GGVN9akao9IB6aKG//AxxmEKss
G+Xjg+6knAZKoeHlExCXjBkWYXKyTSJNT5uDSHC5UhJ4Al1NUOPOQ2WZOSJfFzoq
2XZSrnpOdqJbCK+m06cfhR/QiqJ/sG9V4WXqIpZ7sU8CAfJXhb5H98GwRsl8gzQR
7rO7MXDOJzqm/8Kd5V4RgYhLEy0k51lB/pmT7uPL6/4dMx91EPBI+CN7ZV6cJ/xW
vWR3SbmklvbrngfXh6E35qm+Zz4+EKlMeU0gy0ZsybSKzf/bGzQqHEVf51HJnWie
12Pv3PHZGbz7i7dbP4t4+Y7AtZtADqI1vVWG0wLdsBFwK4ihsiyRouHpjqVUNvZZ
uL8qTNJoyB9GcTZ6ThK4lFTMvj6+H/oFeAdWPzmGl5P99saBoHyDQOmwjq1l9XU4
8dYauab1Y7ju40Wyl6kcqiDVY1ILC7CIyFdOezW9T0JSClu0loO/uE+n3mza3GTN
TbdgNpY5R5e36wnj+cvPZTN0ZEf//DH2USGxiw6P0P8ZGTjUO7GI095qDBf4QUPH
3xejkGnLYsuTdYdMBgAui1pywcXOjfD1EhLe5OsIhi3PTkgfMO2OuODl6y8IrGlk
/6qWLHJkV2qyIG0QWAErmlRfEPrMUtqaS3A0SExaSQeZTzIqDRfW/h5pV6+HZoS2
SzVIg9Ew/pH/SWvacvTW19UK3Jx4TOASP7Qumap9E8RC3XryLsJwKaqYTgpBygGA
LUIyCntYeyLxyS7QXbMArhliSu9Q7IHQhXOobp4FkyUZgFXXnQo3SsRHv5JXlPar
h34e6jSMepT8TFZwwvm54j9Fu6wiwQPBv05NAJhI65NvwSddKDYmEqE+gYNQco/E
YgvjyXd4eaWWpScmqBIEDUn1r1eBFmxQawsIBMKhWl3ntrCKs4DFto8rrN1rXnJa
S/ORKpA0g2hd5Y4ZkUxVqrq4hPRpQVVM+0sVJsC7V3gQrSjta6ut7uIOKiHqztCZ
g/B6ULGpzU7YK+/cXZAF5RfCwIXO7lpN33a55aqKJ/OBNp8sJFLh2bEyCsMy8BcC
sdTokpfPn9pefiqmGoTrmKuOGQlj7mKLziiY6JC8Mlia747diJNfk1npfPioTcTV
QFHWK0gL7PDYsMkCJboAe+aS+DJroWkarEUbVtdmeq1OfTuOGQuP9+vZ1wZ14c1m
ANrTYUeXsy0KD+hsGLE6YN4sNpsn300yoWmR+Aa1lwLZtZlVEflsm0pKViSpEx5G
G6JtkrZJ17dMk8E8qI9j8wq2vCssLiIZoy0OZ8pVAmvac/DCTp8dX+tZ2tutECD/
IPoqLvwDdHrdPBL3Yb2XosAFIyx57qpO06smmMtSSghnqRGpGMC0J0xcc6g+TTFk
FwhZpU/st1NoSiueYbbcGQksM2Mfpw2oJ70hzV3sWViEQORRniOyxdqggnqSgjUj
YcRznfZbrZF68tpnFP0Nog9NIpRJ8KQltyjXm9NU0kUKQN21rL27n2QprBMr3AV9
NR0nQqKdx9OGzVTKnYOKVvtVYixsup4hdQIWy5VX/s8qMhS0N/SO6VKiC93dmohS
iYPk8lMlv0PbF/BYSUJrKykIAFGGX2Sfg1zxuNCSJ3MuP/yW5N2Hufb18UFsG0Oi
RFHeC8VTaPdF6504TLFRFIOBWm+5pY1HuIQKxu4JdDXVusSY1EPdcNeJyhVgseZS
nMYsqba2JQMyx67Kl2ZNlSPXuy9ctR5BuYCa2gjDvjSy5JthQkz+20FQzqaELiwd
2ywS7EQRQkvMii/l9mW06s17w120Y+dUr2rh7uRc0xtoid76YT4Pm16J8EJo6C2R
8iH2danW+rjRLjiOfFVVnDv1vF4HhIGd8iuexeTyxkphK3baIT7yNVzPiEu+WB5j
F9OEAj7rfhFzcbfaJ2loRmUay3pjNDV7lMr9cwK3Ui5XaxWpygMvgqxRfJLiHnDX
sXfU39c7b6BlNiR7Lqa6GQE6u3N4Pa8DMFlOxsbcyoPwepsEt3TLXYj0s902+t4w
qeD9Lg4J/aGq4HN/inQg583hRZra2YqIT0B26nVL6OKVFrDeLHcuWKwfJseW+zNt
9CEOe7nhIV++on2PFT2woSj+0n0tFG0vuOjZ2IO1dK9q8uOo4w/VgzOpJFH8AQMM
8Gphs/TLpSUaLJOU0jSKqLJjJdbOVdRpeZxKJpaVgq75k7PPjbbrQ8oLt67QpBXk
0fhrvRHuh8by7L2ahMLA5OtMdGeIwqUc0KIzmDG6YKgapxm+Nbk6aplHWVef7SkS
j8Cee4S7qssv1cmD9aBAzEhZ8oedfdfub8atY+gBOQT9mzdvMuEXbU27gh760+EY
uXdNPSSdyMKiNyX8lgs75Jgh5KwOjjWkXNzHnUGshy9PVLPAjSWr2I3KoWkdmPP6
Jz2stVlAWRH9O+NNLJ0MiRn4z9y6heZqOSjFcxIeyZe5ADL7BhGkBJzfv9h4IOTf
X+nIugPI5MUIOmATq6hgONCIvj7+XOU1rq4IOoInWHLQBl+6hv/GJwWWLTg2p0HV
r3wTOQ8XmKEhKbLiwfq4DHrHGiHbcyRJGoltDA/r20k1YFKXsdTCoVZamFBsbFAv
jjGE9XQlDa41Lqb9z/JJxeB0DDkzQl84IFxA+fC9m1l7N83YHodhaSOKxJkyFRtB
uhM9fMzmSETxsEqj5W0DN49TTPBzPfgesH9DI0OnUeU+/knWl4eazTw3koio+Xsk
TU/IRgAmUdv4BVbIIqmHMOXeTMeC8NTaHift2U50ZUJnHrI1sLT+GCDuYRhww9HD
LQyDIxGdIS1AEHPH9KNx1luPTB6JSylx3A7QiQaGBcNXE9IAMAhCT/3SJAiImWUV
B5iiZA+DKQzBaEE1mzXYTiFWviMq55iNM9TZPP4P6889DK92PFY4LmdHH6nLeNBx
j2K7eADqXK63s63E3muQD/0v4DrcoGFgUNPwR7+rgGTUxV5EGssoVHCBJi5v1zIQ
5VJz2VucDCcBSqZVsn9g0ng8GP7F2jqUnGxtTfS7StDJgFAzebKQBQlHkEQIUYSs
b1oXGTBgQwRU0dFWLeP8tXpCvd22QkFXmHtv/jbpcJB2Ckj+SsTwF13HfKrixGqH
uQbWav5MICDPd+BluhiRseC2dq90Ds20DQaQ75BnPeywPpM2G5GZErmR1rxG41R3
rjo5ZzVL3V1lvbblUrV66+jFqmSKhKGi/1dUxQ3BMSgBYsZa5kniByA2gLrbVqgy
abyAEN4Dhoxijh+xhNG/Ylm/fdwtHJUi41neO/MwskllhAjImxAZuxePMkqozO3S
5jJ9EcGHt6ClI1oubqLeSI5RtZLWaUGgHsWyvNuWHpTha4oMkSbk8xySMI1Ii+As
IJeVEfde6kQQZ3XXi2To2ScWG45lSlaMxd2UA7sn5B8yJsyWhnPxTyXQONk5yCpp
wq28qulAN1BLcUCU0XGPM/yfcOi9+WFrhLWW0YCFHgrsiXXlE8V5iex4+zBK357y
qfrFPtkntB2ADuL8uXevcQtCY2eKQCaMb08p1nSPBll+4a3Le/7nY5SOSsKYxe3s
E5hxYgV197XhAEFXc65XX5WOYlopQWCg/UIJwZPWLNsOAyaIA4dMqukOW5lpLH0z
3HjLt0eMRuKCf9fO3mRj7Em+G7tQl1IGUviE9wStq0zvoL7Gy+9VkWG0mShxAZ5P
EVb1Q0jaEUnKpNRduW5qGo6wtzCrE/8ZTDN3hKPKyHM6lGWp8Kg9zdpxVLyM/SVb
J8uHZtJYisFYmb8j6KdbO35LQakvtm7RpDT1y6HEE3d0fSPRcJoBuTXNFl0QXWiE
H532+j2OFfvq/v5Mc//kVRIXMMC6PI0kV6AxgidsdsnfPsV9ZQrVlqx3zyg48VsT
Y9mdOzoARm40Go1dvRQ+kPswZjgOtvGKnyP+WjgAxmdaz4BsaMz8MGJG7XfcJv9z
Kliqb2NOcH0ZJJcxl5hTkIReh1y5oxyZRfONdpb5Sai4dmtfUffTRGor2OrMZrpo
EmbZyyBgrJqJ7Xa76mzXrusB6Du56B5gCqfwhKtYNoHrtUkOYp+jjarg8Wsl4dXv
P3bGcEd3RoEjpiG2DRsTp+QWEDdqh66+YKX1U1SdFAMlCPlOokgIbjZDUBgxph8R
9TK47yEZQQG7aY55r0WR6g7/8U0wSpMjuJWPhiuV+EsbrpbIdvpkMjdIBBr5IoyS
E3UkfLL8bleH8jWoIY3wNMhdZ+0CLPjEaTlFTH9fJ/IAebdkjTp++b+pMjvewDFV
zNb3xiZoWywvnwZQdVDprpmGLqojdappmQdQ4+vIqH2RFhe62NOihp+9kYTNxq7Z
Bpp5DpDkvDYSZvlPcOWRj4YBsxUNzoRUyfwuq9Yhw5UnUqRlNOWX4BUmGVVr4ydk
5DvIFb9GyziIUZfDBDuIuMn3zSX+GGL5CeVP5R4GFTRg/WzfMrZ2AbNw0a3dnEcy
JrDfDE4FV+5M8o668/iHmtMsGIiG3RhR+kkakplFTu5vv4zkIVVsRc88V7fUr21+
e3T4ukwIQhI0kev6+lpMjHwOJhFkzxKVZN8H58QoUbPuz6mKpitsfKj2c6+uoUCI
sxpLyC16PIGeok4yivnfjOKOMJwvY90ztIg1RVTLHEItBf9AxNrqxULkDeD47aOq
mBLWYKlwbzKk6yyYifuIaBrqotXf35g2MEiFJEsRp22j+4mSPHN6LlPgSggnTOx9
TLNoc7AtzVDAW4jnRbYDz6ldgnDKgCr6Zc/oRB/oKfPFuAuGirQYQO9lu6RpgxIJ
Z2LgvzUq5qdqGUwymEcSJGVqEWbf3ThdHVLOM/CG2AQZripjljKvS/eifAdsHwgY
x2lCvvT/CFPaReRXb6pYxCDW1IBRcXK9+H1uvUfB3S5eY55ir0VghSn5LC01Qnvt
+9gXReHcVXpQrHL3B0uuzYRSh54kfr0EyA2iq+Ph+sC4gWo07YBPMM4A8ukSk/Yx
og9vP3dBYzGEKwzrzNgQFtYBuEE2T/WHev0kuGsZWCqR9ws/D+uqsp6j2jAP6faQ
CL1zQMIFRM8OE5mqp4Kw/vTK0k688380h0fMu8qJ1ZxxLil7mhubhrLQ7B0be000
rM4HH9aHYQIJn3u23if+WtP1FJ7GA8RVmXVtFK1gGNCJ+A822dr4oTgfHbbPdC/U
PurXKa7pZ9bw/FKhpjBj1WB+GY24S6d/vGkONntwheWZYIToQ69o2ynGeDXAx3I3
v0FPj9QB5NZm34DxYjBIo1amUNbsrBUm1cAf3k6QLSaF11W8LvkQR9jl4PjKXrBh
3UEdXDPVDkpJYctyuJC6DO1lvNZrr57GQSNb/TOTKDd43f46wkIFI+OBqRKPpi7S
bn1umE3l5RXXBTiVrDcV23ookrWkfB4kbsv5PXGd1VMKTrS+juEmiX07/NMjndhF
uXMyEMEad9y0u+xnDwnlbUdPQ7tWkdoC9DyS0KWHG2mEl0WUujV3mht01zQMHPpm
NGmXC53DFl2Z9yQZhOXZ/RqltJtdWzFsIIwzMTCg0eVI9CMU5RWbexBM8WRKAoiI
soJ6O7QCcW/lJqB5eQqbcC3xGuW7zdUYtiho/ciQTIwYcAp/96cGUWfRhmo0ePq8
zuJyb3+48Sp7wC5FgbuzVW1AJOI2DvpZrisacLcxrVD/oSloPD768AhEs5o9QnhL
uPsVoOW/SCtZe45NOY+VZ0EsxOq3WJB/tVwHAUhPC9TXJ23bCpb0Pm9Tcq4UI8V1
hsqKn/I1ethNiuBr+43MgZEOfwP2OCR7lKRzEYDyHrh6itVlf4zTbzfb5ZH20/a6
D947C0ZKUiz86RJjroznMUOUcOaMr36EgDh0L5OYI4cbXbYMR8gcDZX1TxGf0hzU
nouJBRIVe43EbRBpT30AwxSOsnxwnGA9bhY3zFQa9SXxTPGzF63RcCeyqdybprow
o/OR6HFZQ7m0vRZfwOMl9JAd+amhPTl5yGE6lk6xloano622hXMCP6ply41iKlJX
kzFOWfGNcktulSY9CZYrqCD2YE1YNm0KIaKOGB+JXE1hH0IRpDoGA1GZKvaFllRK
/o2BZrAFLAQDzYbyLUYGwQDr9IfJzv7iv1uRGMQzmGDE7qhARinI0Vevdg0LRahJ
ZIkZ3hKo/cIz02DXT9NhsHIHC69zfYN7Toc2zhvyK4ODsCwKVeqynCubrsELWmwY
cqWBmVjW0xcFpLSsMUrngJFFFDURZLMCa/vXE9A6ILlJn9wxv6/uAUMO/QI3hdpz
aQm+asSCP2EjHFWmY7pfdfgvF3kDtTztZFtk0da60vdJHrPomCPkusVLh4uDws5W
GYMC5YuHpTeUKyvqUJA+YhuCEuR6207Q1aCfxcXgRb7uIPev8SdjqzzWdHNzOdOn
DI1QeWn1gCTX07whQIJ3L9ITZM4iOgJKaLM2qT2KbeZhneU20wA2bQJVkyMN0Kk6
992XpihmEsdJ351+l2Ln7/cMnawhj4ag/fYkgbBMKA+bgYnWMjzWBGCtwgRGSAOs
hc/jvvE4XmxIP/3gq62TKXxHQOJJFw56QrhRbzsCi8dcFzBIqO3iWaWzj4NNXdEp
KHd6OJwyqTdNioykPQzXKoo1EX1pN4tI7TDD5I+gSIMRhaIbKAXhQ/vqwa2NHlMb
eHwcc9B1xnqFuzBhKNVSEXVut5fU1CTR0ofrcrx4JdWFh6IK7qmgEv+mXnwJyE+8
NpISdwyBkgimoaHeKZqxlo8YQHjeHCMeouJ9HtakmncGMaz1YImgYV1bbekARXJl
0AZo4sAZlTuq5LA/94koPgWEAVGFvOR163EeObQmQ2wfpp1FGR/nA9WfxrZwzkbP
LHM1bswVO5G4jHRI4sjYF9beX1WdHyHzSPZ40l/UaZozGn69ez7i4R3kGL1a2zeg
/dDXqDODgY8WSJSWo/R0xBzOPQShAj6PmuLLperR4UUrcVTMBIMveS2fYvVf9eU3
ASPdsuJmGeGsf3ACYP4fnaE9Iz7+16edBC3TerE64SqP/2GTkpukWZ+2qkgz2MFw
J5QIt3p7gdvur8743yn+03dHnSZjUJLurDlhCfRE6UqaZR3PYpGtzQ/hckUbpm3W
RWNl/PZwgPMSoQkBLG3s41F/dsPSREfgeL5ZjQR22qYcXY7OqVyotpl/F+Rsz4x2
Q90hLoISa3O70u/kH3DK8gBaLcCs32cHPiVenzQw1k1Ywaqy7C3Bb0NHABixDhHR
dj1EUBqXZwDnKfA0xjHC13q1nHUlaGF5aTp/fdJNvX38Nrl2S2u7rOT/KNtykhld
2ZcDnlTL1c1iEqfZxGlHzcxIxuDb6GtM6ziBnq/hxwr6KA04L2yaFMderRPgsQlb
EdFtuc3Uq5X22cqgZtwP6icdJYrEoreT3nQpRNfTPx95nlKwv7VAcdU0Zmmidl1M
0EKLqpkYEHBZO8YOTh7BICHgd14NZlGp8nMflCvRbCj3l3830ylpk5hN1WP2T2K7
Pp3DGTwbMjNBI7MJq3SEDmbaFC2pS1cL3fHy93BlQDGlcMHMmaKEDW44i/YUiijZ
dXJcSXxfBgNaR34miVHbpb4/4VwiSbiciNAvdQPSLGaUy82PnuWksTpWMZWP9DPz
QPPqASoa/4vLQ/01nLME1UFVJdkhjFvt2aymsYJgq6hyqbsNbb90s7a109mSpYj8
UlIH8GvWczAX84zMrj58e+jrxhkfk0dWODnlAq4d5DsLnRIZDbgPZveqgSB0BUc8
5obytuB/XjS4dFDs3hBj5onvARlG0HnHuj1c5efmllWLRmCvs6KhMAZUXPzs22ha
hhuSeiDM2u+a7JE5jI1KAlZwyfcAqoUj0VP75nZbWEv44bj3V4AuxmhrwEA2nBX4
5WBVWsbE3o0TVnTKAWUPY6Hzblu0aOnJMe7C3Lth7wszWbFknanVcULEciabHoPB
T5snq8pQIpZTnrNEBnzbpCctlZqu85ujx10xS6rqXG3Miy5r0YPinAvv+1p6k0zL
V0ocM/3vNBLDqwf4ZaG6z6jMinEwALlKC7HguW7gfUTwLMXEzX7ty3lz9/OnfAv3
0GL+lmz/QHzBml61xWcgFGsh5WQYfazOygdxe7JDQidRRhGbuaalB+adqezNjvWV
zLahEzDaMSw7YdEvkyS9jtV24qsr42QarRkK1Mztgj10+a9roFmpsKWTJTLG1Pum
OFkSSMlATiy7R+XwtJnuUbZOLp4rus0iDYS6+TRiuUDwYRaOf75lwLf5lh3j+9C+
Sudpb4gIGbPgfc34ecN+8sY7F42Ol0XfmtbQUIJ9K5bCrGuMJR/NYujrWZZJHejO
bD5WuBUL9OlZlPyoFz33qO8o0OgU8xT8uqIL7SXcZiRacWK8z1XzmbQA1w501iZi
RfQf0wRkwhEUWED1a/qcdGAe19UC68W6K3mmyKM1OiDL5+j/sK300spXvO8vidkD
y1/iMvnt0rV8WJDlHySU1WDtYPCma/GU+zE68f3ZGhWb+3hxXHO09XUD6Cesgda4
E4nxCHGOOW2DbG7yjYcW1eRoUbOwyBvyhdGWpUjGv/cmzPlJ2jeJoZK4Q47HS82H
gQZQr5PfczHvbuZPEDTM7VK7zkiXxJ8BRfxJmcCkhbPP/bw0VhOwDHi3EhpKb3hL
CdBYsvR7a2G59b3SE6ZQMb048AXtEK8NKEyYDqTXxr9sZSxh3H9qGt1+vxnwFUTC
s0BzSDmrilCkE4UPKpWhBecY8Lm06QfFKAZaFzK+9Q+24KVLdSV/MkB4VtLJu/Bj
tHhkmKpT0SaBx7zIz7uU8HDSUGDIidyfJyApKHK4Mskjv2fkQ5vHiLKonjDXMFQv
EwSQO1tYl8ne7He7w6MtRE0HSVTyniAOD0gEKMESMMwhMZYCyYLGD5MFAyTr1aF1
YAk/k1MmVL9NJ8wrO2JBFdtOl3sxUy7TwbmjATh1P+DZLrPYPhjsFsSaDR53K4rX
BYzEKBTP7hMZDPjJs2jtUb4Y3n+iHlIQ99GIm4O8IVrrUR3fpeeXv8GMap2BQFqT
LGLhoEeOgxeHpHJx+1uwe7+bO+ixayNbxAkmtxCWB98njXcs4bv9S9vOuhFTD3+j
WAPD32L7vwpVLXrjBJyJ3rMy8bkxCltRtIJ091WAPHo+TZjXYTDiarfUTQaI9Q36
W+wUX052tfSwXQ6RexdJuzUIpKhmhlJWttP6sf6DKV8o9M4oR/4sgmRTwc0qc9eb
TMsV0zYBHgnpBAvO6gbKkZSIUr9mGMd6Y/A8o0btA5A02BcRCmlyu2bXzgkzj9pS
nf0JpE8eU5BbKwZptkKxjcXdMCNeT5UzZVSRohSVGCVJSXtEKurDTps+NmoyExl2
OloyNy72Dpzc0c53VSe6B9mzsLeEApX8Vyc9IyLpe9hNkKLPfU1zhoyHScNjqAr/
IZ6AOAI5wcD6hbvBBXk1TIBNc2d/uuwYPeoCM7Dx2WlpUohw7a4XkJAMx5ZjFVzY
qASZrIPHjsFKhaqc/7y8FKbT8v9LUX7+YQd/dTJqck5VZF1YyjPwMUBb5yIIgYy+
XyqykYnUxjHgBIo6c9rsSKUKkxkdKFk0UmRjAqdK+4rdUx6fNUL/rIz3tKbG9R8S
HTI48ZN76D6/PKiLeiq1VXSd15pMZz3C73vQd3sSww5TVJdfByLWCH9q5KB2FVA+
W2b0XvvLTL6q/BR+r2I/1W9fLXIk8U4QyiIpyGnPbk2q91QztNYAstcW+i2Agqyj
mHEQd+Ue/DJxEGlIveZy4W9Srg/7cAxXJn4YdhN0xMaVk97IvBtLhT8uz5jiMyyV
HRw8YqOr8fdf5Afw0LRowtC0gHahrej1JZkc5nr1sBtCZkataKUXktwuNjB3X+FI
bNmItb9DhpufHA3t8ftjnJe5zErwiJ7K9uKBXbnWzmzv1Pz0Z4kuI4qWhKV9no5k
l4Gs3Fbc+sYrjPa8fBQU+o0JugFBg28fdYGtnvII35gpAK+IFyg7Up8xBJG8Kk1L
1D/iqC0qqzFKV6l33x+7C449gTnUikdWXYSe6nHDRrfz1MqWyy5je1LFfm7QKyhr
eLW4d6UWLWPQ42hGfAIJIceyGI4jvkqEOvLoXT0+Z5BYU1LzTTRQ7yVzrutZcZt9
L6USzjijI3yPNCvhPn2AWJfodEKwgpUD9O8caY9enXHGCG8jPr7bnV74pV2ldRrq
1T6QimZ8K38kcwve7JCIQNP1pImBxicA5F7EGBr489W0RfBLKUAlBoJ5U1iSw+pu
Uhl2EDBmfmw2xQdzJuRsYDOXaTwUfLf4z4oAmMDPfxaOKrb+d4nw1KLnQTGq6JcZ
4UaW5bAtmCyYCPYORS98Ht0m65LIilD8kbBhlLpXhr1RopXm8mgSs/OFHWHFsVK9
JX9P13QDwXqpes+luIoSo8+Dw8mSI1MXUrxCFSEw3dqnbscOuJpJe9bIGFjS4bca
XFifPip3NRfkPtLkcg08qWwEVWzH9975TXJ1+37Gq8KUwv8C5VtBB9+N7Mylquva
yaASZOrSX/AADFe0YKP9A4ZbCMlyBW79Vfky5U1FRtdXcGc8qSfGjBGrU2Lp1k6G
00CzYYSDs+USq+YEcs1iiYvEwQTYjbAXXQJK5epPtzKAH27P2UmlDLWPxouatlo9
u9e3nQNhPhzTKA8ln8dNnYtwDqne2/g+bR+sEjysCJgneoKZ07P3k7rWT6xK2U9B
YT72XWjpmlIe2DRZnYOIPrnNRw4Ms6Qod+1T/JNzSATOxHdY36oRB6nZ4KLX8dlA
XGtARKJvd+W0t0Q0zvg7YDNVxFrDb/iibVQ8ZICFNpy44bbyVkU7/Lv6i8gbOgjC
shoOQ+lbsd2E2RM4DLT2r4GEf8vmCQYJIBKkRTYZVRpWm8/rHT9WL/zH0WL5sWMU
o1AAYvpzoTGpfXqr6IpwsURwOsUlJkQZkWrXRwvBIwGMWCzIQbRyb1Odk4SdEhvU
oCrZwSXqX9eCqSqM+9BkrI63aBO2tAPb1PxAC8/zvg2brtP0Q4Le3R1Bw9qz/vx1
kw49kBGiYGm+rRBaBr11UkinsFIEQuA67Q95BBLV8U0YtibNVPZxX6BZeTQMrqzf
lZI+ZDH/KX9/OtzXef8BijBH3rSjOZHZmwWPYzmt0rkRufVouUuVJv9IQ92IcS71
fPq32pauxC9soFRLnFYMfAuvRerv8kjfhA48smPhNtD24uIfVEATgjDiuqwj5/Fl
MEV82bwhJPGTw9/rFwALD55KNlWI6UfMyZvgsNPxBfWxAaF5Qm8UjZa7cgP8ZaU4
JD05fz/bWBPKt0V72Ednaw==
`pragma protect end_protected
